module CHIP( 	
	clk,
    rst_n,
    in_valid,
    D_re,
    D_im,
    out_valid,
    O_re,
    O_im);

input clk,rst_n;
input in_valid;
input [15:0] D_re,D_im;

output out_valid;
output [25:0] O_re,O_im;

wire   C_clk;
wire   C_rst_n;
wire   C_in_valid;
wire  [15:0] C_D_re,C_D_im;

wire  C_out_valid;
wire  [25:0] C_O_re,C_O_im;

wire BUF_clk;
CLKBUFX20 buf0(.A(C_clk),.Y(BUF_clk));

FFT2048 U_FFT(
    .clk(BUF_clk),
    .rst_n(C_rst_n),
    .in_valid(C_in_valid),
    .D_re(C_D_re), 
    .D_im(C_D_im),
    .out_valid(C_out_valid),
	.O_re(C_O_re),
	.O_im(C_O_im)
);

// Input Pads
PDUSDGZ I_CLK(.PAD(clk), .C(C_clk));
PDUSDGZ I_RESET(.PAD(rst_n), .C(C_rst_n));
PDUSDGZ I_IN_VALID(.PAD(in_valid), .C(C_in_valid));
PDUSDGZ I_D_RE_0  (.PAD(D_re[0]),  .C(C_D_re[0]));
PDUSDGZ I_D_RE_1  (.PAD(D_re[1]),  .C(C_D_re[1]));
PDUSDGZ I_D_RE_2  (.PAD(D_re[2]),  .C(C_D_re[2]));
PDUSDGZ I_D_RE_3  (.PAD(D_re[3]),  .C(C_D_re[3]));
PDUSDGZ I_D_RE_4  (.PAD(D_re[4]),  .C(C_D_re[4]));
PDUSDGZ I_D_RE_5  (.PAD(D_re[5]),  .C(C_D_re[5]));
PDUSDGZ I_D_RE_6  (.PAD(D_re[6]),  .C(C_D_re[6]));
PDUSDGZ I_D_RE_7  (.PAD(D_re[7]),  .C(C_D_re[7]));
PDUSDGZ I_D_RE_8  (.PAD(D_re[8]),  .C(C_D_re[8]));
PDUSDGZ I_D_RE_9  (.PAD(D_re[9]),  .C(C_D_re[9]));
PDUSDGZ I_D_RE_10 (.PAD(D_re[10]), .C(C_D_re[10]));
PDUSDGZ I_D_RE_11 (.PAD(D_re[11]), .C(C_D_re[11]));
PDUSDGZ I_D_RE_12 (.PAD(D_re[12]), .C(C_D_re[12]));
PDUSDGZ I_D_RE_13 (.PAD(D_re[13]), .C(C_D_re[13]));
PDUSDGZ I_D_RE_14 (.PAD(D_re[14]), .C(C_D_re[14]));
PDUSDGZ I_D_RE_15 (.PAD(D_re[15]), .C(C_D_re[15]));
PDUSDGZ I_D_IM_0  (.PAD(D_im[0]),  .C(C_D_im[0]));
PDUSDGZ I_D_IM_1  (.PAD(D_im[1]),  .C(C_D_im[1]));
PDUSDGZ I_D_IM_2  (.PAD(D_im[2]),  .C(C_D_im[2]));
PDUSDGZ I_D_IM_3  (.PAD(D_im[3]),  .C(C_D_im[3]));
PDUSDGZ I_D_IM_4  (.PAD(D_im[4]),  .C(C_D_im[4]));
PDUSDGZ I_D_IM_5  (.PAD(D_im[5]),  .C(C_D_im[5]));
PDUSDGZ I_D_IM_6  (.PAD(D_im[6]),  .C(C_D_im[6]));
PDUSDGZ I_D_IM_7  (.PAD(D_im[7]),  .C(C_D_im[7]));
PDUSDGZ I_D_IM_8  (.PAD(D_im[8]),  .C(C_D_im[8]));
PDUSDGZ I_D_IM_9  (.PAD(D_im[9]),  .C(C_D_im[9]));
PDUSDGZ I_D_IM_10 (.PAD(D_im[10]), .C(C_D_im[10]));
PDUSDGZ I_D_IM_11 (.PAD(D_im[11]), .C(C_D_im[11]));
PDUSDGZ I_D_IM_12 (.PAD(D_im[12]), .C(C_D_im[12]));
PDUSDGZ I_D_IM_13 (.PAD(D_im[13]), .C(C_D_im[13]));
PDUSDGZ I_D_IM_14 (.PAD(D_im[14]), .C(C_D_im[14]));
PDUSDGZ I_D_IM_15 (.PAD(D_im[15]), .C(C_D_im[15]));

// Output Pads
PDD08SDGZ O_OUT_VALID(.OEN(1'b0), .I(C_out_valid), .PAD(out_valid), .C());
PDD08SDGZ O_O_RE_0  (.OEN(1'b0), .I(C_O_re[0]),  .PAD(O_re[0]),  .C());
PDD08SDGZ O_O_RE_1  (.OEN(1'b0), .I(C_O_re[1]),  .PAD(O_re[1]),  .C());
PDD08SDGZ O_O_RE_2  (.OEN(1'b0), .I(C_O_re[2]),  .PAD(O_re[2]),  .C());
PDD08SDGZ O_O_RE_3  (.OEN(1'b0), .I(C_O_re[3]),  .PAD(O_re[3]),  .C());
PDD08SDGZ O_O_RE_4  (.OEN(1'b0), .I(C_O_re[4]),  .PAD(O_re[4]),  .C());
PDD08SDGZ O_O_RE_5  (.OEN(1'b0), .I(C_O_re[5]),  .PAD(O_re[5]),  .C());
PDD08SDGZ O_O_RE_6  (.OEN(1'b0), .I(C_O_re[6]),  .PAD(O_re[6]),  .C());
PDD08SDGZ O_O_RE_7  (.OEN(1'b0), .I(C_O_re[7]),  .PAD(O_re[7]),  .C());
PDD08SDGZ O_O_RE_8  (.OEN(1'b0), .I(C_O_re[8]),  .PAD(O_re[8]),  .C());
PDD08SDGZ O_O_RE_9  (.OEN(1'b0), .I(C_O_re[9]),  .PAD(O_re[9]),  .C());
PDD08SDGZ O_O_RE_10 (.OEN(1'b0), .I(C_O_re[10]), .PAD(O_re[10]), .C());
PDD08SDGZ O_O_RE_11 (.OEN(1'b0), .I(C_O_re[11]), .PAD(O_re[11]), .C());
PDD08SDGZ O_O_RE_12 (.OEN(1'b0), .I(C_O_re[12]), .PAD(O_re[12]), .C());
PDD08SDGZ O_O_RE_13 (.OEN(1'b0), .I(C_O_re[13]), .PAD(O_re[13]), .C());
PDD08SDGZ O_O_RE_14 (.OEN(1'b0), .I(C_O_re[14]), .PAD(O_re[14]), .C());
PDD08SDGZ O_O_RE_15 (.OEN(1'b0), .I(C_O_re[15]), .PAD(O_re[15]), .C());
PDD08SDGZ O_O_RE_16 (.OEN(1'b0), .I(C_O_re[16]), .PAD(O_re[16]), .C());
PDD08SDGZ O_O_RE_17 (.OEN(1'b0), .I(C_O_re[17]), .PAD(O_re[17]), .C());
PDD08SDGZ O_O_RE_18 (.OEN(1'b0), .I(C_O_re[18]), .PAD(O_re[18]), .C());
PDD08SDGZ O_O_RE_19 (.OEN(1'b0), .I(C_O_re[19]), .PAD(O_re[19]), .C());
PDD08SDGZ O_O_RE_20 (.OEN(1'b0), .I(C_O_re[20]), .PAD(O_re[20]), .C());
PDD08SDGZ O_O_RE_21 (.OEN(1'b0), .I(C_O_re[21]), .PAD(O_re[21]), .C());
PDD08SDGZ O_O_RE_22 (.OEN(1'b0), .I(C_O_re[22]), .PAD(O_re[22]), .C());
PDD08SDGZ O_O_RE_23 (.OEN(1'b0), .I(C_O_re[23]), .PAD(O_re[23]), .C());
PDD08SDGZ O_O_RE_24 (.OEN(1'b0), .I(C_O_re[24]), .PAD(O_re[24]), .C());
PDD08SDGZ O_O_RE_25 (.OEN(1'b0), .I(C_O_re[25]), .PAD(O_re[25]), .C());
PDD08SDGZ O_O_IM_0  (.OEN(1'b0), .I(C_O_im[0]),  .PAD(O_im[0]),  .C());
PDD08SDGZ O_O_IM_1  (.OEN(1'b0), .I(C_O_im[1]),  .PAD(O_im[1]),  .C());
PDD08SDGZ O_O_IM_2  (.OEN(1'b0), .I(C_O_im[2]),  .PAD(O_im[2]),  .C());
PDD08SDGZ O_O_IM_3  (.OEN(1'b0), .I(C_O_im[3]),  .PAD(O_im[3]),  .C());
PDD08SDGZ O_O_IM_4  (.OEN(1'b0), .I(C_O_im[4]),  .PAD(O_im[4]),  .C());
PDD08SDGZ O_O_IM_5  (.OEN(1'b0), .I(C_O_im[5]),  .PAD(O_im[5]),  .C());
PDD08SDGZ O_O_IM_6  (.OEN(1'b0), .I(C_O_im[6]),  .PAD(O_im[6]),  .C());
PDD08SDGZ O_O_IM_7  (.OEN(1'b0), .I(C_O_im[7]),  .PAD(O_im[7]),  .C());
PDD08SDGZ O_O_IM_8  (.OEN(1'b0), .I(C_O_im[8]),  .PAD(O_im[8]),  .C());
PDD08SDGZ O_O_IM_9  (.OEN(1'b0), .I(C_O_im[9]),  .PAD(O_im[9]),  .C());
PDD08SDGZ O_O_IM_10 (.OEN(1'b0), .I(C_O_im[10]), .PAD(O_im[10]), .C());
PDD08SDGZ O_O_IM_11 (.OEN(1'b0), .I(C_O_im[11]), .PAD(O_im[11]), .C());
PDD08SDGZ O_O_IM_12 (.OEN(1'b0), .I(C_O_im[12]), .PAD(O_im[12]), .C());
PDD08SDGZ O_O_IM_13 (.OEN(1'b0), .I(C_O_im[13]), .PAD(O_im[13]), .C());
PDD08SDGZ O_O_IM_14 (.OEN(1'b0), .I(C_O_im[14]), .PAD(O_im[14]), .C());
PDD08SDGZ O_O_IM_15 (.OEN(1'b0), .I(C_O_im[15]), .PAD(O_im[15]), .C());
PDD08SDGZ O_O_IM_16 (.OEN(1'b0), .I(C_O_im[16]), .PAD(O_im[16]), .C());
PDD08SDGZ O_O_IM_17 (.OEN(1'b0), .I(C_O_im[17]), .PAD(O_im[17]), .C());
PDD08SDGZ O_O_IM_18 (.OEN(1'b0), .I(C_O_im[18]), .PAD(O_im[18]), .C());
PDD08SDGZ O_O_IM_19 (.OEN(1'b0), .I(C_O_im[19]), .PAD(O_im[19]), .C());
PDD08SDGZ O_O_IM_20 (.OEN(1'b0), .I(C_O_im[20]), .PAD(O_im[20]), .C());
PDD08SDGZ O_O_IM_21 (.OEN(1'b0), .I(C_O_im[21]), .PAD(O_im[21]), .C());
PDD08SDGZ O_O_IM_22 (.OEN(1'b0), .I(C_O_im[22]), .PAD(O_im[22]), .C());
PDD08SDGZ O_O_IM_23 (.OEN(1'b0), .I(C_O_im[23]), .PAD(O_im[23]), .C());
PDD08SDGZ O_O_IM_24 (.OEN(1'b0), .I(C_O_im[24]), .PAD(O_im[24]), .C());
PDD08SDGZ O_O_IM_25 (.OEN(1'b0), .I(C_O_im[25]), .PAD(O_im[25]), .C());


// IO power 
PVDD2DGZ VDDP0 ();
PVSS2DGZ GNDP0 ();
PVDD2DGZ VDDP1 ();
PVSS2DGZ GNDP1 ();
PVDD2DGZ VDDP2 ();
PVSS2DGZ GNDP2 ();
PVDD2DGZ VDDP3 ();
PVSS2DGZ GNDP3 ();
PVDD2DGZ VDDP4 ();
PVSS2DGZ GNDP4 ();
PVDD2DGZ VDDP5 ();
PVSS2DGZ GNDP5 ();
PVDD2DGZ VDDP6 ();
PVSS2DGZ GNDP6 ();
PVDD2DGZ VDDP7 ();
PVSS2DGZ GNDP7 ();
PVDD2DGZ VDDP8 ();
PVSS2DGZ GNDP8 ();
PVDD2DGZ VDDP9 ();
PVSS2DGZ GNDP9 ();
PVDD2DGZ VDDP10 ();
PVSS2DGZ GNDP10 ();
PVDD2DGZ VDDP11 ();
PVSS2DGZ GNDP11 ();


// Core power
PVDD1DGZ VDDC0 ();
PVSS1DGZ GNDC0 ();
PVDD1DGZ VDDC1 ();
PVSS1DGZ GNDC1 ();
PVDD1DGZ VDDC2 ();
PVSS1DGZ GNDC2 ();
PVDD1DGZ VDDC3 ();
PVSS1DGZ GNDC3 ();
PVDD1DGZ VDDC4 ();
PVSS1DGZ GNDC4 ();
PVDD1DGZ VDDC5 ();
PVSS1DGZ GNDC5 ();
PVDD1DGZ VDDC6 ();
PVSS1DGZ GNDC6 ();
PVDD1DGZ VDDC7 ();
PVSS1DGZ GNDC7 ();
PVDD1DGZ VDDC8 ();
PVSS1DGZ GNDC8 ();
PVDD1DGZ VDDC9 ();
PVSS1DGZ GNDC9 ();
PVDD1DGZ VDDC10 ();
PVSS1DGZ GNDC10 ();
PVDD1DGZ VDDC11 ();
PVSS1DGZ GNDC11 ();

endmodule

/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Ultra(TM) in wire load mode
// Version   : O-2018.06-SP1
// Date      : Sat Nov 29 17:13:05 2025
/////////////////////////////////////////////////////////////


module FFT2048 ( D_re, D_im, clk, rst_n, in_valid, O_re, O_im, out_valid );
  input [15:0] D_re;
  input [15:0] D_im;
  output [25:0] O_re;
  output [25:0] O_im;
  input clk, rst_n, in_valid;
  output out_valid;
  wire   A3_WEN, A2_WEN, A1_WEN, A0_WEN, A3_CEN, A2_CEN, A1_CEN, A0_CEN,
         OP_done1, A7_WEN, A6_WEN, A5_WEN, A4_WEN, A7_CEN, A6_CEN, A5_CEN,
         A4_CEN, OP2_done0, S_EN, D_sel_reg_4__0_, out_sel, R7_valid,
         U2_valid_1_, U2_factor_reg, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5191, n5193, n5195, n5197, n5199, n5201,
         n5203, n5205, n5207, n5209, n5211, n5213, n5215, n5217, n5219, n5221,
         n5223, n5225, n5227, n5229, n5231, n5233, n5235, n5237, n5239, n5241,
         n5243, n5245, n5247, n5249, n5251, n5253, n5255, n5257, n5259, n5261,
         n5263, n5265, n5267, n5269, n5271, n5273, n5275, n5277, n5279, n5281,
         n5283, n5285, n5287, n5289, n5291, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5638, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5688,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5750, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
         n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
         n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
         n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
         n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
         n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
         n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
         n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
         n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
         n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
         n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
         n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
         n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
         n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
         n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
         n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
         n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
         n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
         n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
         n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
         n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
         n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
         n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
         n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
         n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337,
         n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
         n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
         n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
         n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
         n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
         n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
         n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
         n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
         n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409,
         n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
         n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
         n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553,
         n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
         n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
         n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
         n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
         n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
         n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
         n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
         n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
         n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
         n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769,
         n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
         n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
         n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
         n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
         n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
         n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817,
         n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
         n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
         n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841,
         n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
         n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
         n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
         n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873,
         n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
         n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889,
         n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
         n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
         n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913,
         n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
         n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
         n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
         n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945,
         n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
         n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961,
         n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
         n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
         n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985,
         n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
         n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
         n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
         n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
         n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
         n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
         n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
         n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
         n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057,
         n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105,
         n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
         n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
         n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129,
         n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137,
         n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
         n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
         n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177,
         n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
         n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
         n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201,
         n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
         n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
         n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225,
         n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
         n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
         n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249,
         n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
         n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
         n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
         n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297,
         n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
         n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
         n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321,
         n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329,
         n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
         n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345,
         n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
         n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
         n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369,
         n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
         n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
         n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
         n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417,
         n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
         n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
         n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441,
         n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449,
         n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
         n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465,
         n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473,
         n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481,
         n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489,
         n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
         n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
         n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
         n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
         n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537,
         n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
         n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
         n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561,
         n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
         n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577,
         n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585,
         n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
         n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633,
         n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
         n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
         n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
         n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
         n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
         n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
         n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
         n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
         n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
         n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
         n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
         n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
         n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753,
         n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761,
         n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
         n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
         n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825,
         n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833,
         n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
         n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
         n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
         n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
         n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873,
         n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
         n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
         n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897,
         n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905,
         n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
         n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921,
         n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929,
         n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
         n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945,
         n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
         n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
         n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969,
         n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
         n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
         n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993,
         n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001,
         n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
         n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017,
         n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
         n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
         n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041,
         n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
         n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
         n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065,
         n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073,
         n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081,
         n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089,
         n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097,
         n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
         n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113,
         n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121,
         n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129,
         n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137,
         n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145,
         n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
         n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161,
         n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169,
         n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
         n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185,
         n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193,
         n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
         n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209,
         n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
         n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
         n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233,
         n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
         n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249,
         n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257,
         n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265,
         n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
         n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281,
         n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289,
         n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
         n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305,
         n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313,
         n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
         n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329,
         n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337,
         n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345,
         n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353,
         n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
         n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369,
         n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377,
         n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385,
         n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393,
         n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401,
         n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409,
         n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
         n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425,
         n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
         n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441,
         n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449,
         n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457,
         n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
         n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473,
         n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481,
         n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
         n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
         n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
         n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513,
         n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521,
         n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529,
         n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
         n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545,
         n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553,
         n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
         n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569,
         n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577,
         n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585,
         n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593,
         n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601,
         n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609,
         n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617,
         n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625,
         n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633,
         n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641,
         n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649,
         n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657,
         n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665,
         n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673,
         n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681,
         n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689,
         n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697,
         n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705,
         n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713,
         n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721,
         n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729,
         n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737,
         n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745,
         n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753,
         n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761,
         n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769,
         n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777,
         n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785,
         n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793,
         n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801,
         n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809,
         n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817,
         n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825,
         n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833,
         n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841,
         n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849,
         n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857,
         n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865,
         n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873,
         n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881,
         n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889,
         n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897,
         n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905,
         n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913,
         n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921,
         n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929,
         n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937,
         n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945,
         n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953,
         n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961,
         n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969,
         n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977,
         n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985,
         n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993,
         n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001,
         n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009,
         n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017,
         n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025,
         n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033,
         n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041,
         n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049,
         n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057,
         n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065,
         n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073,
         n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081,
         n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089,
         n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097,
         n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105,
         n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113,
         n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121,
         n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129,
         n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137,
         n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145,
         n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153,
         n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161,
         n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169,
         n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177,
         n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185,
         n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193,
         n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201,
         n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209,
         n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217,
         n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225,
         n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233,
         n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241,
         n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249,
         n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257,
         n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265,
         n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273,
         n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281,
         n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289,
         n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297,
         n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305,
         n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313,
         n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321,
         n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329,
         n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337,
         n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345,
         n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353,
         n26354, n26355, n26356, n26357, n26358, n26359, n26361, n26362,
         n26363, n26364, n26365, n26366, n26367, n26368, n26369, n26370,
         n26371, n26372, n26373, n26374, n26375, n26376, n26377, n26378,
         n26379, n26380, n26381, n26382, n26383, n26384, n26385, n26386,
         n26387, n26388, n26389, n26390, n26391, n26392, n26393, n26394,
         n26395, n26396, n26397, n26398, n26399, n26400, n26401, n26402,
         n26403, n26404, n26405, n26406, n26407, n26408, n26409, n26410,
         n26411, n26412, n26413, n26414, n26415, n26416, n26417, n26418,
         n26419, n26420, n26421, n26422, n26423, n26424, n26425, n26426,
         n26427, n26428, n26429, n26430, n26431, n26432, n26433, n26434,
         n26435, n26436, n26437, n26438, n26439, n26440, n26441, n26442,
         n26443, n26444, n26445, n26446, n26447, n26448, n26449, n26450,
         n26451, n26452, n26453, n26454, n26455, n26456, n26457, n26458,
         n26459, n26460, n26461, n26462, n26463, n26464, n26465, n26466,
         n26467, n26468, n26469, n26470, n26471, n26472, n26473, n26474,
         n26475, n26476, n26477, n26478, n26479, n26480, n26481, n26482,
         n26483, n26484, n26485, n26486, n26487, n26488, n26489, n26490,
         n26491, n26492, n26493, n26494, n26495, n26496, n26497, n26498,
         n26499, n26500, n26501, n26502, n26503, n26504, n26505, n26506,
         n26507, n26508, n26509, n26510, n26511, n26512, n26513, n26514,
         n26515, n26516, n26517, n26518, n26519, n26520, n26521, n26522,
         n26523, n26524, n26525, n26526, n26527, n26528, n26529, n26530,
         n26531, n26532, n26533, n26534, n26535, n26536, n26537, n26538,
         n26539, n26540, n26541, n26542, n26543, n26544, n26545, n26546,
         n26547, n26548, n26549, n26550, n26551, n26552, n26553, n26554,
         n26555, n26556, n26557, n26558, n26559, n26560, n26561, n26562,
         n26563, n26564, n26565, n26566, n26567, n26568, n26569, n26570,
         n26571, n26572, n26573, n26574, n26575, n26576, n26577, n26578,
         n26579, n26580, n26581, n26582, n26583, n26584, n26585, n26586,
         n26587, n26588, n26589, n26590, n26591, n26592, n26593, n26594,
         n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602,
         n26603, n26604, n26605, n26606, n26607, n26608, n26609, n26610,
         n26611, n26612, n26613, n26614, n26615, n26616, n26617, n26618,
         n26619, n26620, n26621, n26622, n26623, n26624, n26625, n26626,
         n26627, n26628, n26629, n26630, n26631, n26632, n26633, n26634,
         n26635, n26636, n26637, n26638, n26639, n26640, n26641, n26642,
         n26643, n26644, n26645, n26646, n26647, n26648, n26649, n26650,
         n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26658,
         n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666,
         n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674,
         n26675, n26676, n26677, n26678, n26679, n26680, n26681, n26682,
         n26683, n26684, n26685, n26686, n26687, n26688, n26689, n26690,
         n26691, n26692, n26693, n26694, n26695, n26696, n26697, n26698,
         n26699, n26700, n26701, n26702, n26703, n26704, n26705, n26706,
         n26707, n26708, n26709, n26710, n26711, n26712, n26713, n26714,
         n26715, n26716, n26717, n26718, n26719, n26720, n26721, n26722,
         n26723, n26724, n26725, n26726, n26727, n26728, n26729, n26730,
         n26731, n26732, n26733, n26734, n26735, n26736, n26737, n26738,
         n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746,
         n26747, n26748, n26749, n26750, n26751, n26752, n26753, n26754,
         n26755, n26756, n26757, n26758, n26759, n26760, n26761, n26762,
         n26763, n26764, n26765, n26766, n26767, n26768, n26769, n26770,
         n26771, n26772, n26773, n26774, n26775, n26776, n26777, n26778,
         n26779, n26780, n26781, n26782, n26783, n26784, n26785, n26786,
         n26787, n26788, n26789, n26790, n26791, n26792, n26793, n26794,
         n26795, n26796, n26797, n26798, n26799, n26800, n26801, n26802,
         n26803, n26804, n26805, n26806, n26807, n26808, n26809, n26810,
         n26811, n26812, n26813, n26814, n26815, n26816, n26817, n26818,
         n26819, n26820, n26821, n26822, n26823, n26824, n26825, n26826,
         n26827, n26828, n26829, n26830, n26831, n26832, n26833, n26834,
         n26835, n26836, n26837, n26838, n26839, n26840, n26841, n26842,
         n26843, n26844, n26845, n26846, n26847, n26848, n26849, n26850,
         n26851, n26852, n26853, n26854, n26855, n26856, n26857, n26858,
         n26859, n26860, n26861, n26862, n26863, n26864, n26865, n26866,
         n26867, n26868, n26869, n26870, n26871, n26872, n26873, n26874,
         n26875, n26876, n26877, n26878, n26879, n26880, n26881, n26882,
         n26883, n26884, n26885, n26886, n26887, n26888, n26889, n26890,
         n26891, n26892, n26893, n26894, n26895, n26896, n26897, n26898,
         n26899, n26900, n26901, n26902, n26903, n26904, n26905, n26906,
         n26907, n26908, n26909, n26910, n26911, n26912, n26913, n26914,
         n26915, n26916, n26917, n26918, n26919, n26920, n26921, n26922,
         n26923, n26924, n26925, n26926, n26927, n26928, n26929, n26930,
         n26931, n26932, n26933, n26934, n26935, n26936, n26937, n26938,
         n26939, n26940, n26941, n26942, n26943, n26944, n26945, n26946,
         n26947, n26948, n26949, n26950, n26951, n26952, n26953, n26954,
         n26955, n26956, n26957, n26958, n26959, n26960, n26961, n26962,
         n26963, n26964, n26965, n26966, n26967, n26968, n26969, n26970,
         n26971, n26972, n26973, n26974, n26975, n26976, n26977, n26978,
         n26979, n26980, n26981, n26982, n26983, n26984, n26985, n26986,
         n26987, n26988, n26989, n26990, n26991, n26992, n26993, n26994,
         n26995, n26996, n26997, n26998, n26999, n27000, n27001, n27002,
         n27003, n27004, n27005, n27006, n27007, n27008, n27009, n27010,
         n27011, n27012, n27013, n27014, n27015, n27016, n27017, n27018,
         n27019, n27020, n27021, n27022, n27023, n27024, n27025, n27026,
         n27027, n27028, n27029, n27030, n27031, n27032, n27033, n27034,
         n27035, n27036, n27037, n27038, n27039, n27040, n27041, n27042,
         n27043, n27044, n27045, n27046, n27047, n27048, n27049, n27050,
         n27051, n27052, n27053, n27054, n27055, n27056, n27057, n27058,
         n27059, n27060, n27061, n27062, n27063, n27064, n27065, n27066,
         n27067, n27068, n27069, n27070, n27071, n27072, n27073, n27074,
         n27075, n27076, n27077, n27078, n27079, n27080, n27081, n27082,
         n27083, n27084, n27085, n27086, n27087, n27088, n27089, n27090,
         n27091, n27092, n27093, n27094, n27095, n27096, n27097, n27098,
         n27099, n27100, n27101, n27102, n27103, n27104, n27105, n27106,
         n27107, n27108, n27109, n27110, n27111, n27112, n27113, n27114,
         n27115, n27116, n27117, n27118, n27119, n27120, n27121, n27122,
         n27123, n27124, n27125, n27126, n27127, n27128, n27129, n27130,
         n27131, n27132, n27133, n27134, n27135, n27136, n27137, n27138,
         n27139, n27140, n27141, n27142, n27143, n27144, n27145, n27146,
         n27147, n27148, n27149, n27150, n27151, n27152, n27153, n27154,
         n27155, n27156, n27157, n27158, n27159, n27160, n27161, n27162,
         n27163, n27164, n27165, n27166, n27167, n27168, n27169, n27170,
         n27171, n27172, n27173, n27174, n27175, n27176, n27177, n27178,
         n27179, n27180, n27181, n27182, n27183, n27184, n27185, n27186,
         n27187, n27188, n27189, n27190, n27191, n27192, n27193, n27194,
         n27195, n27196, n27197, n27198, n27199, n27200, n27201, n27202,
         n27203, n27204, n27205, n27206, n27207, n27208, n27209, n27210,
         n27211, n27212, n27213, n27214, n27215, n27216, n27217, n27218,
         n27219, n27220, n27221, n27222, n27223, n27224, n27225, n27226,
         n27227, n27228, n27229, n27230, n27231, n27232, n27233, n27234,
         n27235, n27236, n27237, n27238, n27239, n27240, n27241, n27242,
         n27243, n27244, n27245, n27246, n27247, n27248, n27249, n27250,
         n27251, n27252, n27253, n27254, n27255, n27256, n27257, n27258,
         n27259, n27260, n27261, n27262, n27263, n27264, n27265, n27266,
         n27267, n27268, n27269, n27270, n27271, n27272, n27273, n27274,
         n27275, n27276, n27277, n27278, n27279, n27280, n27281, n27282,
         n27283, n27284, n27285, n27286, n27287, n27288, n27289, n27290,
         n27291, n27292, n27293, n27294, n27295, n27296, n27297, n27298,
         n27299, n27300, n27301, n27302, n27303, n27304, n27305, n27306,
         n27307, n27308, n27309, n27310, n27311, n27312, n27313, n27314,
         n27315, n27316, n27317, n27318, n27319, n27320, n27321, n27322,
         n27323, n27324, n27325, n27326, n27327, n27328, n27329, n27330,
         n27331, n27332, n27333, n27334, n27335, n27336, n27337, n27338,
         n27339, n27340, n27341, n27342, n27343, n27344, n27345, n27346,
         n27347, n27348, n27349, n27350, n27351, n27352, n27353, n27354,
         n27355, n27356, n27357, n27358, n27359, n27360, n27361, n27362,
         n27363, n27364, n27365, n27366, n27367, n27368, n27369, n27370,
         n27371, n27372, n27373, n27374, n27375, n27376, n27377, n27378,
         n27379, n27380, n27381, n27382, n27383, n27384, n27385, n27386,
         n27387, n27388, n27389, n27390, n27391, n27392, n27393, n27394,
         n27395, n27396, n27397, n27398, n27399, n27400, n27401, n27402,
         n27403, n27404, n27405, n27406, n27407, n27408, n27409, n27410,
         n27411, n27412, n27413, n27414, n27415, n27416, n27417, n27418,
         n27419, n27420, n27421, n27422, n27423, n27424, n27425, n27426,
         n27427, n27428, n27429, n27430, n27431, n27432, n27433, n27434,
         n27435, n27436, n27437, n27438, n27439, n27440, n27441, n27442,
         n27443, n27444, n27445, n27446, n27447, n27448, n27449, n27450,
         n27451, n27452, n27453, n27454, n27455, n27456, n27457, n27458,
         n27459, n27460, n27461, n27462, n27463, n27464, n27465, n27466,
         n27467, n27468, n27469, n27470, n27471, n27472, n27473, n27474,
         n27475, n27476, n27477, n27478, n27479, n27480, n27481, n27482,
         n27483, n27484, n27485, n27486, n27487, n27488, n27489, n27490,
         n27491, n27492, n27493, n27494, n27495, n27496, n27497, n27498,
         n27499, n27500, n27501, n27502, n27503, n27504, n27505, n27506,
         n27507, n27508, n27509, n27510, n27511, n27512, n27513, n27514,
         n27515, n27516, n27517, n27518, n27519, n27520, n27521, n27522,
         n27523, n27524, n27525, n27526, n27527, n27528, n27529, n27530,
         n27531, n27532, n27533, n27534, n27535, n27536, n27537, n27538,
         n27539, n27540, n27541, n27542, n27543, n27544, n27545, n27546,
         n27547, n27548, n27549, n27550, n27551, n27552, n27553, n27554,
         n27555, n27556, n27557, n27558, n27559, n27560, n27561, n27562,
         n27563, n27564, n27565, n27566, n27567, n27568, n27569, n27570,
         n27571, n27572, n27573, n27574, n27575, n27576, n27577, n27578,
         n27579, n27580, n27581, n27582, n27583, n27584, n27585, n27586,
         n27587, n27588, n27589, n27590, n27591, n27592, n27593, n27594,
         n27595, n27596, n27597, n27598, n27599, n27600, n27601, n27602,
         n27603, n27604, n27605, n27606, n27607, n27608, n27609, n27610,
         n27611, n27612, n27613, n27614, n27615, n27616, n27617, n27618,
         n27619, n27620, n27621, n27622, n27623, n27624, n27625, n27626,
         n27627, n27628, n27629, n27630, n27631, n27632, n27633, n27634,
         n27635, n27636, n27637, n27638, n27639, n27640, n27641, n27642,
         n27643, n27644, n27645, n27646, n27647, n27648, n27649, n27650,
         n27651, n27652, n27653, n27654, n27655, n27656, n27657, n27658,
         n27659, n27660, n27661, n27662, n27663, n27664, n27665, n27666,
         n27667, n27668, n27669, n27670, n27671, n27672, n27673, n27674,
         n27675, n27676, n27677, n27678, n27679, n27680, n27681, n27682,
         n27683, n27684, n27685, n27686, n27687, n27688, n27689, n27690,
         n27691, n27692, n27693, n27694, n27695, n27696, n27697, n27698,
         n27699, n27700, n27701, n27702, n27703, n27704, n27705, n27706,
         n27707, n27708, n27709, n27710, n27711, n27712, n27713, n27714,
         n27715, n27716, n27717, n27718, n27719, n27720, n27721, n27722,
         n27723, n27724, n27725, n27726, n27727, n27728, n27729, n27730,
         n27731, n27732, n27733, n27734, n27735, n27736, n27737, n27738,
         n27739, n27740, n27741, n27742, n27743, n27744, n27745, n27746,
         n27747, n27748, n27749, n27750, n27751, n27752, n27753, n27754,
         n27755, n27756, n27757, n27758, n27759, n27760, n27761, n27762,
         n27763, n27764, n27765, n27766, n27767, n27768, n27769, n27770,
         n27771, n27772, n27773, n27774, n27775, n27776, n27777, n27778,
         n27779, n27780, n27781, n27782, n27783, n27784, n27785, n27786,
         n27787, n27788, n27789, n27790, n27791, n27792, n27793, n27794,
         n27795, n27796, n27797, n27798, n27799, n27800, n27801, n27802,
         n27803, n27804, n27805, n27806, n27807, n27808, n27809, n27810,
         n27811, n27812, n27813, n27814, n27815, n27816, n27817, n27818,
         n27819, n27820, n27821, n27822, n27823, n27824, n27825, n27826,
         n27827, n27828, n27829, n27830, n27831, n27832, n27833, n27834,
         n27835, n27836, n27837, n27838, n27839, n27840, n27841, n27842,
         n27843, n27844, n27845, n27846, n27847, n27848, n27849, n27850,
         n27851, n27852, n27853, n27854, n27855, n27856, n27857, n27858,
         n27859, n27860, n27861, n27862, n27863, n27864, n27865, n27866,
         n27867, n27868, n27869, n27870, n27871, n27872, n27873, n27874,
         n27875, n27876, n27877, n27878, n27879, n27880, n27881, n27882,
         n27883, n27884, n27885, n27886, n27887, n27888, n27889, n27890,
         n27891, n27892, n27893, n27894, n27895, n27896, n27897, n27898,
         n27899, n27900, n27901, n27902, n27903, n27904, n27905, n27906,
         n27907, n27908, n27909, n27910, n27911, n27912, n27913, n27914,
         n27915, n27916, n27917, n27918, n27919, n27920, n27921, n27922,
         n27923, n27924, n27925, n27926, n27927, n27928, n27929, n27930,
         n27931, n27932, n27933, n27934, n27935, n27936, n27937, n27938,
         n27939, n27940, n27941, n27942, n27943, n27944, n27945, n27946,
         n27947, n27948, n27949, n27950, n27951, n27952, n27953, n27954,
         n27955, n27956, n27957, n27958, n27959, n27960, n27961, n27962,
         n27963, n27964, n27965, n27966, n27967, n27968, n27969, n27970,
         n27971, n27972, n27973, n27974, n27975, n27976, n27977, n27978,
         n27979, n27980, n27981, n27982, n27983, n27984, n27985, n27986,
         n27987, n27988, n27989, n27990, n27991, n27992, n27993, n27994,
         n27995, n27996, n27997, n27998, n27999, n28000, n28001, n28002,
         n28003, n28004, n28005, n28006, n28007, n28008, n28009, n28010,
         n28011, n28012, n28013, n28014, n28015, n28016, n28017, n28018,
         n28019, n28020, n28021, n28022, n28023, n28024, n28025, n28026,
         n28027, n28028, n28029, n28030, n28031, n28032, n28033, n28034,
         n28035, n28036, n28037, n28038, n28039, n28040, n28041, n28042,
         n28043, n28044, n28045, n28046, n28047, n28048, n28049, n28050,
         n28051, n28052, n28053, n28054, n28055, n28056, n28057, n28058,
         n28059, n28060, n28061, n28062, n28063, n28064, n28065, n28066,
         n28067, n28068, n28069, n28070, n28071, n28072, n28073, n28074,
         n28075, n28076, n28077, n28078, n28079, n28080, n28081, n28082,
         n28083, n28084, n28085, n28086, n28087, n28088, n28089, n28090,
         n28091, n28092, n28093, n28094, n28095, n28096, n28097, n28098,
         n28099, n28100, n28101, n28102, n28103, n28104, n28105, n28106,
         n28107, n28108, n28109, n28110, n28111, n28112, n28113, n28114,
         n28115, n28116, n28117, n28118, n28119, n28120, n28121, n28122,
         n28123, n28124, n28125, n28126, n28127, n28128, n28129, n28130,
         n28131, n28132, n28133, n28134, n28135, n28136, n28137, n28138,
         n28139, n28140, n28141, n28142, n28143, n28144, n28145, n28146,
         n28147, n28148, n28149, n28150, n28151, n28152, n28153, n28154,
         n28155, n28156, n28157, n28158, n28159, n28160, n28161, n28162,
         n28163, n28164, n28165, n28166, n28167, n28168, n28169, n28170,
         n28171, n28172, n28173, n28174, n28175, n28176, n28177, n28178,
         n28179, n28180, n28181, n28182, n28183, n28184, n28185, n28186,
         n28187, n28188, n28189, n28190, n28191, n28192, n28193, n28194,
         n28195, n28196, n28197, n28198, n28199, n28200, n28201, n28202,
         n28203, n28204, n28205, n28206, n28207, n28208, n28209, n28210,
         n28211, n28212, n28213, n28214, n28215, n28216, n28217, n28218,
         n28219, n28220, n28221, n28222, n28223, n28224, n28225, n28226,
         n28227, n28228, n28229, n28230, n28231, n28232, n28233, n28234,
         n28235, n28236, n28237, n28238, n28239, n28240, n28241, n28242,
         n28243, n28244, n28245, n28246, n28247, n28248, n28249, n28250,
         n28251, n28252, n28253, n28254, n28255, n28256, n28257, n28258,
         n28259, n28260, n28261, n28262, n28263, n28264, n28265, n28266,
         n28267, n28268, n28269, n28270, n28271, n28272, n28273, n28274,
         n28275, n28276, n28277, n28278, n28279, n28280, n28281, n28282,
         n28283, n28284, n28285, n28286, n28287, n28288, n28289, n28290,
         n28291, n28292, n28293, n28294, n28295, n28296, n28297, n28298,
         n28299, n28300, n28301, n28302, n28303, n28304, n28305, n28306,
         n28307, n28308, n28309, n28310, n28311, n28312, n28313, n28314,
         n28315, n28316, n28317, n28318, n28319, n28320, n28321, n28322,
         n28323, n28324, n28325, n28326, n28327, n28328, n28329, n28330,
         n28331, n28332, n28333, n28334, n28335, n28336, n28337, n28338,
         n28339, n28340, n28341, n28342, n28343, n28344, n28345, n28346,
         n28347, n28348, n28349, n28350, n28351, n28352, n28353, n28354,
         n28355, n28356, n28357, n28358, n28359, n28360, n28361, n28362,
         n28363, n28364, n28365, n28366, n28367, n28368, n28369, n28370,
         n28371, n28372, n28373, n28374, n28375, n28376, n28377, n28378,
         n28379, n28380, n28381, n28382, n28383, n28384, n28385, n28386,
         n28387, n28388, n28389, n28390, n28391, n28392, n28393, n28394,
         n28395, n28396, n28397, n28398, n28399, n28400, n28401, n28402,
         n28403, n28404, n28405, n28406, n28407, n28408, n28409, n28410,
         n28411, n28412, n28413, n28414, n28415, n28416, n28417, n28418,
         n28419, n28420, n28421, n28422, n28423, n28424, n28425, n28426,
         n28427, n28428, n28429, n28430, n28431, n28432, n28433, n28434,
         n28435, n28436, n28437, n28438, n28439, n28440, n28441, n28442,
         n28443, n28444, n28445, n28446, n28447, n28448, n28449, n28450,
         n28451, n28452, n28453, n28454, n28455, n28456, n28457, n28458,
         n28459, n28460, n28461, n28462, n28463, n28464, n28465, n28466,
         n28467, n28468, n28469, n28470, n28471, n28472, n28473, n28474,
         n28475, n28476, n28477, n28478, n28479, n28480, n28481, n28482,
         n28483, n28484, n28485, n28486, n28487, n28488, n28489, n28490,
         n28491, n28492, n28493, n28494, n28495, n28496, n28497, n28498,
         n28499, n28500, n28501, n28502, n28503, n28504, n28505, n28506,
         n28507, n28508, n28509, n28510, n28511, n28512, n28513, n28514,
         n28515, n28516, n28517, n28518, n28519, n28520, n28521, n28522,
         n28523, n28524, n28525, n28526, n28527, n28528, n28529, n28530,
         n28531, n28532, n28533, n28534, n28535, n28536, n28537, n28538,
         n28539, n28540, n28541, n28542, n28543, n28544, n28545, n28546,
         n28547, n28548, n28549, n28550, n28551, n28552, n28553, n28554,
         n28555, n28556, n28557, n28558, n28559, n28560, n28561, n28562,
         n28563, n28564, n28565, n28566, n28567, n28568, n28569, n28570,
         n28571, n28572, n28573, n28574, n28575, n28576, n28577, n28578,
         n28579, n28580, n28581, n28582, n28583, n28584, n28585, n28586,
         n28587, n28588, n28589, n28590, n28591, n28592, n28593, n28594,
         n28595, n28596, n28597, n28598, n28599, n28600, n28601, n28602,
         n28603, n28604, n28605, n28606, n28607, n28608, n28609, n28610,
         n28611, n28612, n28613, n28614, n28615, n28616, n28617, n28618,
         n28619, n28620, n28621, n28622, n28623, n28624, n28625, n28626,
         n28627, n28628, n28629, n28630, n28631, n28632, n28633, n28634,
         n28635, n28636, n28637, n28638, n28639, n28640, n28641, n28642,
         n28643, n28644, n28645, n28646, n28647, n28648, n28649, n28650,
         n28651, n28652, n28653, n28654, n28655, n28656, n28657, n28658,
         n28659, n28660, n28661, n28662, n28663, n28664, n28665, n28666,
         n28667, n28668, n28669, n28670, n28671, n28672, n28673, n28674,
         n28675, n28676, n28677, n28678, n28679, n28680, n28681, n28682,
         n28683, n28684, n28685, n28686, n28687, n28688, n28689, n28690,
         n28691, n28692, n28693, n28694, n28695, n28696, n28697, n28698,
         n28699, n28700, n28701, n28702, n28703, n28704, n28705, n28706,
         n28707, n28708, n28709, n28710, n28711, n28712, n28713, n28714,
         n28715, n28716, n28717, n28718, n28719, n28720, n28721, n28722,
         n28723, n28724, n28725, n28726, n28727, n28728, n28729, n28730,
         n28731, n28732, n28733, n28734, n28735, n28736, n28737, n28738,
         n28739, n28740, n28741, n28742, n28743, n28744, n28745, n28746,
         n28747, n28748, n28749, n28750, n28751, n28752, n28753, n28754,
         n28755, n28756, n28757, n28758, n28759, n28760, n28761, n28762,
         n28763, n28764, n28765, n28766, n28767, n28768, n28769, n28770,
         n28771, n28772, n28773, n28774, n28775, n28776, n28777, n28778,
         n28779, n28780, n28781, n28782, n28783, n28784, n28785, n28786,
         n28787, n28788, n28789, n28790, n28791, n28792, n28793, n28794,
         n28795, n28796, n28797, n28798, n28799, n28800, n28801, n28802,
         n28803, n28804, n28805, n28806, n28807, n28808, n28809, n28810,
         n28811, n28812, n28813, n28814, n28815, n28816, n28817, n28818,
         n28819, n28820, n28821, n28822, n28823, n28824, n28825, n28826,
         n28827, n28828, n28829, n28830, n28831, n28832, n28833, n28834,
         n28835, n28836, n28837, n28838, n28839, n28840, n28841, n28842,
         n28843, n28844, n28845, n28846, n28847, n28848, n28849, n28850,
         n28851, n28852, n28853, n28854, n28855, n28856, n28857, n28858,
         n28859, n28860, n28861, n28862, n28863, n28864, n28865, n28866,
         n28867, n28868, n28869, n28870, n28871, n28872, n28873, n28874,
         n28875, n28876, n28877, n28878, n28879, n28880, n28881, n28882,
         n28883, n28884, n28885, n28886, n28887, n28888, n28889, n28890,
         n28891, n28892, n28893, n28894, n28895, n28896, n28897, n28898,
         n28899, n28900, n28901, n28902, n28903, n28904, n28905, n28906,
         n28907, n28908, n28909, n28910, n28911, n28912, n28913, n28914,
         n28915, n28916, n28917, n28918, n28919, n28920, n28921, n28922,
         n28923, n28924, n28925, n28926, n28927, n28928, n28929, n28930,
         n28931, n28932, n28933, n28934, n28935, n28936, n28937, n28938,
         n28939, n28940, n28941, n28942, n28943, n28944, n28945, n28946,
         n28947, n28948, n28949, n28950, n28951, n28952, n28953, n28954,
         n28955, n28956, n28957, n28958, n28959, n28960, n28961, n28962,
         n28963, n28964, n28965, n28966, n28967, n28968, n28969, n28970,
         n28971, n28972, n28973, n28974, n28975, n28976, n28977, n28978,
         n28979, n28980, n28981, n28982, n28983, n28984, n28985, n28986,
         n28987, n28988, n28989, n28990, n28991, n28992, n28993, n28994,
         n28995, n28996, n28997, n28998, n28999, n29000, n29001, n29002,
         n29003, n29004, n29005, n29006, n29007, n29008, n29009, n29010,
         n29011, n29012, n29013, n29014, n29015, n29016, n29017, n29018,
         n29019, n29020, n29021, n29022, n29023, n29024, n29025, n29026,
         n29027, n29028, n29029, n29030, n29031, n29032, n29033, n29034,
         n29035, n29036, n29037, n29038, n29039, n29040, n29041, n29042,
         n29043, n29044, n29045, n29046, n29047, n29048, n29049, n29050,
         n29051, n29052, n29053, n29054, n29055, n29056, n29057, n29058,
         n29059, n29060, n29061, n29062, n29063, n29064, n29065, n29066,
         n29067, n29068, n29069, n29070, n29071, n29072, n29073, n29074,
         n29075, n29076, n29077, n29078, n29079, n29080, n29081, n29082,
         n29083, n29084, n29085, n29086, n29087, n29088, n29089, n29090,
         n29091, n29092, n29093, n29094, n29095, n29096, n29097, n29098,
         n29099, n29100, n29101, n29102, n29103, n29104, n29105, n29106,
         n29107, n29108, n29109, n29110, n29111, n29112, n29113, n29114,
         n29115, n29116, n29117, n29118, n29119, n29120, n29121, n29122,
         n29123, n29124, n29125, n29126, n29127, n29128, n29129, n29130,
         n29131, n29132, n29133, n29134, n29135, n29136, n29137, n29138,
         n29139, n29140, n29141, n29142, n29143, n29144, n29145, n29146,
         n29147, n29148, n29149, n29150, n29151, n29152, n29153, n29154,
         n29155, n29156, n29157, n29158, n29159, n29160, n29161, n29162,
         n29163, n29164, n29165, n29166, n29167, n29168, n29169, n29170,
         n29171, n29172, n29173, n29174, n29175, n29176, n29177, n29178,
         n29179, n29180, n29181, n29182, n29183, n29184, n29185, n29186,
         n29187, n29188, n29189, n29190, n29191, n29192, n29193, n29194,
         n29195, n29196, n29197, n29198, n29199, n29200, n29201, n29202,
         n29203, n29204, n29205, n29206, n29207, n29208, n29209, n29210,
         n29211, n29212, n29213, n29214, n29215, n29216, n29217, n29218,
         n29219, n29220, n29221, n29222, n29223, n29224, n29225, n29226,
         n29227, n29228, n29229, n29230, n29231, n29232, n29233, n29234,
         n29235, n29236, n29237, n29238, n29239, n29240, n29241, n29242,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106,
         SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108,
         SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110,
         SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112,
         SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114,
         SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116,
         SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118,
         SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120,
         SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122,
         SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124,
         SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126,
         SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128,
         SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130,
         SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132,
         SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134,
         SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136,
         SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138,
         SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140,
         SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142,
         SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144,
         SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146,
         SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148,
         SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150,
         SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152,
         SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154,
         SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156,
         SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158,
         SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160,
         SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162,
         SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164,
         SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166,
         SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168,
         SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170,
         SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172,
         SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174,
         SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176,
         SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178,
         SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180,
         SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182,
         SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184,
         SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186,
         SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188,
         SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190,
         SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192,
         SYNOPSYS_UNCONNECTED_193, SYNOPSYS_UNCONNECTED_194,
         SYNOPSYS_UNCONNECTED_195, SYNOPSYS_UNCONNECTED_196,
         SYNOPSYS_UNCONNECTED_197, SYNOPSYS_UNCONNECTED_198,
         SYNOPSYS_UNCONNECTED_199, SYNOPSYS_UNCONNECTED_200,
         SYNOPSYS_UNCONNECTED_201, SYNOPSYS_UNCONNECTED_202,
         SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_204,
         SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_206,
         SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_208,
         SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_210,
         SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_212,
         SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_214,
         SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_216,
         SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_218,
         SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_220,
         SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_222,
         SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_224,
         SYNOPSYS_UNCONNECTED_225, SYNOPSYS_UNCONNECTED_226,
         SYNOPSYS_UNCONNECTED_227, SYNOPSYS_UNCONNECTED_228,
         SYNOPSYS_UNCONNECTED_229, SYNOPSYS_UNCONNECTED_230,
         SYNOPSYS_UNCONNECTED_231, SYNOPSYS_UNCONNECTED_232,
         SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_234,
         SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_236,
         SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_238,
         SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_240,
         SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_242,
         SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_244,
         SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_246,
         SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_248,
         SYNOPSYS_UNCONNECTED_249, SYNOPSYS_UNCONNECTED_250,
         SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_252,
         SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_254,
         SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256,
         SYNOPSYS_UNCONNECTED_257, SYNOPSYS_UNCONNECTED_258,
         SYNOPSYS_UNCONNECTED_259, SYNOPSYS_UNCONNECTED_260,
         SYNOPSYS_UNCONNECTED_261, SYNOPSYS_UNCONNECTED_262,
         SYNOPSYS_UNCONNECTED_263, SYNOPSYS_UNCONNECTED_264,
         SYNOPSYS_UNCONNECTED_265, SYNOPSYS_UNCONNECTED_266,
         SYNOPSYS_UNCONNECTED_267, SYNOPSYS_UNCONNECTED_268,
         SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_270,
         SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_272,
         SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_274,
         SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_276,
         SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_278,
         SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_280,
         SYNOPSYS_UNCONNECTED_281, SYNOPSYS_UNCONNECTED_282,
         SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_284,
         SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_286,
         SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_288,
         SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290,
         SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292,
         SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294,
         SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296,
         SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298,
         SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300,
         SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302,
         SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304,
         SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306,
         SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308,
         SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310,
         SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312,
         SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314,
         SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_316,
         SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_318,
         SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_320,
         SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_322,
         SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_324,
         SYNOPSYS_UNCONNECTED_325, SYNOPSYS_UNCONNECTED_326,
         SYNOPSYS_UNCONNECTED_327, SYNOPSYS_UNCONNECTED_328,
         SYNOPSYS_UNCONNECTED_329, SYNOPSYS_UNCONNECTED_330,
         SYNOPSYS_UNCONNECTED_331, SYNOPSYS_UNCONNECTED_332,
         SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_334,
         SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_336,
         SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_338,
         SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340,
         SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342,
         SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344,
         SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346,
         SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348,
         SYNOPSYS_UNCONNECTED_349, SYNOPSYS_UNCONNECTED_350,
         SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_352,
         SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354,
         SYNOPSYS_UNCONNECTED_355, SYNOPSYS_UNCONNECTED_356,
         SYNOPSYS_UNCONNECTED_357, SYNOPSYS_UNCONNECTED_358,
         SYNOPSYS_UNCONNECTED_359, SYNOPSYS_UNCONNECTED_360,
         SYNOPSYS_UNCONNECTED_361, SYNOPSYS_UNCONNECTED_362,
         SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364,
         SYNOPSYS_UNCONNECTED_365, SYNOPSYS_UNCONNECTED_366,
         SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_368,
         SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370,
         SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372,
         SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374,
         SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_376,
         SYNOPSYS_UNCONNECTED_377, SYNOPSYS_UNCONNECTED_378,
         SYNOPSYS_UNCONNECTED_379, SYNOPSYS_UNCONNECTED_380,
         SYNOPSYS_UNCONNECTED_381, SYNOPSYS_UNCONNECTED_382,
         SYNOPSYS_UNCONNECTED_383, SYNOPSYS_UNCONNECTED_384,
         SYNOPSYS_UNCONNECTED_385, SYNOPSYS_UNCONNECTED_386,
         SYNOPSYS_UNCONNECTED_387, SYNOPSYS_UNCONNECTED_388,
         SYNOPSYS_UNCONNECTED_389, SYNOPSYS_UNCONNECTED_390,
         SYNOPSYS_UNCONNECTED_391, SYNOPSYS_UNCONNECTED_392,
         SYNOPSYS_UNCONNECTED_393, SYNOPSYS_UNCONNECTED_394,
         SYNOPSYS_UNCONNECTED_395, SYNOPSYS_UNCONNECTED_396,
         SYNOPSYS_UNCONNECTED_397, SYNOPSYS_UNCONNECTED_398,
         SYNOPSYS_UNCONNECTED_399, SYNOPSYS_UNCONNECTED_400,
         SYNOPSYS_UNCONNECTED_401, SYNOPSYS_UNCONNECTED_402,
         SYNOPSYS_UNCONNECTED_403, SYNOPSYS_UNCONNECTED_404,
         SYNOPSYS_UNCONNECTED_405, SYNOPSYS_UNCONNECTED_406,
         SYNOPSYS_UNCONNECTED_407, SYNOPSYS_UNCONNECTED_408,
         SYNOPSYS_UNCONNECTED_409, SYNOPSYS_UNCONNECTED_410,
         SYNOPSYS_UNCONNECTED_411, SYNOPSYS_UNCONNECTED_412,
         SYNOPSYS_UNCONNECTED_413, SYNOPSYS_UNCONNECTED_414,
         SYNOPSYS_UNCONNECTED_415, SYNOPSYS_UNCONNECTED_416,
         SYNOPSYS_UNCONNECTED_417, SYNOPSYS_UNCONNECTED_418,
         SYNOPSYS_UNCONNECTED_419, SYNOPSYS_UNCONNECTED_420,
         SYNOPSYS_UNCONNECTED_421, SYNOPSYS_UNCONNECTED_422,
         SYNOPSYS_UNCONNECTED_423, SYNOPSYS_UNCONNECTED_424,
         SYNOPSYS_UNCONNECTED_425, SYNOPSYS_UNCONNECTED_426,
         SYNOPSYS_UNCONNECTED_427, SYNOPSYS_UNCONNECTED_428,
         SYNOPSYS_UNCONNECTED_429, SYNOPSYS_UNCONNECTED_430,
         SYNOPSYS_UNCONNECTED_431, SYNOPSYS_UNCONNECTED_432,
         SYNOPSYS_UNCONNECTED_433, SYNOPSYS_UNCONNECTED_434,
         SYNOPSYS_UNCONNECTED_435, SYNOPSYS_UNCONNECTED_436,
         SYNOPSYS_UNCONNECTED_437, SYNOPSYS_UNCONNECTED_438,
         SYNOPSYS_UNCONNECTED_439, SYNOPSYS_UNCONNECTED_440,
         SYNOPSYS_UNCONNECTED_441, SYNOPSYS_UNCONNECTED_442,
         SYNOPSYS_UNCONNECTED_443, SYNOPSYS_UNCONNECTED_444,
         SYNOPSYS_UNCONNECTED_445, SYNOPSYS_UNCONNECTED_446,
         SYNOPSYS_UNCONNECTED_447, SYNOPSYS_UNCONNECTED_448,
         SYNOPSYS_UNCONNECTED_449, SYNOPSYS_UNCONNECTED_450,
         SYNOPSYS_UNCONNECTED_451, SYNOPSYS_UNCONNECTED_452,
         SYNOPSYS_UNCONNECTED_453, SYNOPSYS_UNCONNECTED_454,
         SYNOPSYS_UNCONNECTED_455, SYNOPSYS_UNCONNECTED_456,
         SYNOPSYS_UNCONNECTED_457, SYNOPSYS_UNCONNECTED_458,
         SYNOPSYS_UNCONNECTED_459, SYNOPSYS_UNCONNECTED_460,
         SYNOPSYS_UNCONNECTED_461;
  wire   [9:0] ram_sel_reg;
  wire   [2:0] cs;
  wire   [11:0] cnt;
  wire   [31:0] buffer;
  wire   [4:0] A_sel_reg;
  wire   [3:0] B_sel_reg;
  wire   [9:0] C_sel_reg;
  wire   [51:0] A0_d;
  wire   [51:0] A1_d;
  wire   [51:0] A2_d;
  wire   [51:0] A3_d;
  wire   [51:0] A4_d;
  wire   [51:0] A5_d;
  wire   [51:0] A6_d;
  wire   [51:0] A7_d;
  wire   [7:0] A0_addr;
  wire   [7:0] A1_addr;
  wire   [39:0] Q0_addr;
  wire   [39:0] Q1_addr;
  wire   [7:0] A2_addr;
  wire   [39:0] Q2_addr;
  wire   [39:0] Q3_addr;
  wire   [7:0] A3_addr;
  wire   [51:0] AOPA;
  wire   [51:0] AOPB;
  wire   [51:0] AOPC;
  wire   [51:0] AOPD;
  wire   [51:0] BOPA;
  wire   [51:0] BOPB;
  wire   [51:0] BOPC;
  wire   [51:0] BOPD;
  wire   [30:0] W0;
  wire   [30:0] W1;
  wire   [30:0] W2;
  wire   [30:0] W3;
  wire   [53:0] Q0;
  wire   [53:0] Q1;
  wire   [53:0] Q2;
  wire   [53:0] Q3;
  wire   [53:0] Q4;
  wire   [53:0] Q5;
  wire   [53:0] Q6;
  wire   [53:0] Q7;
  wire   [51:0] CQ0;
  wire   [51:0] CQ1;
  wire   [5:1] B0_addr;
  wire   [6:0] B1_addr;
  wire   [3:1] B2_addr;
  wire   [51:0] DATA0;
  wire   [31:0] T1_rom3_q;
  wire   [31:0] T1_rom2_q;
  wire   [31:0] T1_rom1_q;
  wire   [7:0] T1_rom_addr;
  wire   [31:0] T1_rom0_q;
  wire   [27:0] U0_pipe15;
  wire   [27:0] U0_pipe14;
  wire   [27:0] U0_pipe13;
  wire   [27:0] U0_pipe12;
  wire   [27:0] U0_pipe11;
  wire   [27:0] U0_pipe10;
  wire   [27:0] U0_pipe9;
  wire   [27:0] U0_pipe8;
  wire   [27:0] U0_pipe7;
  wire   [27:0] U0_pipe6;
  wire   [27:0] U0_pipe5;
  wire   [27:0] U0_pipe4;
  wire   [27:0] U0_pipe3;
  wire   [27:0] U0_pipe2;
  wire   [27:0] U0_pipe1;
  wire   [27:0] U0_pipe0;
  wire   [25:0] U2_pipe3;
  wire   [25:0] U2_pipe2;
  wire   [25:0] U2_pipe1;
  wire   [25:0] U2_pipe0;
  wire   [25:0] U2_A_i_d;
  wire   [25:0] U2_A_r_d;
  wire   [25:0] U2_B_i;
  wire   [25:0] U2_B_r;
  wire   [27:0] U1_pipe15;
  wire   [27:0] U1_pipe14;
  wire   [27:0] U1_pipe13;
  wire   [27:0] U1_pipe12;
  wire   [27:0] U1_pipe11;
  wire   [27:0] U1_pipe10;
  wire   [27:0] U1_pipe9;
  wire   [27:0] U1_pipe8;
  wire   [27:0] U1_pipe7;
  wire   [27:0] U1_pipe6;
  wire   [27:0] U1_pipe5;
  wire   [27:0] U1_pipe4;
  wire   [27:0] U1_pipe3;
  wire   [27:0] U1_pipe2;
  wire   [27:0] U1_pipe1;
  wire   [27:0] U1_pipe0;
  wire   [25:0] U1_A_i_d0;
  wire   [25:0] U1_A_r_d0;
  wire   [1:0] U1_valid;
  wire   [40:0] U0_U0_y2;
  wire   [40:0] U0_U0_y1;
  wire   [40:0] U0_U0_y0;
  wire   [16:2] U0_U0_z2;
  wire   [16:0] U0_U0_z1;
  wire   [26:0] U0_U0_z0;
  wire   [39:0] U2_U0_y2;
  wire   [39:0] U2_U0_y1;
  wire   [39:0] U2_U0_y0;
  wire   [16:1] U2_U0_z2;
  wire   [16:0] U2_U0_z1;
  wire   [26:0] U2_U0_z0;
  wire   [40:0] U1_U2_y2;
  wire   [40:0] U1_U2_y1;
  wire   [40:0] U1_U2_y0;
  wire   [16:1] U1_U2_z2;
  wire   [16:0] U1_U2_z1;
  wire   [26:0] U1_U2_z0;
  wire   [40:0] U1_U1_y2;
  wire   [40:0] U1_U1_y1;
  wire   [40:0] U1_U1_y0;
  wire   [16:1] U1_U1_z2;
  wire   [16:0] U1_U1_z1;
  wire   [26:0] U1_U1_z0;
  wire   [40:0] U1_U0_y2;
  wire   [40:0] U1_U0_y1;
  wire   [40:0] U1_U0_y0;
  wire   [26:0] U1_U0_z0;
  wire   [40:0] U0_U2_y2;
  wire   [40:0] U0_U2_y1;
  wire   [40:0] U0_U2_y0;
  wire   [26:0] U0_U2_z0;
  wire   [40:0] U0_U1_y2;
  wire   [40:0] U0_U1_y1;
  wire   [40:0] U0_U1_y0;
  wire   [26:0] U0_U1_z0;
  tri   [51:0] B0_q;
  tri   [51:0] B1_q;
  tri   [51:0] B2_q;
  tri   [51:0] B3_q;
  tri   [51:0] B4_q;
  tri   [51:0] B5_q;
  tri   [51:0] B6_q;
  tri   [51:0] B7_q;

  DRAM_256_52 DS0 ( .QA({SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_46, 
        SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_30, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_51, 
        SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_49, 
        SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_45, 
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_1}), .AA(A0_addr), .DA(
        A0_d), .QB(B0_q), .AB({n29093, n29109, B0_addr[5], n6928, n7124, 
        n29096, B0_addr[1], n6929}), .DB({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CLKA(
        clk), .CENA(A0_CEN), .OENA(1'b0), .WENA(A0_WEN), .CLKB(clk), .CENB(
        n7119), .OENB(1'b0), .WENB(1'b1) );
  DRAM_256_52 DS1 ( .QA({SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_98, 
        SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_95, 
        SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_93, 
        SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_91, 
        SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_89, 
        SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_87, 
        SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_84, 
        SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_82, 
        SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_80, 
        SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_78, 
        SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_76, 
        SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_73, 
        SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_71, 
        SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_69, 
        SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_67, 
        SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_65, 
        SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_62, 
        SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_60, 
        SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_58, 
        SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_56, 
        SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_54, 
        SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_103, 
        SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_101, 
        SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_97, 
        SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_75, 
        SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_53}), .AA(A1_addr), .DA(
        A1_d), .QB(B1_q), .AB({n29093, B1_addr[6], B0_addr[5], n29095, n7124, 
        B1_addr[2], B0_addr[1], B1_addr[0]}), .DB({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CLKA(clk), .CENA(A1_CEN), .OENA(1'b0), .WENA(A1_WEN), .CLKB(clk), .CENB(
        n7119), .OENB(1'b0), .WENB(1'b1) );
  DRAM_256_52 DS2 ( .QA({SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_150, 
        SYNOPSYS_UNCONNECTED_148, SYNOPSYS_UNCONNECTED_147, 
        SYNOPSYS_UNCONNECTED_146, SYNOPSYS_UNCONNECTED_145, 
        SYNOPSYS_UNCONNECTED_144, SYNOPSYS_UNCONNECTED_143, 
        SYNOPSYS_UNCONNECTED_142, SYNOPSYS_UNCONNECTED_141, 
        SYNOPSYS_UNCONNECTED_140, SYNOPSYS_UNCONNECTED_139, 
        SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_136, 
        SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_134, 
        SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_132, 
        SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_130, 
        SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_128, 
        SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_125, 
        SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_123, 
        SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_121, 
        SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_119, 
        SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_117, 
        SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_114, 
        SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_112, 
        SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_110, 
        SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_108, 
        SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_106, 
        SYNOPSYS_UNCONNECTED_156, SYNOPSYS_UNCONNECTED_155, 
        SYNOPSYS_UNCONNECTED_154, SYNOPSYS_UNCONNECTED_153, 
        SYNOPSYS_UNCONNECTED_152, SYNOPSYS_UNCONNECTED_149, 
        SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_127, 
        SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_105}), .AA(A2_addr), 
        .DA(A2_d), .QB(B2_q), .AB({n29094, n29109, n29108, n6928, n7135, 
        n29096, B2_addr[1], n6929}), .DB({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CLKA(
        clk), .CENA(A2_CEN), .OENA(1'b0), .WENA(A2_WEN), .CLKB(clk), .CENB(
        n7119), .OENB(1'b0), .WENB(1'b1) );
  DRAM_256_52 DS3 ( .QA({SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_202, 
        SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_199, 
        SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_197, 
        SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_195, 
        SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_193, 
        SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_191, 
        SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_188, 
        SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_186, 
        SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_184, 
        SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_182, 
        SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_180, 
        SYNOPSYS_UNCONNECTED_178, SYNOPSYS_UNCONNECTED_177, 
        SYNOPSYS_UNCONNECTED_176, SYNOPSYS_UNCONNECTED_175, 
        SYNOPSYS_UNCONNECTED_174, SYNOPSYS_UNCONNECTED_173, 
        SYNOPSYS_UNCONNECTED_172, SYNOPSYS_UNCONNECTED_171, 
        SYNOPSYS_UNCONNECTED_170, SYNOPSYS_UNCONNECTED_169, 
        SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_166, 
        SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_164, 
        SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_162, 
        SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_160, 
        SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_158, 
        SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_207, 
        SYNOPSYS_UNCONNECTED_206, SYNOPSYS_UNCONNECTED_205, 
        SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_201, 
        SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_179, 
        SYNOPSYS_UNCONNECTED_168, SYNOPSYS_UNCONNECTED_157}), .AA(A3_addr), 
        .DA(A3_d), .QB(B3_q), .AB({n29094, B1_addr[6], n29108, n29095, n7135, 
        B1_addr[2], B2_addr[1], B1_addr[0]}), .DB({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CLKA(clk), .CENA(A3_CEN), .OENA(1'b0), .WENA(A3_WEN), .CLKB(clk), .CENB(
        n7119), .OENB(1'b0), .WENB(1'b1) );
  DRAM_256_52 DS4 ( .QA({SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_254, 
        SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_251, 
        SYNOPSYS_UNCONNECTED_250, SYNOPSYS_UNCONNECTED_249, 
        SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_247, 
        SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_245, 
        SYNOPSYS_UNCONNECTED_244, SYNOPSYS_UNCONNECTED_243, 
        SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_240, 
        SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_238, 
        SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_236, 
        SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_234, 
        SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_232, 
        SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_229, 
        SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_227, 
        SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_225, 
        SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_223, 
        SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_221, 
        SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_218, 
        SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_216, 
        SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_214, 
        SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_212, 
        SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_210, 
        SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_259, 
        SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_257, 
        SYNOPSYS_UNCONNECTED_256, SYNOPSYS_UNCONNECTED_253, 
        SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_231, 
        SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_209}), .AA(A0_addr), 
        .DA(A4_d), .QB(B4_q), .AB({n29093, n29109, B0_addr[5], n6928, n7124, 
        n29096, B0_addr[1], n6929}), .DB({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CLKA(
        clk), .CENA(A4_CEN), .OENA(1'b0), .WENA(A4_WEN), .CLKB(clk), .CENB(
        n7119), .OENB(1'b0), .WENB(1'b1) );
  DRAM_256_52 DS5 ( .QA({SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_306, 
        SYNOPSYS_UNCONNECTED_304, SYNOPSYS_UNCONNECTED_303, 
        SYNOPSYS_UNCONNECTED_302, SYNOPSYS_UNCONNECTED_301, 
        SYNOPSYS_UNCONNECTED_300, SYNOPSYS_UNCONNECTED_299, 
        SYNOPSYS_UNCONNECTED_298, SYNOPSYS_UNCONNECTED_297, 
        SYNOPSYS_UNCONNECTED_296, SYNOPSYS_UNCONNECTED_295, 
        SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_292, 
        SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_290, 
        SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_288, 
        SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_286, 
        SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_284, 
        SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_281, 
        SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_279, 
        SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_277, 
        SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_275, 
        SYNOPSYS_UNCONNECTED_274, SYNOPSYS_UNCONNECTED_273, 
        SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_270, 
        SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_268, 
        SYNOPSYS_UNCONNECTED_267, SYNOPSYS_UNCONNECTED_266, 
        SYNOPSYS_UNCONNECTED_265, SYNOPSYS_UNCONNECTED_264, 
        SYNOPSYS_UNCONNECTED_263, SYNOPSYS_UNCONNECTED_262, 
        SYNOPSYS_UNCONNECTED_312, SYNOPSYS_UNCONNECTED_311, 
        SYNOPSYS_UNCONNECTED_310, SYNOPSYS_UNCONNECTED_309, 
        SYNOPSYS_UNCONNECTED_308, SYNOPSYS_UNCONNECTED_305, 
        SYNOPSYS_UNCONNECTED_294, SYNOPSYS_UNCONNECTED_283, 
        SYNOPSYS_UNCONNECTED_272, SYNOPSYS_UNCONNECTED_261}), .AA(A1_addr), 
        .DA(A5_d), .QB(B5_q), .AB({n29093, B1_addr[6], B0_addr[5], n29095, 
        n7124, B1_addr[2], B0_addr[1], B1_addr[0]}), .DB({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .CLKA(clk), .CENA(A5_CEN), .OENA(1'b0), .WENA(A5_WEN), .CLKB(
        clk), .CENB(n7119), .OENB(1'b0), .WENB(1'b1) );
  DRAM_256_52 DS6 ( .QA({SYNOPSYS_UNCONNECTED_359, SYNOPSYS_UNCONNECTED_358, 
        SYNOPSYS_UNCONNECTED_356, SYNOPSYS_UNCONNECTED_355, 
        SYNOPSYS_UNCONNECTED_354, SYNOPSYS_UNCONNECTED_353, 
        SYNOPSYS_UNCONNECTED_352, SYNOPSYS_UNCONNECTED_351, 
        SYNOPSYS_UNCONNECTED_350, SYNOPSYS_UNCONNECTED_349, 
        SYNOPSYS_UNCONNECTED_348, SYNOPSYS_UNCONNECTED_347, 
        SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_344, 
        SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_342, 
        SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_340, 
        SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_338, 
        SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_336, 
        SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_333, 
        SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_331, 
        SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_329, 
        SYNOPSYS_UNCONNECTED_328, SYNOPSYS_UNCONNECTED_327, 
        SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_325, 
        SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_322, 
        SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_320, 
        SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_318, 
        SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_316, 
        SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_314, 
        SYNOPSYS_UNCONNECTED_364, SYNOPSYS_UNCONNECTED_363, 
        SYNOPSYS_UNCONNECTED_362, SYNOPSYS_UNCONNECTED_361, 
        SYNOPSYS_UNCONNECTED_360, SYNOPSYS_UNCONNECTED_357, 
        SYNOPSYS_UNCONNECTED_346, SYNOPSYS_UNCONNECTED_335, 
        SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_313}), .AA(A2_addr), 
        .DA(A6_d), .QB(B6_q), .AB({n29094, n29109, n29108, n6928, n7135, 
        n29096, B2_addr[1], n6929}), .DB({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CLKA(
        clk), .CENA(A6_CEN), .OENA(1'b0), .WENA(A6_WEN), .CLKB(clk), .CENB(
        n7119), .OENB(1'b0), .WENB(1'b1) );
  DRAM_256_52 DS7 ( .QA({SYNOPSYS_UNCONNECTED_411, SYNOPSYS_UNCONNECTED_410, 
        SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_407, 
        SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_405, 
        SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_403, 
        SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_401, 
        SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_399, 
        SYNOPSYS_UNCONNECTED_397, SYNOPSYS_UNCONNECTED_396, 
        SYNOPSYS_UNCONNECTED_395, SYNOPSYS_UNCONNECTED_394, 
        SYNOPSYS_UNCONNECTED_393, SYNOPSYS_UNCONNECTED_392, 
        SYNOPSYS_UNCONNECTED_391, SYNOPSYS_UNCONNECTED_390, 
        SYNOPSYS_UNCONNECTED_389, SYNOPSYS_UNCONNECTED_388, 
        SYNOPSYS_UNCONNECTED_386, SYNOPSYS_UNCONNECTED_385, 
        SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_383, 
        SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_381, 
        SYNOPSYS_UNCONNECTED_380, SYNOPSYS_UNCONNECTED_379, 
        SYNOPSYS_UNCONNECTED_378, SYNOPSYS_UNCONNECTED_377, 
        SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_374, 
        SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_372, 
        SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_370, 
        SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_368, 
        SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_366, 
        SYNOPSYS_UNCONNECTED_416, SYNOPSYS_UNCONNECTED_415, 
        SYNOPSYS_UNCONNECTED_414, SYNOPSYS_UNCONNECTED_413, 
        SYNOPSYS_UNCONNECTED_412, SYNOPSYS_UNCONNECTED_409, 
        SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_387, 
        SYNOPSYS_UNCONNECTED_376, SYNOPSYS_UNCONNECTED_365}), .AA(A3_addr), 
        .DA(A7_d), .QB(B7_q), .AB({n29094, B1_addr[6], n29108, n29095, n7135, 
        B1_addr[2], B2_addr[1], B1_addr[0]}), .DB({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CLKA(clk), .CENA(A7_CEN), .OENA(1'b0), .WENA(A7_WEN), .CLKB(clk), .CENB(
        n7119), .OENB(1'b0), .WENB(1'b1) );
  R2_Wp T1_Wp3 ( .Q(T1_rom3_q), .A(cnt[8:0]), .CLK(clk), .CEN(1'b0) );
  ROM_W3p T1_Wp2 ( .Q(T1_rom2_q), .A({n7132, n7131, T1_rom_addr[5:3], n7078, 
        T1_rom_addr[1:0]}), .CLK(clk), .CEN(1'b0) );
  ROM_W2p T1_Wp1 ( .Q(T1_rom1_q), .A({n7132, n7131, T1_rom_addr[5:3], n7078, 
        n7122, n7121}), .CLK(clk), .CEN(1'b0) );
  ROM_Wp T1_Wp0 ( .Q(T1_rom0_q), .A({n7132, n7131, T1_rom_addr[5:3], n7078, 
        n7122, n7121}), .CLK(clk), .CEN(1'b0) );
  DFFSX1 R_EN_reg ( .D(n11971), .CK(clk), .SN(rst_n), .Q(n28698) );
  DFFSX1 S_EN_reg ( .D(n29241), .CK(clk), .SN(rst_n), .Q(n28986), .QN(S_EN) );
  DFFSX1 cnt_reg_10_ ( .D(n5688), .CK(clk), .SN(rst_n), .Q(n29107), .QN(
        cnt[10]) );
  DFFSX1 valid1_reg_2_ ( .D(n5694), .CK(clk), .SN(rst_n), .Q(n29092) );
  DFFSX1 valid1_reg_1_ ( .D(n29092), .CK(clk), .SN(rst_n), .Q(n28702) );
  DFFSX1 cnt_reg_11_ ( .D(n5680), .CK(clk), .SN(rst_n), .Q(n29012), .QN(
        cnt[11]) );
  DFFSX1 cnt_reg_1_ ( .D(n5678), .CK(clk), .SN(rst_n), .Q(n28705), .QN(cnt[1])
         );
  DFFSX1 cnt_reg_2_ ( .D(n5677), .CK(clk), .SN(rst_n), .Q(n28674), .QN(cnt[2])
         );
  DFFSX4 T1_W3_reg_9_ ( .D(n29113), .CK(clk), .SN(rst_n), .Q(n8045), .QN(W3[9]) );
  DFFSX2 T1_W3_reg_6_ ( .D(n29116), .CK(clk), .SN(rst_n), .Q(n8037), .QN(W3[6]) );
  DFFSX4 T1_W3_reg_5_ ( .D(n29117), .CK(clk), .SN(rst_n), .Q(n8022), .QN(W3[5]) );
  DFFSX4 T1_W3_reg_4_ ( .D(n29118), .CK(clk), .SN(rst_n), .Q(n8030), .QN(W3[4]) );
  DFFSX4 T1_W3_reg_3_ ( .D(n29119), .CK(clk), .SN(rst_n), .Q(n8021), .QN(W3[3]) );
  DFFSX1 T1_W3_reg_31_ ( .D(n29120), .CK(clk), .SN(rst_n), .Q(n7986) );
  DFFSX1 T1_W3_reg_30_ ( .D(n29121), .CK(clk), .SN(rst_n), .QN(W3[30]) );
  DFFSX1 T1_W3_reg_29_ ( .D(n29123), .CK(clk), .SN(rst_n), .QN(W3[29]) );
  DFFSX1 T1_W3_reg_28_ ( .D(n29124), .CK(clk), .SN(rst_n), .QN(W3[28]) );
  DFFSX1 T1_W3_reg_27_ ( .D(n29125), .CK(clk), .SN(rst_n), .QN(W3[27]) );
  DFFSX1 T1_W3_reg_26_ ( .D(n29126), .CK(clk), .SN(rst_n), .QN(W3[26]) );
  DFFSX1 T1_W3_reg_24_ ( .D(n29128), .CK(clk), .SN(rst_n), .QN(W3[24]) );
  DFFSX2 T1_W3_reg_22_ ( .D(n29130), .CK(clk), .SN(rst_n), .QN(W3[22]) );
  DFFSX2 T1_W3_reg_21_ ( .D(n29131), .CK(clk), .SN(rst_n), .QN(W3[21]) );
  DFFSX2 T1_W3_reg_20_ ( .D(n29132), .CK(clk), .SN(rst_n), .QN(W3[20]) );
  DFFSX4 T1_W3_reg_1_ ( .D(n29133), .CK(clk), .SN(rst_n), .Q(n6908), .QN(W3[1]) );
  DFFSX2 T1_W3_reg_18_ ( .D(n29135), .CK(clk), .SN(rst_n), .QN(W3[18]) );
  DFFSX2 T1_W3_reg_16_ ( .D(n29137), .CK(clk), .SN(rst_n), .QN(W3[16]) );
  DFFSX1 T1_W3_reg_14_ ( .D(n29139), .CK(clk), .SN(rst_n), .Q(n7982), .QN(
        W3[14]) );
  DFFSX1 T1_W3_reg_12_ ( .D(n29141), .CK(clk), .SN(rst_n), .Q(n7984), .QN(
        W3[12]) );
  DFFSX1 T1_W3_reg_10_ ( .D(n29143), .CK(clk), .SN(rst_n), .Q(n7985), .QN(
        W3[10]) );
  DFFSX1 cnt_reg_9_ ( .D(n5638), .CK(clk), .SN(rst_n), .Q(n28758), .QN(cnt[9])
         );
  DFFSX1 out_start_reg ( .D(n5695), .CK(clk), .SN(rst_n), .Q(n28699) );
  DFFSX1 out_start0_reg ( .D(n28699), .CK(clk), .SN(rst_n), .Q(n29091) );
  DFFSX4 T1_W0_reg_9_ ( .D(n29209), .CK(clk), .SN(rst_n), .Q(n8048), .QN(W0[9]) );
  DFFSX4 T1_W0_reg_8_ ( .D(n29210), .CK(clk), .SN(rst_n), .Q(n7998), .QN(W0[8]) );
  DFFSX4 T1_W0_reg_7_ ( .D(n29211), .CK(clk), .SN(rst_n), .Q(n8043), .QN(W0[7]) );
  DFFSX4 T1_W0_reg_6_ ( .D(n29212), .CK(clk), .SN(rst_n), .Q(n8039), .QN(W0[6]) );
  DFFSX4 T1_W0_reg_5_ ( .D(n29213), .CK(clk), .SN(rst_n), .Q(n7945), .QN(W0[5]) );
  DFFSX4 T1_W0_reg_4_ ( .D(n29214), .CK(clk), .SN(rst_n), .Q(n8014), .QN(W0[4]) );
  DFFSX4 T1_W0_reg_3_ ( .D(n29215), .CK(clk), .SN(rst_n), .Q(n8026), .QN(W0[3]) );
  DFFSX1 T1_W0_reg_31_ ( .D(n29216), .CK(clk), .SN(rst_n), .Q(n7987), .QN(
        n6898) );
  DFFSX1 T1_W0_reg_30_ ( .D(n29217), .CK(clk), .SN(rst_n), .QN(W0[30]) );
  DFFSX2 T1_W0_reg_29_ ( .D(n29219), .CK(clk), .SN(rst_n), .QN(W0[29]) );
  DFFSX2 T1_W0_reg_28_ ( .D(n29220), .CK(clk), .SN(rst_n), .QN(W0[28]) );
  DFFSX2 T1_W0_reg_27_ ( .D(n29221), .CK(clk), .SN(rst_n), .QN(W0[27]) );
  DFFSX4 T1_W0_reg_26_ ( .D(n29222), .CK(clk), .SN(rst_n), .QN(W0[26]) );
  DFFSX4 T1_W0_reg_24_ ( .D(n29224), .CK(clk), .SN(rst_n), .QN(W0[24]) );
  DFFSX4 T1_W0_reg_22_ ( .D(n29226), .CK(clk), .SN(rst_n), .QN(W0[22]) );
  DFFSX4 T1_W0_reg_21_ ( .D(n29227), .CK(clk), .SN(rst_n), .QN(W0[21]) );
  DFFSX4 T1_W0_reg_20_ ( .D(n29228), .CK(clk), .SN(rst_n), .QN(W0[20]) );
  DFFSX4 T1_W0_reg_1_ ( .D(n29229), .CK(clk), .SN(rst_n), .Q(n8029), .QN(W0[1]) );
  DFFSX4 T1_W0_reg_18_ ( .D(n29231), .CK(clk), .SN(rst_n), .QN(W0[18]) );
  DFFSX4 T1_W0_reg_17_ ( .D(n29232), .CK(clk), .SN(rst_n), .QN(W0[17]) );
  DFFSX4 T1_W0_reg_16_ ( .D(n29233), .CK(clk), .SN(rst_n), .QN(W0[16]) );
  DFFSX1 T1_W0_reg_15_ ( .D(n29234), .CK(clk), .SN(rst_n), .Q(n8006), .QN(
        n6897) );
  DFFSX4 T1_W0_reg_13_ ( .D(n29236), .CK(clk), .SN(rst_n), .Q(n8005), .QN(
        W0[13]) );
  DFFSX4 T1_W0_reg_12_ ( .D(n29237), .CK(clk), .SN(rst_n), .Q(n7973), .QN(
        W0[12]) );
  DFFSX4 T1_W0_reg_11_ ( .D(n29238), .CK(clk), .SN(rst_n), .Q(n8025), .QN(
        W0[11]) );
  DFFSX4 T1_W0_reg_10_ ( .D(n29239), .CK(clk), .SN(rst_n), .Q(n7951), .QN(
        W0[10]) );
  DFFSX4 T1_W0_reg_0_ ( .D(n29240), .CK(clk), .SN(rst_n), .Q(n8013), .QN(W0[0]) );
  DFFSX4 T1_W1_reg_8_ ( .D(n29178), .CK(clk), .SN(rst_n), .Q(n8017), .QN(W1[8]) );
  DFFSX4 T1_W1_reg_7_ ( .D(n29179), .CK(clk), .SN(rst_n), .Q(n7950), .QN(W1[7]) );
  DFFSX4 T1_W1_reg_6_ ( .D(n29180), .CK(clk), .SN(rst_n), .Q(n8038), .QN(W1[6]) );
  DFFSX4 T1_W1_reg_5_ ( .D(n29181), .CK(clk), .SN(rst_n), .Q(n7949), .QN(W1[5]) );
  DFFSX4 T1_W1_reg_4_ ( .D(n29182), .CK(clk), .SN(rst_n), .Q(n8020), .QN(W1[4]) );
  DFFSX4 T1_W1_reg_3_ ( .D(n29183), .CK(clk), .SN(rst_n), .Q(n7996), .QN(W1[3]) );
  DFFSX1 T1_W1_reg_31_ ( .D(n29184), .CK(clk), .SN(rst_n), .Q(n7976), .QN(
        n6933) );
  DFFSX1 T1_W1_reg_30_ ( .D(n29185), .CK(clk), .SN(rst_n), .QN(W1[30]) );
  DFFSX4 T1_W1_reg_2_ ( .D(n29186), .CK(clk), .SN(rst_n), .Q(n8041), .QN(W1[2]) );
  DFFSX1 T1_W1_reg_29_ ( .D(n29187), .CK(clk), .SN(rst_n), .QN(W1[29]) );
  DFFSX2 T1_W1_reg_28_ ( .D(n29188), .CK(clk), .SN(rst_n), .QN(W1[28]) );
  DFFSX2 T1_W1_reg_26_ ( .D(n29190), .CK(clk), .SN(rst_n), .QN(W1[26]) );
  DFFSX4 T1_W1_reg_22_ ( .D(n29194), .CK(clk), .SN(rst_n), .QN(W1[22]) );
  DFFSX4 T1_W1_reg_21_ ( .D(n29195), .CK(clk), .SN(rst_n), .QN(W1[21]) );
  DFFSX4 T1_W1_reg_20_ ( .D(n29196), .CK(clk), .SN(rst_n), .QN(W1[20]) );
  DFFSX4 T1_W1_reg_1_ ( .D(n29197), .CK(clk), .SN(rst_n), .Q(n8040), .QN(W1[1]) );
  DFFSX4 T1_W1_reg_17_ ( .D(n29200), .CK(clk), .SN(rst_n), .QN(W1[17]) );
  DFFSX4 T1_W1_reg_16_ ( .D(n29201), .CK(clk), .SN(rst_n), .QN(W1[16]) );
  DFFSX1 T1_W1_reg_15_ ( .D(n29202), .CK(clk), .SN(rst_n), .Q(n7959), .QN(
        W1[15]) );
  DFFSX4 T1_W1_reg_13_ ( .D(n29204), .CK(clk), .SN(rst_n), .Q(n8007), .QN(
        W1[13]) );
  DFFSX4 T1_W1_reg_0_ ( .D(n29208), .CK(clk), .SN(rst_n), .Q(n8009), .QN(W1[0]) );
  DFFSX4 T1_W2_reg_9_ ( .D(n29145), .CK(clk), .SN(rst_n), .Q(n8047), .QN(W2[9]) );
  DFFSX4 T1_W2_reg_8_ ( .D(n29146), .CK(clk), .SN(rst_n), .Q(n8011), .QN(W2[8]) );
  DFFSX4 T1_W2_reg_7_ ( .D(n29147), .CK(clk), .SN(rst_n), .Q(n8042), .QN(W2[7]) );
  DFFSX4 T1_W2_reg_6_ ( .D(n29148), .CK(clk), .SN(rst_n), .Q(n7946), .QN(W2[6]) );
  DFFSX4 T1_W2_reg_5_ ( .D(n29149), .CK(clk), .SN(rst_n), .Q(n7942), .QN(W2[5]) );
  DFFSX4 T1_W2_reg_4_ ( .D(n29150), .CK(clk), .SN(rst_n), .Q(n7980), .QN(W2[4]) );
  DFFSX4 T1_W2_reg_3_ ( .D(n29151), .CK(clk), .SN(rst_n), .Q(n8027), .QN(W2[3]) );
  DFFSX1 T1_W2_reg_31_ ( .D(n29152), .CK(clk), .SN(rst_n), .Q(n7978), .QN(
        n6943) );
  DFFSX1 T1_W2_reg_30_ ( .D(n29153), .CK(clk), .SN(rst_n), .QN(W2[30]) );
  DFFSX4 T1_W2_reg_2_ ( .D(n29154), .CK(clk), .SN(rst_n), .Q(n7947), .QN(W2[2]) );
  DFFSX2 T1_W2_reg_29_ ( .D(n29155), .CK(clk), .SN(rst_n), .QN(W2[29]) );
  DFFSX2 T1_W2_reg_28_ ( .D(n29156), .CK(clk), .SN(rst_n), .QN(W2[28]) );
  DFFSX4 T1_W2_reg_25_ ( .D(n29159), .CK(clk), .SN(rst_n), .QN(W2[25]) );
  DFFSX4 T1_W2_reg_24_ ( .D(n29160), .CK(clk), .SN(rst_n), .QN(W2[24]) );
  DFFSX4 T1_W2_reg_22_ ( .D(n29162), .CK(clk), .SN(rst_n), .QN(W2[22]) );
  DFFSX4 T1_W2_reg_21_ ( .D(n29163), .CK(clk), .SN(rst_n), .Q(n5758), .QN(
        W2[21]) );
  DFFSX4 T1_W2_reg_20_ ( .D(n29164), .CK(clk), .SN(rst_n), .QN(W2[20]) );
  DFFSX4 T1_W2_reg_1_ ( .D(n29165), .CK(clk), .SN(rst_n), .Q(n8028), .QN(W2[1]) );
  DFFSX4 T1_W2_reg_19_ ( .D(n29166), .CK(clk), .SN(rst_n), .QN(W2[19]) );
  DFFSX4 T1_W2_reg_18_ ( .D(n29167), .CK(clk), .SN(rst_n), .QN(W2[18]) );
  DFFSX4 T1_W2_reg_17_ ( .D(n29168), .CK(clk), .SN(rst_n), .QN(W2[17]) );
  DFFSX4 T1_W2_reg_16_ ( .D(n29169), .CK(clk), .SN(rst_n), .QN(W2[16]) );
  DFFSX4 T1_W2_reg_13_ ( .D(n29172), .CK(clk), .SN(rst_n), .Q(n8031), .QN(
        W2[13]) );
  DFFSX4 T1_W2_reg_10_ ( .D(n29175), .CK(clk), .SN(rst_n), .Q(n7974), .QN(
        W2[10]) );
  DFFSX4 T1_W2_reg_0_ ( .D(n29176), .CK(clk), .SN(rst_n), .Q(n8008), .QN(W2[0]) );
  DFFSX1 valid_reg_2_ ( .D(n5693), .CK(clk), .SN(rst_n), .Q(n29090) );
  DFFSX1 valid_reg_1_ ( .D(n29090), .CK(clk), .SN(rst_n), .Q(n28701) );
  DFFSX1 U1_valid_reg_0_ ( .D(n28701), .CK(clk), .SN(rst_n), .Q(n8053), .QN(
        U1_valid[0]) );
  DFFSX1 Q3_addr_reg_4__0_ ( .D(n5536), .CK(clk), .SN(rst_n), .QN(Q3_addr[32])
         );
  DFFSX1 Q3_addr_reg_4__1_ ( .D(n5535), .CK(clk), .SN(rst_n), .QN(Q3_addr[33])
         );
  DFFSX1 Q3_addr_reg_4__2_ ( .D(n5534), .CK(clk), .SN(rst_n), .QN(Q3_addr[34])
         );
  DFFSX1 Q3_addr_reg_4__3_ ( .D(n5533), .CK(clk), .SN(rst_n), .QN(Q3_addr[35])
         );
  DFFSX1 Q3_addr_reg_4__4_ ( .D(n5532), .CK(clk), .SN(rst_n), .QN(Q3_addr[36])
         );
  DFFSX1 Q3_addr_reg_4__5_ ( .D(n5531), .CK(clk), .SN(rst_n), .QN(Q3_addr[37])
         );
  DFFSX1 Q1_addr_reg_4__0_ ( .D(n5530), .CK(clk), .SN(rst_n), .QN(Q1_addr[32])
         );
  DFFSX1 Q1_addr_reg_3__0_ ( .D(n5529), .CK(clk), .SN(rst_n), .QN(Q1_addr[24])
         );
  DFFSX1 Q1_addr_reg_2__0_ ( .D(n5528), .CK(clk), .SN(rst_n), .QN(Q1_addr[16])
         );
  DFFSX1 Q1_addr_reg_1__0_ ( .D(n5527), .CK(clk), .SN(rst_n), .QN(Q1_addr[8])
         );
  DFFSX1 Q1_addr_reg_0__0_ ( .D(n5526), .CK(clk), .SN(rst_n), .Q(n28752), .QN(
        Q1_addr[0]) );
  DFFSX1 Q1_addr_reg_4__1_ ( .D(n5525), .CK(clk), .SN(rst_n), .QN(Q1_addr[33])
         );
  DFFSX1 Q1_addr_reg_3__1_ ( .D(n5524), .CK(clk), .SN(rst_n), .QN(Q1_addr[25])
         );
  DFFSX1 Q1_addr_reg_2__1_ ( .D(n5523), .CK(clk), .SN(rst_n), .QN(Q1_addr[17])
         );
  DFFSX1 Q1_addr_reg_1__1_ ( .D(n5522), .CK(clk), .SN(rst_n), .QN(Q1_addr[9])
         );
  DFFSX1 Q1_addr_reg_0__1_ ( .D(n5521), .CK(clk), .SN(rst_n), .Q(n28753), .QN(
        Q1_addr[1]) );
  DFFSX1 Q1_addr_reg_4__2_ ( .D(n5520), .CK(clk), .SN(rst_n), .QN(Q1_addr[34])
         );
  DFFSX1 Q1_addr_reg_3__2_ ( .D(n5519), .CK(clk), .SN(rst_n), .QN(Q1_addr[26])
         );
  DFFSX1 Q1_addr_reg_2__2_ ( .D(n5518), .CK(clk), .SN(rst_n), .QN(Q1_addr[18])
         );
  DFFSX1 Q1_addr_reg_1__2_ ( .D(n5517), .CK(clk), .SN(rst_n), .QN(Q1_addr[10])
         );
  DFFSX1 Q1_addr_reg_0__2_ ( .D(n5516), .CK(clk), .SN(rst_n), .Q(n28755), .QN(
        Q1_addr[2]) );
  DFFSX1 Q1_addr_reg_4__3_ ( .D(n5515), .CK(clk), .SN(rst_n), .QN(Q1_addr[35])
         );
  DFFSX1 Q1_addr_reg_3__3_ ( .D(n5514), .CK(clk), .SN(rst_n), .QN(Q1_addr[27])
         );
  DFFSX1 Q1_addr_reg_2__3_ ( .D(n5513), .CK(clk), .SN(rst_n), .QN(Q1_addr[19])
         );
  DFFSX1 Q1_addr_reg_1__3_ ( .D(n5512), .CK(clk), .SN(rst_n), .QN(Q1_addr[11])
         );
  DFFSX1 Q1_addr_reg_0__3_ ( .D(n5511), .CK(clk), .SN(rst_n), .Q(n28756), .QN(
        Q1_addr[3]) );
  DFFSX1 Q1_addr_reg_4__4_ ( .D(n5510), .CK(clk), .SN(rst_n), .QN(Q1_addr[36])
         );
  DFFSX1 Q1_addr_reg_3__4_ ( .D(n5509), .CK(clk), .SN(rst_n), .QN(Q1_addr[28])
         );
  DFFSX1 Q1_addr_reg_2__4_ ( .D(n5508), .CK(clk), .SN(rst_n), .QN(Q1_addr[20])
         );
  DFFSX1 Q1_addr_reg_1__4_ ( .D(n5507), .CK(clk), .SN(rst_n), .QN(Q1_addr[12])
         );
  DFFSX1 Q1_addr_reg_0__4_ ( .D(n5506), .CK(clk), .SN(rst_n), .Q(n28754), .QN(
        Q1_addr[4]) );
  DFFSX1 Q0_addr_reg_4__0_ ( .D(n5505), .CK(clk), .SN(rst_n), .QN(Q0_addr[32])
         );
  DFFSX1 Q0_addr_reg_3__0_ ( .D(n5504), .CK(clk), .SN(rst_n), .QN(Q0_addr[24])
         );
  DFFSX1 Q0_addr_reg_4__1_ ( .D(n5503), .CK(clk), .SN(rst_n), .QN(Q0_addr[33])
         );
  DFFSX1 Q0_addr_reg_3__1_ ( .D(n5502), .CK(clk), .SN(rst_n), .QN(Q0_addr[25])
         );
  DFFSX1 Q0_addr_reg_4__2_ ( .D(n5501), .CK(clk), .SN(rst_n), .QN(Q0_addr[34])
         );
  DFFSX1 Q0_addr_reg_3__2_ ( .D(n5500), .CK(clk), .SN(rst_n), .QN(Q0_addr[26])
         );
  DFFSX1 Q0_addr_reg_4__3_ ( .D(n5499), .CK(clk), .SN(rst_n), .QN(Q0_addr[35])
         );
  DFFSX1 Q0_addr_reg_3__3_ ( .D(n5498), .CK(clk), .SN(rst_n), .QN(Q0_addr[27])
         );
  DFFSX1 Q3_addr_reg_3__0_ ( .D(n5497), .CK(clk), .SN(rst_n), .QN(Q3_addr[24])
         );
  DFFSX1 Q3_addr_reg_2__0_ ( .D(n5496), .CK(clk), .SN(rst_n), .QN(Q3_addr[16])
         );
  DFFSX1 Q3_addr_reg_1__0_ ( .D(n5495), .CK(clk), .SN(rst_n), .QN(Q3_addr[8])
         );
  DFFSX1 Q3_addr_reg_0__0_ ( .D(n5494), .CK(clk), .SN(rst_n), .QN(Q3_addr[0])
         );
  DFFSX1 Q3_addr_reg_3__1_ ( .D(n5493), .CK(clk), .SN(rst_n), .QN(Q3_addr[25])
         );
  DFFSX1 Q3_addr_reg_2__1_ ( .D(n5492), .CK(clk), .SN(rst_n), .QN(Q3_addr[17])
         );
  DFFSX1 Q3_addr_reg_1__1_ ( .D(n5491), .CK(clk), .SN(rst_n), .QN(Q3_addr[9])
         );
  DFFSX1 Q3_addr_reg_0__1_ ( .D(n5490), .CK(clk), .SN(rst_n), .QN(Q3_addr[1])
         );
  DFFSX1 Q3_addr_reg_3__2_ ( .D(n5489), .CK(clk), .SN(rst_n), .QN(Q3_addr[26])
         );
  DFFSX1 Q3_addr_reg_2__2_ ( .D(n5488), .CK(clk), .SN(rst_n), .QN(Q3_addr[18])
         );
  DFFSX1 Q3_addr_reg_1__2_ ( .D(n5487), .CK(clk), .SN(rst_n), .QN(Q3_addr[10])
         );
  DFFSX1 Q3_addr_reg_0__2_ ( .D(n5486), .CK(clk), .SN(rst_n), .QN(Q3_addr[2])
         );
  DFFSX1 Q3_addr_reg_3__3_ ( .D(n5485), .CK(clk), .SN(rst_n), .QN(Q3_addr[27])
         );
  DFFSX1 Q3_addr_reg_2__3_ ( .D(n5484), .CK(clk), .SN(rst_n), .QN(Q3_addr[19])
         );
  DFFSX1 Q3_addr_reg_1__3_ ( .D(n5483), .CK(clk), .SN(rst_n), .QN(Q3_addr[11])
         );
  DFFSX1 Q3_addr_reg_0__3_ ( .D(n5482), .CK(clk), .SN(rst_n), .QN(Q3_addr[3])
         );
  DFFSX1 Q3_addr_reg_3__4_ ( .D(n5481), .CK(clk), .SN(rst_n), .QN(Q3_addr[28])
         );
  DFFSX1 Q3_addr_reg_2__4_ ( .D(n5480), .CK(clk), .SN(rst_n), .QN(Q3_addr[20])
         );
  DFFSX1 Q3_addr_reg_1__4_ ( .D(n5479), .CK(clk), .SN(rst_n), .QN(Q3_addr[12])
         );
  DFFSX1 Q3_addr_reg_0__4_ ( .D(n5478), .CK(clk), .SN(rst_n), .QN(Q3_addr[4])
         );
  DFFSX1 Q3_addr_reg_3__5_ ( .D(n5477), .CK(clk), .SN(rst_n), .QN(Q3_addr[29])
         );
  DFFSX1 Q3_addr_reg_2__5_ ( .D(n5476), .CK(clk), .SN(rst_n), .QN(Q3_addr[21])
         );
  DFFSX1 Q3_addr_reg_1__5_ ( .D(n5475), .CK(clk), .SN(rst_n), .QN(Q3_addr[13])
         );
  DFFSX1 Q3_addr_reg_0__5_ ( .D(n5474), .CK(clk), .SN(rst_n), .QN(Q3_addr[5])
         );
  DFFSX1 Q2_addr_reg_4__0_ ( .D(n5473), .CK(clk), .SN(rst_n), .QN(Q2_addr[32])
         );
  DFFSX1 Q2_addr_reg_3__0_ ( .D(n5472), .CK(clk), .SN(rst_n), .QN(Q2_addr[24])
         );
  DFFSX1 Q2_addr_reg_2__0_ ( .D(n5471), .CK(clk), .SN(rst_n), .QN(Q2_addr[16])
         );
  DFFSX1 Q2_addr_reg_1__0_ ( .D(n5470), .CK(clk), .SN(rst_n), .QN(Q2_addr[8])
         );
  DFFSX1 Q2_addr_reg_0__0_ ( .D(n5469), .CK(clk), .SN(rst_n), .QN(Q2_addr[0])
         );
  DFFSX1 Q2_addr_reg_4__1_ ( .D(n5468), .CK(clk), .SN(rst_n), .QN(Q2_addr[33])
         );
  DFFSX1 Q2_addr_reg_3__1_ ( .D(n5467), .CK(clk), .SN(rst_n), .QN(Q2_addr[25])
         );
  DFFSX1 Q2_addr_reg_2__1_ ( .D(n5466), .CK(clk), .SN(rst_n), .QN(Q2_addr[17])
         );
  DFFSX1 Q2_addr_reg_1__1_ ( .D(n5465), .CK(clk), .SN(rst_n), .QN(Q2_addr[9])
         );
  DFFSX1 Q2_addr_reg_0__1_ ( .D(n5464), .CK(clk), .SN(rst_n), .QN(Q2_addr[1])
         );
  DFFSX1 Q2_addr_reg_4__2_ ( .D(n5463), .CK(clk), .SN(rst_n), .QN(Q2_addr[34])
         );
  DFFSX1 Q2_addr_reg_3__2_ ( .D(n5462), .CK(clk), .SN(rst_n), .QN(Q2_addr[26])
         );
  DFFSX1 Q2_addr_reg_2__2_ ( .D(n5461), .CK(clk), .SN(rst_n), .QN(Q2_addr[18])
         );
  DFFSX1 Q2_addr_reg_1__2_ ( .D(n5460), .CK(clk), .SN(rst_n), .QN(Q2_addr[10])
         );
  DFFSX1 Q2_addr_reg_0__2_ ( .D(n5459), .CK(clk), .SN(rst_n), .QN(Q2_addr[2])
         );
  DFFSX1 Q2_addr_reg_4__3_ ( .D(n5458), .CK(clk), .SN(rst_n), .QN(Q2_addr[35])
         );
  DFFSX1 Q2_addr_reg_3__3_ ( .D(n5457), .CK(clk), .SN(rst_n), .QN(Q2_addr[27])
         );
  DFFSX1 Q2_addr_reg_2__3_ ( .D(n5456), .CK(clk), .SN(rst_n), .QN(Q2_addr[19])
         );
  DFFSX1 Q2_addr_reg_1__3_ ( .D(n5455), .CK(clk), .SN(rst_n), .QN(Q2_addr[11])
         );
  DFFSX1 Q2_addr_reg_0__3_ ( .D(n5454), .CK(clk), .SN(rst_n), .QN(Q2_addr[3])
         );
  DFFSX1 Q2_addr_reg_4__5_ ( .D(n5453), .CK(clk), .SN(rst_n), .QN(Q2_addr[37])
         );
  DFFSX1 Q2_addr_reg_3__5_ ( .D(n5452), .CK(clk), .SN(rst_n), .QN(Q2_addr[29])
         );
  DFFSX1 Q2_addr_reg_2__5_ ( .D(n5451), .CK(clk), .SN(rst_n), .QN(Q2_addr[21])
         );
  DFFSX1 Q2_addr_reg_1__5_ ( .D(n5450), .CK(clk), .SN(rst_n), .QN(Q2_addr[13])
         );
  DFFSX1 Q2_addr_reg_0__5_ ( .D(n5449), .CK(clk), .SN(rst_n), .QN(Q2_addr[5])
         );
  DFFSX1 Q0_addr_reg_2__0_ ( .D(n5448), .CK(clk), .SN(rst_n), .QN(Q0_addr[16])
         );
  DFFSX1 Q0_addr_reg_1__0_ ( .D(n5447), .CK(clk), .SN(rst_n), .QN(Q0_addr[8])
         );
  DFFSX1 Q0_addr_reg_0__0_ ( .D(n5446), .CK(clk), .SN(rst_n), .QN(Q0_addr[0])
         );
  DFFSX1 Q0_addr_reg_2__1_ ( .D(n5445), .CK(clk), .SN(rst_n), .QN(Q0_addr[17])
         );
  DFFSX1 Q0_addr_reg_1__1_ ( .D(n5444), .CK(clk), .SN(rst_n), .QN(Q0_addr[9])
         );
  DFFSX1 Q0_addr_reg_0__1_ ( .D(n5443), .CK(clk), .SN(rst_n), .QN(Q0_addr[1])
         );
  DFFSX1 Q0_addr_reg_2__2_ ( .D(n5442), .CK(clk), .SN(rst_n), .QN(Q0_addr[18])
         );
  DFFSX1 Q0_addr_reg_1__2_ ( .D(n5441), .CK(clk), .SN(rst_n), .QN(Q0_addr[10])
         );
  DFFSX1 Q0_addr_reg_0__2_ ( .D(n5440), .CK(clk), .SN(rst_n), .QN(Q0_addr[2])
         );
  DFFSX1 Q0_addr_reg_2__3_ ( .D(n5439), .CK(clk), .SN(rst_n), .QN(Q0_addr[19])
         );
  DFFSX1 Q0_addr_reg_1__3_ ( .D(n5438), .CK(clk), .SN(rst_n), .QN(Q0_addr[11])
         );
  DFFSX1 Q0_addr_reg_0__3_ ( .D(n5437), .CK(clk), .SN(rst_n), .QN(Q0_addr[3])
         );
  DFFSX1 ram_sel_reg_reg_4__0_ ( .D(n5436), .CK(clk), .SN(rst_n), .Q(n28759), 
        .QN(ram_sel_reg[8]) );
  DFFSX1 ram_sel_reg_reg_3__0_ ( .D(n5435), .CK(clk), .SN(rst_n), .QN(
        ram_sel_reg[6]) );
  DFFSX1 ram_sel_reg_reg_2__0_ ( .D(n5434), .CK(clk), .SN(rst_n), .QN(
        ram_sel_reg[4]) );
  DFFSX1 ram_sel_reg_reg_1__0_ ( .D(n5433), .CK(clk), .SN(rst_n), .QN(
        ram_sel_reg[2]) );
  DFFSX1 ram_sel_reg_reg_0__0_ ( .D(n5432), .CK(clk), .SN(rst_n), .QN(
        ram_sel_reg[0]) );
  DFFSX1 ram_sel_reg_reg_4__1_ ( .D(n5431), .CK(clk), .SN(rst_n), .QN(
        ram_sel_reg[9]) );
  DFFSX1 ram_sel_reg_reg_3__1_ ( .D(n5430), .CK(clk), .SN(rst_n), .QN(
        ram_sel_reg[7]) );
  DFFSX1 ram_sel_reg_reg_2__1_ ( .D(n5429), .CK(clk), .SN(rst_n), .QN(
        ram_sel_reg[5]) );
  DFFSX1 ram_sel_reg_reg_1__1_ ( .D(n5428), .CK(clk), .SN(rst_n), .QN(
        ram_sel_reg[3]) );
  DFFSX1 ram_sel_reg_reg_0__1_ ( .D(n5427), .CK(clk), .SN(rst_n), .QN(
        ram_sel_reg[1]) );
  DFFSX1 D_sel_reg_reg_4__0_ ( .D(n5426), .CK(clk), .SN(rst_n), .Q(n28678), 
        .QN(D_sel_reg_4__0_) );
  DFFSX1 B_sel_reg_reg_3__0_ ( .D(n5425), .CK(clk), .SN(rst_n), .QN(
        B_sel_reg[3]) );
  DFFSX1 B_sel_reg_reg_2__0_ ( .D(n5424), .CK(clk), .SN(rst_n), .QN(
        B_sel_reg[2]) );
  DFFSX1 B_sel_reg_reg_1__0_ ( .D(n5423), .CK(clk), .SN(rst_n), .QN(
        B_sel_reg[1]) );
  DFFSX1 B_sel_reg_reg_0__0_ ( .D(n5422), .CK(clk), .SN(rst_n), .Q(n28675), 
        .QN(B_sel_reg[0]) );
  DFFSX1 A_sel_reg_reg_4__1_ ( .D(n5421), .CK(clk), .SN(rst_n), .Q(n28672), 
        .QN(A_sel_reg[4]) );
  DFFSX1 A_sel_reg_reg_3__1_ ( .D(n5420), .CK(clk), .SN(rst_n), .QN(
        A_sel_reg[3]) );
  DFFSX1 A_sel_reg_reg_2__1_ ( .D(n5419), .CK(clk), .SN(rst_n), .QN(
        A_sel_reg[2]) );
  DFFSX1 A_sel_reg_reg_1__1_ ( .D(n5418), .CK(clk), .SN(rst_n), .QN(
        A_sel_reg[1]) );
  DFFSX1 A_sel_reg_reg_0__1_ ( .D(n5417), .CK(clk), .SN(rst_n), .QN(
        A_sel_reg[0]) );
  DFFSX1 C_sel_reg_reg_4__0_ ( .D(n5416), .CK(clk), .SN(rst_n), .Q(n28677), 
        .QN(C_sel_reg[8]) );
  DFFSX1 C_sel_reg_reg_3__0_ ( .D(n5415), .CK(clk), .SN(rst_n), .QN(
        C_sel_reg[6]) );
  DFFSX1 C_sel_reg_reg_2__0_ ( .D(n5414), .CK(clk), .SN(rst_n), .QN(
        C_sel_reg[4]) );
  DFFSX1 C_sel_reg_reg_1__0_ ( .D(n5413), .CK(clk), .SN(rst_n), .QN(
        C_sel_reg[2]) );
  DFFSX1 C_sel_reg_reg_4__1_ ( .D(n5411), .CK(clk), .SN(rst_n), .Q(n28671), 
        .QN(C_sel_reg[9]) );
  DFFSX1 C_sel_reg_reg_3__1_ ( .D(n5410), .CK(clk), .SN(rst_n), .QN(
        C_sel_reg[7]) );
  DFFSX1 C_sel_reg_reg_2__1_ ( .D(n5409), .CK(clk), .SN(rst_n), .QN(
        C_sel_reg[5]) );
  DFFSX1 C_sel_reg_reg_1__1_ ( .D(n5408), .CK(clk), .SN(rst_n), .QN(
        C_sel_reg[3]) );
  DFFSX1 C_sel_reg_reg_0__1_ ( .D(n5407), .CK(clk), .SN(rst_n), .QN(
        C_sel_reg[1]) );
  DFFSX1 T1_factor_reg ( .D(n5696), .CK(clk), .SN(rst_n), .Q(n29089) );
  DFFSX4 U2_factor_reg_reg ( .D(n29089), .CK(clk), .SN(rst_n), .Q(n29106), 
        .QN(U2_factor_reg) );
  DFFSX1 Q3_addr_reg_4__6_ ( .D(n5404), .CK(clk), .SN(rst_n), .QN(Q3_addr[38])
         );
  DFFSX1 Q3_addr_reg_3__6_ ( .D(n5403), .CK(clk), .SN(rst_n), .QN(Q3_addr[30])
         );
  DFFSX1 Q3_addr_reg_2__6_ ( .D(n5402), .CK(clk), .SN(rst_n), .QN(Q3_addr[22])
         );
  DFFSX1 Q3_addr_reg_1__6_ ( .D(n5401), .CK(clk), .SN(rst_n), .QN(Q3_addr[14])
         );
  DFFSX1 Q3_addr_reg_0__6_ ( .D(n5400), .CK(clk), .SN(rst_n), .QN(Q3_addr[6])
         );
  DFFSX1 Q1_addr_reg_4__6_ ( .D(n5399), .CK(clk), .SN(rst_n), .QN(Q1_addr[38])
         );
  DFFSX1 Q1_addr_reg_3__6_ ( .D(n5398), .CK(clk), .SN(rst_n), .QN(Q1_addr[30])
         );
  DFFSX1 Q1_addr_reg_2__6_ ( .D(n5397), .CK(clk), .SN(rst_n), .QN(Q1_addr[22])
         );
  DFFSX1 Q1_addr_reg_1__6_ ( .D(n5396), .CK(clk), .SN(rst_n), .QN(Q1_addr[14])
         );
  DFFSX1 Q1_addr_reg_0__6_ ( .D(n5395), .CK(clk), .SN(rst_n), .Q(n28919), .QN(
        Q1_addr[6]) );
  DFFSX1 Q1_addr_reg_4__7_ ( .D(n5394), .CK(clk), .SN(rst_n), .QN(Q1_addr[39])
         );
  DFFSX1 Q1_addr_reg_3__7_ ( .D(n5393), .CK(clk), .SN(rst_n), .QN(Q1_addr[31])
         );
  DFFSX1 Q1_addr_reg_2__7_ ( .D(n5392), .CK(clk), .SN(rst_n), .QN(Q1_addr[23])
         );
  DFFSX1 Q1_addr_reg_1__7_ ( .D(n5391), .CK(clk), .SN(rst_n), .QN(Q1_addr[15])
         );
  DFFSX1 Q1_addr_reg_0__7_ ( .D(n5390), .CK(clk), .SN(rst_n), .Q(n28920), .QN(
        Q1_addr[7]) );
  DFFSX1 Q0_addr_reg_4__7_ ( .D(n5389), .CK(clk), .SN(rst_n), .QN(Q0_addr[39])
         );
  DFFSX1 Q0_addr_reg_3__7_ ( .D(n5388), .CK(clk), .SN(rst_n), .QN(Q0_addr[31])
         );
  DFFSX1 Q0_addr_reg_2__7_ ( .D(n5387), .CK(clk), .SN(rst_n), .QN(Q0_addr[23])
         );
  DFFSX1 Q0_addr_reg_1__7_ ( .D(n5386), .CK(clk), .SN(rst_n), .QN(Q0_addr[15])
         );
  DFFSX1 Q0_addr_reg_0__7_ ( .D(n5385), .CK(clk), .SN(rst_n), .QN(Q0_addr[7])
         );
  DFFSX1 Q1_addr_reg_4__5_ ( .D(n5384), .CK(clk), .SN(rst_n), .QN(Q1_addr[37])
         );
  DFFSX1 Q1_addr_reg_3__5_ ( .D(n5383), .CK(clk), .SN(rst_n), .QN(Q1_addr[29])
         );
  DFFSX1 Q1_addr_reg_2__5_ ( .D(n5382), .CK(clk), .SN(rst_n), .QN(Q1_addr[21])
         );
  DFFSX1 Q1_addr_reg_1__5_ ( .D(n5381), .CK(clk), .SN(rst_n), .QN(Q1_addr[13])
         );
  DFFSX1 Q1_addr_reg_0__5_ ( .D(n5380), .CK(clk), .SN(rst_n), .Q(n28757), .QN(
        Q1_addr[5]) );
  DFFSX1 Q0_addr_reg_4__5_ ( .D(n5379), .CK(clk), .SN(rst_n), .QN(Q0_addr[37])
         );
  DFFSX1 Q0_addr_reg_3__5_ ( .D(n5378), .CK(clk), .SN(rst_n), .QN(Q0_addr[29])
         );
  DFFSX1 Q0_addr_reg_2__5_ ( .D(n5377), .CK(clk), .SN(rst_n), .QN(Q0_addr[21])
         );
  DFFSX1 Q0_addr_reg_1__5_ ( .D(n5376), .CK(clk), .SN(rst_n), .QN(Q0_addr[13])
         );
  DFFSX1 Q0_addr_reg_0__5_ ( .D(n5375), .CK(clk), .SN(rst_n), .QN(Q0_addr[5])
         );
  DFFSX1 Q0_addr_reg_4__4_ ( .D(n5374), .CK(clk), .SN(rst_n), .QN(Q0_addr[36])
         );
  DFFSX1 Q0_addr_reg_3__4_ ( .D(n5373), .CK(clk), .SN(rst_n), .QN(Q0_addr[28])
         );
  DFFSX1 Q0_addr_reg_2__4_ ( .D(n5372), .CK(clk), .SN(rst_n), .QN(Q0_addr[20])
         );
  DFFSX1 Q0_addr_reg_1__4_ ( .D(n5371), .CK(clk), .SN(rst_n), .QN(Q0_addr[12])
         );
  DFFSX1 Q0_addr_reg_0__4_ ( .D(n5370), .CK(clk), .SN(rst_n), .QN(Q0_addr[4])
         );
  DFFSX1 Q2_addr_reg_4__4_ ( .D(n5369), .CK(clk), .SN(rst_n), .QN(Q2_addr[36])
         );
  DFFSX1 Q2_addr_reg_3__4_ ( .D(n5368), .CK(clk), .SN(rst_n), .QN(Q2_addr[28])
         );
  DFFSX1 Q2_addr_reg_2__4_ ( .D(n5367), .CK(clk), .SN(rst_n), .QN(Q2_addr[20])
         );
  DFFSX1 Q2_addr_reg_1__4_ ( .D(n5366), .CK(clk), .SN(rst_n), .QN(Q2_addr[12])
         );
  DFFSX1 Q2_addr_reg_0__4_ ( .D(n5365), .CK(clk), .SN(rst_n), .QN(Q2_addr[4])
         );
  DFFSX1 Q0_addr_reg_4__6_ ( .D(n5364), .CK(clk), .SN(rst_n), .QN(Q0_addr[38])
         );
  DFFSX1 Q0_addr_reg_3__6_ ( .D(n5363), .CK(clk), .SN(rst_n), .QN(Q0_addr[30])
         );
  DFFSX1 Q0_addr_reg_2__6_ ( .D(n5362), .CK(clk), .SN(rst_n), .QN(Q0_addr[22])
         );
  DFFSX1 Q0_addr_reg_1__6_ ( .D(n5361), .CK(clk), .SN(rst_n), .QN(Q0_addr[14])
         );
  DFFSX1 Q0_addr_reg_0__6_ ( .D(n5360), .CK(clk), .SN(rst_n), .QN(Q0_addr[6])
         );
  DFFSX1 Q2_addr_reg_4__6_ ( .D(n5359), .CK(clk), .SN(rst_n), .QN(Q2_addr[38])
         );
  DFFSX1 Q2_addr_reg_3__6_ ( .D(n5358), .CK(clk), .SN(rst_n), .QN(Q2_addr[30])
         );
  DFFSX1 Q2_addr_reg_2__6_ ( .D(n5357), .CK(clk), .SN(rst_n), .QN(Q2_addr[22])
         );
  DFFSX1 Q2_addr_reg_1__6_ ( .D(n5356), .CK(clk), .SN(rst_n), .QN(Q2_addr[14])
         );
  DFFSX1 Q2_addr_reg_0__6_ ( .D(n5355), .CK(clk), .SN(rst_n), .QN(Q2_addr[6])
         );
  DFFSX1 Q3_addr_reg_4__7_ ( .D(n5354), .CK(clk), .SN(rst_n), .QN(Q3_addr[39])
         );
  DFFSX1 Q3_addr_reg_3__7_ ( .D(n5353), .CK(clk), .SN(rst_n), .QN(Q3_addr[31])
         );
  DFFSX1 Q3_addr_reg_2__7_ ( .D(n5352), .CK(clk), .SN(rst_n), .QN(Q3_addr[23])
         );
  DFFSX1 Q3_addr_reg_1__7_ ( .D(n5351), .CK(clk), .SN(rst_n), .QN(Q3_addr[15])
         );
  DFFSX1 Q3_addr_reg_0__7_ ( .D(n5350), .CK(clk), .SN(rst_n), .QN(Q3_addr[7])
         );
  DFFSX1 Q2_addr_reg_4__7_ ( .D(n5349), .CK(clk), .SN(rst_n), .QN(Q2_addr[39])
         );
  DFFSX1 Q2_addr_reg_3__7_ ( .D(n5348), .CK(clk), .SN(rst_n), .QN(Q2_addr[31])
         );
  DFFSX1 Q2_addr_reg_2__7_ ( .D(n5347), .CK(clk), .SN(rst_n), .QN(Q2_addr[23])
         );
  DFFSX1 Q2_addr_reg_1__7_ ( .D(n5346), .CK(clk), .SN(rst_n), .QN(Q2_addr[15])
         );
  DFFSX1 Q2_addr_reg_0__7_ ( .D(n5345), .CK(clk), .SN(rst_n), .QN(Q2_addr[7])
         );
  DFFSX1 U1_A_i_d0_reg_9_ ( .D(n29036), .CK(clk), .SN(rst_n), .QN(U1_A_i_d0[9]) );
  DFFSX1 U1_A_i_d0_reg_8_ ( .D(n29035), .CK(clk), .SN(rst_n), .QN(U1_A_i_d0[8]) );
  DFFSX1 U1_A_i_d0_reg_7_ ( .D(n29034), .CK(clk), .SN(rst_n), .QN(U1_A_i_d0[7]) );
  DFFSX1 U1_A_i_d0_reg_6_ ( .D(n29033), .CK(clk), .SN(rst_n), .Q(n7068), .QN(
        U1_A_i_d0[6]) );
  DFFSX1 U1_A_i_d0_reg_5_ ( .D(n29017), .CK(clk), .SN(rst_n), .QN(U1_A_i_d0[5]) );
  DFFSX1 U1_A_r_d0_reg_25_ ( .D(n28749), .CK(clk), .SN(rst_n), .Q(n29007), 
        .QN(U1_A_r_d0[25]) );
  DFFSX1 U1_A_r_d0_reg_24_ ( .D(n28687), .CK(clk), .SN(rst_n), .QN(
        U1_A_r_d0[24]) );
  DFFSX1 U1_A_i_d0_reg_4_ ( .D(n29011), .CK(clk), .SN(rst_n), .QN(U1_A_i_d0[4]) );
  DFFSX1 U1_A_r_d0_reg_23_ ( .D(n28684), .CK(clk), .SN(rst_n), .Q(n7074), .QN(
        U1_A_r_d0[23]) );
  DFFSX1 U1_A_r_d0_reg_22_ ( .D(n28710), .CK(clk), .SN(rst_n), .QN(
        U1_A_r_d0[22]) );
  DFFSX1 U1_A_r_d0_reg_21_ ( .D(n28685), .CK(clk), .SN(rst_n), .QN(
        U1_A_r_d0[21]) );
  DFFSX1 U1_A_r_d0_reg_20_ ( .D(n28708), .CK(clk), .SN(rst_n), .Q(n7082), .QN(
        U1_A_r_d0[20]) );
  DFFSX1 U1_A_r_d0_reg_19_ ( .D(n28686), .CK(clk), .SN(rst_n), .Q(n5760), .QN(
        U1_A_r_d0[19]) );
  DFFSX1 U1_A_r_d0_reg_18_ ( .D(n28711), .CK(clk), .SN(rst_n), .Q(n7071), .QN(
        U1_A_r_d0[18]) );
  DFFSX1 U1_A_r_d0_reg_17_ ( .D(n28688), .CK(clk), .SN(rst_n), .QN(
        U1_A_r_d0[17]) );
  DFFSX1 U1_A_r_d0_reg_16_ ( .D(n28712), .CK(clk), .SN(rst_n), .Q(n7070), .QN(
        U1_A_r_d0[16]) );
  DFFSX1 U1_A_r_d0_reg_15_ ( .D(n28746), .CK(clk), .SN(rst_n), .QN(
        U1_A_r_d0[15]) );
  DFFSX1 U1_A_r_d0_reg_14_ ( .D(n28683), .CK(clk), .SN(rst_n), .QN(
        U1_A_r_d0[14]) );
  DFFSX1 U1_A_i_d0_reg_3_ ( .D(n29032), .CK(clk), .SN(rst_n), .QN(U1_A_i_d0[3]) );
  DFFSX1 U1_A_r_d0_reg_13_ ( .D(n28681), .CK(clk), .SN(rst_n), .QN(
        U1_A_r_d0[13]) );
  DFFSX1 U1_A_r_d0_reg_12_ ( .D(n28713), .CK(clk), .SN(rst_n), .QN(
        U1_A_r_d0[12]) );
  DFFSX1 U1_A_r_d0_reg_11_ ( .D(n28747), .CK(clk), .SN(rst_n), .QN(
        U1_A_r_d0[11]) );
  DFFSX1 U1_A_r_d0_reg_10_ ( .D(n28748), .CK(clk), .SN(rst_n), .Q(n7065), .QN(
        U1_A_r_d0[10]) );
  DFFSX1 U1_A_r_d0_reg_9_ ( .D(n6932), .CK(clk), .SN(rst_n), .QN(U1_A_r_d0[9])
         );
  DFFSX1 U1_A_r_d0_reg_8_ ( .D(n6910), .CK(clk), .SN(rst_n), .QN(U1_A_r_d0[8])
         );
  DFFSX1 U1_A_r_d0_reg_7_ ( .D(n29100), .CK(clk), .SN(rst_n), .QN(U1_A_r_d0[7]) );
  DFFSX1 U1_A_r_d0_reg_6_ ( .D(n28750), .CK(clk), .SN(rst_n), .Q(n7063), .QN(
        U1_A_r_d0[6]) );
  DFFSX1 U1_A_r_d0_reg_5_ ( .D(n29105), .CK(clk), .SN(rst_n), .QN(U1_A_r_d0[5]) );
  DFFSX1 U1_A_r_d0_reg_4_ ( .D(n29104), .CK(clk), .SN(rst_n), .QN(U1_A_r_d0[4]) );
  DFFSX1 U1_A_i_d0_reg_2_ ( .D(n29016), .CK(clk), .SN(rst_n), .QN(U1_A_i_d0[2]) );
  DFFSX1 U1_A_r_d0_reg_3_ ( .D(n29103), .CK(clk), .SN(rst_n), .QN(U1_A_r_d0[3]) );
  DFFSX1 U1_A_r_d0_reg_2_ ( .D(n29102), .CK(clk), .SN(rst_n), .QN(U1_A_r_d0[2]) );
  DFFSX1 U1_A_r_d0_reg_0_ ( .D(n28751), .CK(clk), .SN(rst_n), .QN(U1_A_r_d0[0]) );
  DFFSX1 U1_A_i_d0_reg_25_ ( .D(n29031), .CK(clk), .SN(rst_n), .Q(n29008), 
        .QN(U1_A_i_d0[25]) );
  DFFSX1 U1_A_i_d0_reg_24_ ( .D(n29030), .CK(clk), .SN(rst_n), .Q(n7076), .QN(
        U1_A_i_d0[24]) );
  DFFSX1 U1_A_i_d0_reg_23_ ( .D(n29029), .CK(clk), .SN(rst_n), .Q(n8156), .QN(
        U1_A_i_d0[23]) );
  DFFSX1 U1_A_i_d0_reg_22_ ( .D(n29028), .CK(clk), .SN(rst_n), .Q(n5757), .QN(
        U1_A_i_d0[22]) );
  DFFSX1 U1_A_i_d0_reg_21_ ( .D(n29027), .CK(clk), .SN(rst_n), .Q(n7072), .QN(
        U1_A_i_d0[21]) );
  DFFSX1 U1_A_i_d0_reg_20_ ( .D(n29026), .CK(clk), .SN(rst_n), .Q(n7081), .QN(
        U1_A_i_d0[20]) );
  DFFSX1 U1_A_i_d0_reg_1_ ( .D(n29013), .CK(clk), .SN(rst_n), .QN(U1_A_i_d0[1]) );
  DFFSX1 U1_A_i_d0_reg_19_ ( .D(n29025), .CK(clk), .SN(rst_n), .Q(n5782), .QN(
        U1_A_i_d0[19]) );
  DFFSX1 U1_A_i_d0_reg_18_ ( .D(n29024), .CK(clk), .SN(rst_n), .Q(n8173), .QN(
        U1_A_i_d0[18]) );
  DFFSX1 U1_A_i_d0_reg_17_ ( .D(n29023), .CK(clk), .SN(rst_n), .Q(n5783), .QN(
        U1_A_i_d0[17]) );
  DFFSX1 U1_A_i_d0_reg_16_ ( .D(n29022), .CK(clk), .SN(rst_n), .Q(n7069), .QN(
        U1_A_i_d0[16]) );
  DFFSX1 U1_A_i_d0_reg_15_ ( .D(n29015), .CK(clk), .SN(rst_n), .Q(n7077), .QN(
        U1_A_i_d0[15]) );
  DFFSX1 U1_A_i_d0_reg_14_ ( .D(n29021), .CK(clk), .SN(rst_n), .Q(n7073), .QN(
        U1_A_i_d0[14]) );
  DFFSX1 U1_A_i_d0_reg_13_ ( .D(n29014), .CK(clk), .SN(rst_n), .QN(
        U1_A_i_d0[13]) );
  DFFSX1 U1_A_i_d0_reg_12_ ( .D(n29020), .CK(clk), .SN(rst_n), .Q(n5787), .QN(
        U1_A_i_d0[12]) );
  DFFSX1 U1_A_i_d0_reg_11_ ( .D(n29019), .CK(clk), .SN(rst_n), .QN(
        U1_A_i_d0[11]) );
  DFFSX1 U1_A_i_d0_reg_10_ ( .D(n29018), .CK(clk), .SN(rst_n), .Q(n7064), .QN(
        U1_A_i_d0[10]) );
  DFFSX1 U1_A_i_d0_reg_0_ ( .D(n28676), .CK(clk), .SN(rst_n), .QN(U1_A_i_d0[0]) );
  DFFSX1 U2_A_i_d_reg_9_ ( .D(n29088), .CK(clk), .SN(rst_n), .QN(U2_A_i_d[9])
         );
  DFFSX1 DATA0_reg_9_ ( .D(n5291), .CK(clk), .SN(rst_n), .QN(DATA0[9]) );
  DFFSX1 U2_A_i_d_reg_8_ ( .D(n29087), .CK(clk), .SN(rst_n), .QN(U2_A_i_d[8])
         );
  DFFSX1 DATA0_reg_8_ ( .D(n5289), .CK(clk), .SN(rst_n), .QN(DATA0[8]) );
  DFFSX1 U2_A_i_d_reg_7_ ( .D(n29086), .CK(clk), .SN(rst_n), .QN(U2_A_i_d[7])
         );
  DFFSX1 DATA0_reg_7_ ( .D(n5287), .CK(clk), .SN(rst_n), .QN(DATA0[7]) );
  DFFSX1 U2_A_i_d_reg_6_ ( .D(n29085), .CK(clk), .SN(rst_n), .Q(n5773), .QN(
        U2_A_i_d[6]) );
  DFFSX1 DATA0_reg_6_ ( .D(n5285), .CK(clk), .SN(rst_n), .QN(DATA0[6]) );
  DFFSX1 U2_A_i_d_reg_5_ ( .D(n29084), .CK(clk), .SN(rst_n), .QN(U2_A_i_d[5])
         );
  DFFSX1 DATA0_reg_5_ ( .D(n5283), .CK(clk), .SN(rst_n), .QN(DATA0[5]) );
  DFFSX1 U2_A_r_d_reg_25_ ( .D(n29083), .CK(clk), .SN(rst_n), .Q(n29010), .QN(
        U2_A_r_d[25]) );
  DFFSX1 DATA0_reg_51_ ( .D(n5281), .CK(clk), .SN(rst_n), .QN(DATA0[51]) );
  DFFSX1 U2_A_r_d_reg_24_ ( .D(n29082), .CK(clk), .SN(rst_n), .QN(U2_A_r_d[24]) );
  DFFSX1 DATA0_reg_50_ ( .D(n5279), .CK(clk), .SN(rst_n), .QN(DATA0[50]) );
  DFFSX1 U2_A_i_d_reg_4_ ( .D(n29081), .CK(clk), .SN(rst_n), .QN(U2_A_i_d[4])
         );
  DFFSX1 DATA0_reg_4_ ( .D(n5277), .CK(clk), .SN(rst_n), .QN(DATA0[4]) );
  DFFSX1 U2_A_r_d_reg_23_ ( .D(n29080), .CK(clk), .SN(rst_n), .QN(U2_A_r_d[23]) );
  DFFSX1 DATA0_reg_49_ ( .D(n5275), .CK(clk), .SN(rst_n), .QN(DATA0[49]) );
  DFFSX1 U2_A_r_d_reg_22_ ( .D(n29079), .CK(clk), .SN(rst_n), .QN(U2_A_r_d[22]) );
  DFFSX1 DATA0_reg_48_ ( .D(n5273), .CK(clk), .SN(rst_n), .QN(DATA0[48]) );
  DFFSX1 U2_A_r_d_reg_21_ ( .D(n29078), .CK(clk), .SN(rst_n), .Q(n7075), .QN(
        U2_A_r_d[21]) );
  DFFSX1 DATA0_reg_47_ ( .D(n5271), .CK(clk), .SN(rst_n), .QN(DATA0[47]) );
  DFFSX1 U2_A_r_d_reg_20_ ( .D(n29077), .CK(clk), .SN(rst_n), .Q(n8077), .QN(
        U2_A_r_d[20]) );
  DFFSX1 DATA0_reg_46_ ( .D(n5269), .CK(clk), .SN(rst_n), .QN(DATA0[46]) );
  DFFSX1 U2_A_r_d_reg_19_ ( .D(n29076), .CK(clk), .SN(rst_n), .QN(U2_A_r_d[19]) );
  DFFSX1 DATA0_reg_45_ ( .D(n5267), .CK(clk), .SN(rst_n), .QN(DATA0[45]) );
  DFFSX1 U2_A_r_d_reg_18_ ( .D(n29075), .CK(clk), .SN(rst_n), .QN(U2_A_r_d[18]) );
  DFFSX1 DATA0_reg_44_ ( .D(n5265), .CK(clk), .SN(rst_n), .QN(DATA0[44]) );
  DFFSX1 U2_A_r_d_reg_17_ ( .D(n29074), .CK(clk), .SN(rst_n), .QN(U2_A_r_d[17]) );
  DFFSX1 DATA0_reg_43_ ( .D(n5263), .CK(clk), .SN(rst_n), .QN(DATA0[43]) );
  DFFSX1 U2_A_r_d_reg_16_ ( .D(n29073), .CK(clk), .SN(rst_n), .QN(U2_A_r_d[16]) );
  DFFSX1 DATA0_reg_42_ ( .D(n5261), .CK(clk), .SN(rst_n), .QN(DATA0[42]) );
  DFFSX1 U2_A_r_d_reg_15_ ( .D(n29072), .CK(clk), .SN(rst_n), .QN(U2_A_r_d[15]) );
  DFFSX1 DATA0_reg_41_ ( .D(n5259), .CK(clk), .SN(rst_n), .QN(DATA0[41]) );
  DFFSX1 U2_A_r_d_reg_14_ ( .D(n29071), .CK(clk), .SN(rst_n), .QN(U2_A_r_d[14]) );
  DFFSX1 DATA0_reg_40_ ( .D(n5257), .CK(clk), .SN(rst_n), .QN(DATA0[40]) );
  DFFSX1 U2_A_i_d_reg_3_ ( .D(n29070), .CK(clk), .SN(rst_n), .QN(U2_A_i_d[3])
         );
  DFFSX1 DATA0_reg_3_ ( .D(n5255), .CK(clk), .SN(rst_n), .QN(DATA0[3]) );
  DFFSX1 U2_A_r_d_reg_13_ ( .D(n29069), .CK(clk), .SN(rst_n), .QN(U2_A_r_d[13]) );
  DFFSX1 DATA0_reg_39_ ( .D(n5253), .CK(clk), .SN(rst_n), .QN(DATA0[39]) );
  DFFSX1 U2_A_r_d_reg_12_ ( .D(n29068), .CK(clk), .SN(rst_n), .QN(U2_A_r_d[12]) );
  DFFSX1 DATA0_reg_38_ ( .D(n5251), .CK(clk), .SN(rst_n), .QN(DATA0[38]) );
  DFFSX1 U2_A_r_d_reg_11_ ( .D(n29067), .CK(clk), .SN(rst_n), .QN(U2_A_r_d[11]) );
  DFFSX1 DATA0_reg_37_ ( .D(n5249), .CK(clk), .SN(rst_n), .QN(DATA0[37]) );
  DFFSX1 U2_A_r_d_reg_10_ ( .D(n29066), .CK(clk), .SN(rst_n), .QN(U2_A_r_d[10]) );
  DFFSX1 DATA0_reg_36_ ( .D(n5247), .CK(clk), .SN(rst_n), .QN(DATA0[36]) );
  DFFSX1 U2_A_r_d_reg_9_ ( .D(n29065), .CK(clk), .SN(rst_n), .QN(U2_A_r_d[9])
         );
  DFFSX1 DATA0_reg_35_ ( .D(n5245), .CK(clk), .SN(rst_n), .QN(DATA0[35]) );
  DFFSX1 U2_A_r_d_reg_8_ ( .D(n29064), .CK(clk), .SN(rst_n), .QN(U2_A_r_d[8])
         );
  DFFSX1 DATA0_reg_34_ ( .D(n5243), .CK(clk), .SN(rst_n), .QN(DATA0[34]) );
  DFFSX1 U2_A_r_d_reg_7_ ( .D(n29063), .CK(clk), .SN(rst_n), .QN(U2_A_r_d[7])
         );
  DFFSX1 DATA0_reg_33_ ( .D(n5241), .CK(clk), .SN(rst_n), .QN(DATA0[33]) );
  DFFSX1 U2_A_r_d_reg_6_ ( .D(n29062), .CK(clk), .SN(rst_n), .Q(n5776), .QN(
        U2_A_r_d[6]) );
  DFFSX1 DATA0_reg_32_ ( .D(n5239), .CK(clk), .SN(rst_n), .QN(DATA0[32]) );
  DFFSX1 U2_A_r_d_reg_5_ ( .D(n29061), .CK(clk), .SN(rst_n), .QN(U2_A_r_d[5])
         );
  DFFSX1 DATA0_reg_31_ ( .D(n5237), .CK(clk), .SN(rst_n), .QN(DATA0[31]) );
  DFFSX1 U2_A_r_d_reg_4_ ( .D(n29060), .CK(clk), .SN(rst_n), .Q(n7067), .QN(
        U2_A_r_d[4]) );
  DFFSX1 DATA0_reg_30_ ( .D(n5235), .CK(clk), .SN(rst_n), .QN(DATA0[30]) );
  DFFSX1 U2_A_i_d_reg_2_ ( .D(n29059), .CK(clk), .SN(rst_n), .QN(U2_A_i_d[2])
         );
  DFFSX1 DATA0_reg_2_ ( .D(n5233), .CK(clk), .SN(rst_n), .QN(DATA0[2]) );
  DFFSX1 U2_A_r_d_reg_3_ ( .D(n29058), .CK(clk), .SN(rst_n), .QN(U2_A_r_d[3])
         );
  DFFSX1 DATA0_reg_29_ ( .D(n5231), .CK(clk), .SN(rst_n), .QN(DATA0[29]) );
  DFFSX1 U2_A_r_d_reg_2_ ( .D(n29057), .CK(clk), .SN(rst_n), .QN(U2_A_r_d[2])
         );
  DFFSX1 DATA0_reg_28_ ( .D(n5229), .CK(clk), .SN(rst_n), .QN(DATA0[28]) );
  DFFSX1 U2_A_r_d_reg_1_ ( .D(n29056), .CK(clk), .SN(rst_n), .QN(U2_A_r_d[1])
         );
  DFFSX1 DATA0_reg_27_ ( .D(n5227), .CK(clk), .SN(rst_n), .QN(DATA0[27]) );
  DFFSX1 U2_A_r_d_reg_0_ ( .D(n29055), .CK(clk), .SN(rst_n), .QN(U2_A_r_d[0])
         );
  DFFSX1 DATA0_reg_26_ ( .D(n5225), .CK(clk), .SN(rst_n), .QN(DATA0[26]) );
  DFFSX1 U2_A_i_d_reg_25_ ( .D(n29054), .CK(clk), .SN(rst_n), .Q(n29009), .QN(
        U2_A_i_d[25]) );
  DFFSX1 DATA0_reg_25_ ( .D(n5223), .CK(clk), .SN(rst_n), .QN(DATA0[25]) );
  DFFSX1 U2_A_i_d_reg_24_ ( .D(n29053), .CK(clk), .SN(rst_n), .QN(U2_A_i_d[24]) );
  DFFSX1 DATA0_reg_24_ ( .D(n5221), .CK(clk), .SN(rst_n), .QN(DATA0[24]) );
  DFFSX1 U2_A_i_d_reg_23_ ( .D(n29052), .CK(clk), .SN(rst_n), .QN(U2_A_i_d[23]) );
  DFFSX1 DATA0_reg_23_ ( .D(n5219), .CK(clk), .SN(rst_n), .QN(DATA0[23]) );
  DFFSX1 U2_A_i_d_reg_22_ ( .D(n29051), .CK(clk), .SN(rst_n), .QN(U2_A_i_d[22]) );
  DFFSX1 DATA0_reg_22_ ( .D(n5217), .CK(clk), .SN(rst_n), .QN(DATA0[22]) );
  DFFSX1 U2_A_i_d_reg_21_ ( .D(n29050), .CK(clk), .SN(rst_n), .QN(U2_A_i_d[21]) );
  DFFSX1 DATA0_reg_21_ ( .D(n5215), .CK(clk), .SN(rst_n), .QN(DATA0[21]) );
  DFFSX1 U2_A_i_d_reg_20_ ( .D(n29049), .CK(clk), .SN(rst_n), .QN(U2_A_i_d[20]) );
  DFFSX1 DATA0_reg_20_ ( .D(n5213), .CK(clk), .SN(rst_n), .QN(DATA0[20]) );
  DFFSX1 U2_A_i_d_reg_1_ ( .D(n29048), .CK(clk), .SN(rst_n), .QN(U2_A_i_d[1])
         );
  DFFSX1 DATA0_reg_1_ ( .D(n5211), .CK(clk), .SN(rst_n), .QN(DATA0[1]) );
  DFFSX1 U2_A_i_d_reg_19_ ( .D(n29047), .CK(clk), .SN(rst_n), .QN(U2_A_i_d[19]) );
  DFFSX1 DATA0_reg_19_ ( .D(n5209), .CK(clk), .SN(rst_n), .QN(DATA0[19]) );
  DFFSX1 U2_A_i_d_reg_18_ ( .D(n29046), .CK(clk), .SN(rst_n), .Q(n5780), .QN(
        U2_A_i_d[18]) );
  DFFSX1 DATA0_reg_18_ ( .D(n5207), .CK(clk), .SN(rst_n), .QN(DATA0[18]) );
  DFFSX1 U2_A_i_d_reg_17_ ( .D(n29045), .CK(clk), .SN(rst_n), .QN(U2_A_i_d[17]) );
  DFFSX1 DATA0_reg_17_ ( .D(n5205), .CK(clk), .SN(rst_n), .QN(DATA0[17]) );
  DFFSX1 U2_A_i_d_reg_16_ ( .D(n29044), .CK(clk), .SN(rst_n), .Q(n7079), .QN(
        U2_A_i_d[16]) );
  DFFSX1 DATA0_reg_16_ ( .D(n5203), .CK(clk), .SN(rst_n), .QN(DATA0[16]) );
  DFFSX1 U2_A_i_d_reg_15_ ( .D(n29043), .CK(clk), .SN(rst_n), .QN(U2_A_i_d[15]) );
  DFFSX1 DATA0_reg_15_ ( .D(n5201), .CK(clk), .SN(rst_n), .QN(DATA0[15]) );
  DFFSX1 U2_A_i_d_reg_14_ ( .D(n29042), .CK(clk), .SN(rst_n), .Q(n5781), .QN(
        U2_A_i_d[14]) );
  DFFSX1 DATA0_reg_14_ ( .D(n5199), .CK(clk), .SN(rst_n), .QN(DATA0[14]) );
  DFFSX1 U2_A_i_d_reg_13_ ( .D(n29041), .CK(clk), .SN(rst_n), .QN(U2_A_i_d[13]) );
  DFFSX1 DATA0_reg_13_ ( .D(n5197), .CK(clk), .SN(rst_n), .QN(DATA0[13]) );
  DFFSX1 U2_A_i_d_reg_12_ ( .D(n29040), .CK(clk), .SN(rst_n), .Q(n7080), .QN(
        U2_A_i_d[12]) );
  DFFSX1 DATA0_reg_12_ ( .D(n5195), .CK(clk), .SN(rst_n), .QN(DATA0[12]) );
  DFFSX1 U2_A_i_d_reg_11_ ( .D(n29039), .CK(clk), .SN(rst_n), .QN(U2_A_i_d[11]) );
  DFFSX1 DATA0_reg_11_ ( .D(n5193), .CK(clk), .SN(rst_n), .QN(DATA0[11]) );
  DFFSX1 U2_A_i_d_reg_10_ ( .D(n29038), .CK(clk), .SN(rst_n), .QN(U2_A_i_d[10]) );
  DFFSX1 DATA0_reg_10_ ( .D(n5191), .CK(clk), .SN(rst_n), .QN(DATA0[10]) );
  DFFSX1 U2_A_i_d_reg_0_ ( .D(n29037), .CK(clk), .SN(rst_n), .QN(U2_A_i_d[0])
         );
  DFFSX1 DATA0_reg_0_ ( .D(n5189), .CK(clk), .SN(rst_n), .QN(DATA0[0]) );
  DFFSX1 buffer_reg_31_ ( .D(n5188), .CK(clk), .SN(rst_n), .QN(buffer[31]) );
  DFFSX1 buffer_reg_30_ ( .D(n5187), .CK(clk), .SN(rst_n), .QN(buffer[30]) );
  DFFSX1 buffer_reg_29_ ( .D(n5186), .CK(clk), .SN(rst_n), .QN(buffer[29]) );
  DFFSX1 buffer_reg_28_ ( .D(n5185), .CK(clk), .SN(rst_n), .QN(buffer[28]) );
  DFFSX1 buffer_reg_27_ ( .D(n5184), .CK(clk), .SN(rst_n), .QN(buffer[27]) );
  DFFSX1 buffer_reg_26_ ( .D(n5183), .CK(clk), .SN(rst_n), .QN(buffer[26]) );
  DFFSX1 buffer_reg_25_ ( .D(n5182), .CK(clk), .SN(rst_n), .QN(buffer[25]) );
  DFFSX1 buffer_reg_24_ ( .D(n5181), .CK(clk), .SN(rst_n), .QN(buffer[24]) );
  DFFSX1 buffer_reg_23_ ( .D(n5180), .CK(clk), .SN(rst_n), .QN(buffer[23]) );
  DFFSX1 buffer_reg_22_ ( .D(n5179), .CK(clk), .SN(rst_n), .QN(buffer[22]) );
  DFFSX1 buffer_reg_21_ ( .D(n5178), .CK(clk), .SN(rst_n), .QN(buffer[21]) );
  DFFSX1 buffer_reg_20_ ( .D(n5177), .CK(clk), .SN(rst_n), .QN(buffer[20]) );
  DFFSX1 buffer_reg_19_ ( .D(n5176), .CK(clk), .SN(rst_n), .QN(buffer[19]) );
  DFFSX1 buffer_reg_18_ ( .D(n5175), .CK(clk), .SN(rst_n), .QN(buffer[18]) );
  DFFSX1 buffer_reg_17_ ( .D(n5174), .CK(clk), .SN(rst_n), .QN(buffer[17]) );
  DFFSX1 buffer_reg_16_ ( .D(n5173), .CK(clk), .SN(rst_n), .QN(buffer[16]) );
  DFFSX1 buffer_reg_15_ ( .D(n5172), .CK(clk), .SN(rst_n), .QN(buffer[15]) );
  DFFSX1 buffer_reg_14_ ( .D(n5171), .CK(clk), .SN(rst_n), .QN(buffer[14]) );
  DFFSX1 buffer_reg_13_ ( .D(n5170), .CK(clk), .SN(rst_n), .QN(buffer[13]) );
  DFFSX1 buffer_reg_12_ ( .D(n5169), .CK(clk), .SN(rst_n), .QN(buffer[12]) );
  DFFSX1 buffer_reg_11_ ( .D(n5168), .CK(clk), .SN(rst_n), .QN(buffer[11]) );
  DFFSX1 buffer_reg_10_ ( .D(n5167), .CK(clk), .SN(rst_n), .QN(buffer[10]) );
  DFFSX1 buffer_reg_9_ ( .D(n5166), .CK(clk), .SN(rst_n), .QN(buffer[9]) );
  DFFSX1 buffer_reg_8_ ( .D(n5165), .CK(clk), .SN(rst_n), .QN(buffer[8]) );
  DFFSX1 buffer_reg_7_ ( .D(n5164), .CK(clk), .SN(rst_n), .QN(buffer[7]) );
  DFFSX1 buffer_reg_6_ ( .D(n5163), .CK(clk), .SN(rst_n), .QN(buffer[6]) );
  DFFSX1 buffer_reg_5_ ( .D(n5162), .CK(clk), .SN(rst_n), .QN(buffer[5]) );
  DFFSX1 buffer_reg_4_ ( .D(n5161), .CK(clk), .SN(rst_n), .QN(buffer[4]) );
  DFFSX1 buffer_reg_3_ ( .D(n5160), .CK(clk), .SN(rst_n), .QN(buffer[3]) );
  DFFSX1 buffer_reg_2_ ( .D(n5159), .CK(clk), .SN(rst_n), .QN(buffer[2]) );
  DFFSX1 buffer_reg_1_ ( .D(n5158), .CK(clk), .SN(rst_n), .QN(buffer[1]) );
  DFFSX1 buffer_reg_0_ ( .D(n5157), .CK(clk), .SN(rst_n), .QN(buffer[0]) );
  DFFSX1 out_sel_reg ( .D(n5156), .CK(clk), .SN(rst_n), .QN(out_sel) );
  DFFSX1 U1_pipe0_reg_4_ ( .D(n5155), .CK(clk), .SN(rst_n), .QN(U1_pipe0[4])
         );
  DFFSX1 U1_pipe1_reg_23_ ( .D(n5154), .CK(clk), .SN(rst_n), .QN(U1_pipe1[23])
         );
  DFFSX1 U1_pipe1_reg_22_ ( .D(n5153), .CK(clk), .SN(rst_n), .QN(U1_pipe1[22])
         );
  DFFSX1 U1_pipe1_reg_21_ ( .D(n5152), .CK(clk), .SN(rst_n), .QN(U1_pipe1[21])
         );
  DFFSX1 U1_pipe1_reg_20_ ( .D(n5151), .CK(clk), .SN(rst_n), .QN(U1_pipe1[20])
         );
  DFFSX1 U1_pipe1_reg_19_ ( .D(n5150), .CK(clk), .SN(rst_n), .QN(U1_pipe1[19])
         );
  DFFSX1 U1_pipe1_reg_18_ ( .D(n5149), .CK(clk), .SN(rst_n), .QN(U1_pipe1[18])
         );
  DFFSX1 U1_pipe1_reg_17_ ( .D(n5148), .CK(clk), .SN(rst_n), .QN(U1_pipe1[17])
         );
  DFFSX1 U1_pipe1_reg_16_ ( .D(n5147), .CK(clk), .SN(rst_n), .QN(U1_pipe1[16])
         );
  DFFSX1 U1_pipe1_reg_15_ ( .D(n5146), .CK(clk), .SN(rst_n), .QN(U1_pipe1[15])
         );
  DFFSX1 U1_pipe1_reg_14_ ( .D(n5145), .CK(clk), .SN(rst_n), .QN(U1_pipe1[14])
         );
  DFFSX1 U1_pipe1_reg_13_ ( .D(n5144), .CK(clk), .SN(rst_n), .QN(U1_pipe1[13])
         );
  DFFSX1 U1_pipe1_reg_12_ ( .D(n5143), .CK(clk), .SN(rst_n), .QN(U1_pipe1[12])
         );
  DFFSX1 U1_pipe1_reg_11_ ( .D(n5142), .CK(clk), .SN(rst_n), .QN(U1_pipe1[11])
         );
  DFFSX1 U1_pipe1_reg_10_ ( .D(n5141), .CK(clk), .SN(rst_n), .QN(U1_pipe1[10])
         );
  DFFSX1 U1_pipe1_reg_9_ ( .D(n5140), .CK(clk), .SN(rst_n), .QN(U1_pipe1[9])
         );
  DFFSX1 U1_pipe1_reg_8_ ( .D(n5139), .CK(clk), .SN(rst_n), .QN(U1_pipe1[8])
         );
  DFFSX1 U1_pipe1_reg_7_ ( .D(n5138), .CK(clk), .SN(rst_n), .QN(U1_pipe1[7])
         );
  DFFSX1 U1_pipe1_reg_6_ ( .D(n5137), .CK(clk), .SN(rst_n), .QN(U1_pipe1[6])
         );
  DFFSX1 U1_pipe1_reg_5_ ( .D(n5136), .CK(clk), .SN(rst_n), .QN(U1_pipe1[5])
         );
  DFFSX1 U1_pipe1_reg_4_ ( .D(n5135), .CK(clk), .SN(rst_n), .QN(U1_pipe1[4])
         );
  DFFSX1 U1_pipe1_reg_3_ ( .D(n5134), .CK(clk), .SN(rst_n), .QN(U1_pipe1[3])
         );
  DFFSX1 U1_pipe1_reg_2_ ( .D(n5133), .CK(clk), .SN(rst_n), .QN(U1_pipe1[2])
         );
  DFFSX1 U1_pipe1_reg_1_ ( .D(n5132), .CK(clk), .SN(rst_n), .QN(U1_pipe1[1])
         );
  DFFSX1 U1_pipe1_reg_0_ ( .D(n5131), .CK(clk), .SN(rst_n), .QN(U1_pipe1[0])
         );
  DFFSX1 U1_pipe0_reg_24_ ( .D(n5127), .CK(clk), .SN(rst_n), .QN(U1_pipe0[24])
         );
  DFFSX1 U1_pipe0_reg_23_ ( .D(n5126), .CK(clk), .SN(rst_n), .QN(U1_pipe0[23])
         );
  DFFSX1 U1_pipe0_reg_22_ ( .D(n5125), .CK(clk), .SN(rst_n), .QN(U1_pipe0[22])
         );
  DFFSX1 U1_pipe0_reg_21_ ( .D(n5124), .CK(clk), .SN(rst_n), .QN(U1_pipe0[21])
         );
  DFFSX1 U1_pipe0_reg_20_ ( .D(n5123), .CK(clk), .SN(rst_n), .QN(U1_pipe0[20])
         );
  DFFSX1 U1_pipe0_reg_19_ ( .D(n5122), .CK(clk), .SN(rst_n), .QN(U1_pipe0[19])
         );
  DFFSX1 U1_pipe0_reg_18_ ( .D(n5121), .CK(clk), .SN(rst_n), .QN(U1_pipe0[18])
         );
  DFFSX1 U1_pipe0_reg_17_ ( .D(n5120), .CK(clk), .SN(rst_n), .QN(U1_pipe0[17])
         );
  DFFSX1 U1_pipe0_reg_16_ ( .D(n5119), .CK(clk), .SN(rst_n), .QN(U1_pipe0[16])
         );
  DFFSX1 U1_pipe0_reg_15_ ( .D(n5118), .CK(clk), .SN(rst_n), .QN(U1_pipe0[15])
         );
  DFFSX1 U1_pipe0_reg_14_ ( .D(n5117), .CK(clk), .SN(rst_n), .QN(U1_pipe0[14])
         );
  DFFSX1 U1_pipe0_reg_13_ ( .D(n5116), .CK(clk), .SN(rst_n), .QN(U1_pipe0[13])
         );
  DFFSX1 U1_pipe0_reg_12_ ( .D(n5115), .CK(clk), .SN(rst_n), .QN(U1_pipe0[12])
         );
  DFFSX1 U1_pipe0_reg_11_ ( .D(n5114), .CK(clk), .SN(rst_n), .QN(U1_pipe0[11])
         );
  DFFSX1 U1_pipe0_reg_10_ ( .D(n5113), .CK(clk), .SN(rst_n), .QN(U1_pipe0[10])
         );
  DFFSX1 U1_pipe0_reg_9_ ( .D(n5112), .CK(clk), .SN(rst_n), .QN(U1_pipe0[9])
         );
  DFFSX1 U1_pipe0_reg_8_ ( .D(n5111), .CK(clk), .SN(rst_n), .QN(U1_pipe0[8])
         );
  DFFSX1 U1_pipe0_reg_7_ ( .D(n5110), .CK(clk), .SN(rst_n), .QN(U1_pipe0[7])
         );
  DFFSX1 U1_pipe0_reg_6_ ( .D(n5109), .CK(clk), .SN(rst_n), .QN(U1_pipe0[6])
         );
  DFFSX1 U1_pipe0_reg_5_ ( .D(n5108), .CK(clk), .SN(rst_n), .QN(U1_pipe0[5])
         );
  DFFSX1 U1_pipe0_reg_3_ ( .D(n5107), .CK(clk), .SN(rst_n), .QN(U1_pipe0[3])
         );
  DFFSX1 U1_pipe5_reg_10_ ( .D(n5106), .CK(clk), .SN(rst_n), .QN(U1_pipe5[10])
         );
  DFFSX1 U1_pipe5_reg_9_ ( .D(n5105), .CK(clk), .SN(rst_n), .QN(U1_pipe5[9])
         );
  DFFSX1 U1_pipe5_reg_8_ ( .D(n5104), .CK(clk), .SN(rst_n), .QN(U1_pipe5[8])
         );
  DFFSX1 U1_pipe5_reg_7_ ( .D(n5103), .CK(clk), .SN(rst_n), .QN(U1_pipe5[7])
         );
  DFFSX1 U1_pipe5_reg_6_ ( .D(n5102), .CK(clk), .SN(rst_n), .QN(U1_pipe5[6])
         );
  DFFSX1 U1_pipe5_reg_5_ ( .D(n5101), .CK(clk), .SN(rst_n), .QN(U1_pipe5[5])
         );
  DFFSX1 U1_pipe5_reg_4_ ( .D(n5100), .CK(clk), .SN(rst_n), .QN(U1_pipe5[4])
         );
  DFFSX1 U1_pipe5_reg_3_ ( .D(n5099), .CK(clk), .SN(rst_n), .QN(U1_pipe5[3])
         );
  DFFSX1 U1_pipe5_reg_2_ ( .D(n5098), .CK(clk), .SN(rst_n), .QN(U1_pipe5[2])
         );
  DFFSX1 U1_pipe5_reg_1_ ( .D(n5097), .CK(clk), .SN(rst_n), .QN(U1_pipe5[1])
         );
  DFFSX1 U1_pipe5_reg_0_ ( .D(n5096), .CK(clk), .SN(rst_n), .QN(U1_pipe5[0])
         );
  DFFSX1 U1_pipe4_reg_25_ ( .D(n5093), .CK(clk), .SN(rst_n), .QN(U1_pipe4[25])
         );
  DFFSX1 U1_pipe4_reg_24_ ( .D(n5092), .CK(clk), .SN(rst_n), .QN(U1_pipe4[24])
         );
  DFFSX1 U1_pipe4_reg_22_ ( .D(n5090), .CK(clk), .SN(rst_n), .QN(U1_pipe4[22])
         );
  DFFSX1 U1_pipe4_reg_21_ ( .D(n5089), .CK(clk), .SN(rst_n), .QN(U1_pipe4[21])
         );
  DFFSX1 U1_pipe4_reg_20_ ( .D(n5088), .CK(clk), .SN(rst_n), .QN(U1_pipe4[20])
         );
  DFFSX1 U1_pipe4_reg_19_ ( .D(n5087), .CK(clk), .SN(rst_n), .QN(U1_pipe4[19])
         );
  DFFSX1 U1_pipe4_reg_18_ ( .D(n5086), .CK(clk), .SN(rst_n), .QN(U1_pipe4[18])
         );
  DFFSX1 U1_pipe4_reg_17_ ( .D(n5085), .CK(clk), .SN(rst_n), .QN(U1_pipe4[17])
         );
  DFFSX1 U1_pipe4_reg_16_ ( .D(n5084), .CK(clk), .SN(rst_n), .QN(U1_pipe4[16])
         );
  DFFSX1 U1_pipe4_reg_15_ ( .D(n5083), .CK(clk), .SN(rst_n), .QN(U1_pipe4[15])
         );
  DFFSX1 U1_pipe4_reg_14_ ( .D(n5082), .CK(clk), .SN(rst_n), .QN(U1_pipe4[14])
         );
  DFFSX1 U1_pipe4_reg_13_ ( .D(n5081), .CK(clk), .SN(rst_n), .QN(U1_pipe4[13])
         );
  DFFSX1 U1_pipe4_reg_12_ ( .D(n5080), .CK(clk), .SN(rst_n), .QN(U1_pipe4[12])
         );
  DFFSX1 U1_pipe4_reg_11_ ( .D(n5079), .CK(clk), .SN(rst_n), .QN(U1_pipe4[11])
         );
  DFFSX1 U1_pipe4_reg_10_ ( .D(n5078), .CK(clk), .SN(rst_n), .QN(U1_pipe4[10])
         );
  DFFSX1 U1_pipe4_reg_9_ ( .D(n5077), .CK(clk), .SN(rst_n), .QN(U1_pipe4[9])
         );
  DFFSX1 U1_pipe4_reg_8_ ( .D(n5076), .CK(clk), .SN(rst_n), .QN(U1_pipe4[8])
         );
  DFFSX1 U1_pipe4_reg_7_ ( .D(n5075), .CK(clk), .SN(rst_n), .QN(U1_pipe4[7])
         );
  DFFSX1 U1_pipe4_reg_6_ ( .D(n5074), .CK(clk), .SN(rst_n), .QN(U1_pipe4[6])
         );
  DFFSX1 U1_pipe4_reg_5_ ( .D(n5073), .CK(clk), .SN(rst_n), .QN(U1_pipe4[5])
         );
  DFFSX1 U1_pipe4_reg_4_ ( .D(n5072), .CK(clk), .SN(rst_n), .QN(U1_pipe4[4])
         );
  DFFSX1 U1_pipe4_reg_3_ ( .D(n5071), .CK(clk), .SN(rst_n), .QN(U1_pipe4[3])
         );
  DFFSX1 U1_pipe4_reg_2_ ( .D(n5070), .CK(clk), .SN(rst_n), .QN(U1_pipe4[2])
         );
  DFFSX1 U1_pipe4_reg_1_ ( .D(n5069), .CK(clk), .SN(rst_n), .Q(n28893), .QN(
        U1_pipe4[1]) );
  DFFSX1 U1_pipe4_reg_0_ ( .D(n5068), .CK(clk), .SN(rst_n), .QN(U1_pipe4[0])
         );
  DFFSX1 U1_pipe3_reg_27_ ( .D(n5067), .CK(clk), .SN(rst_n), .QN(U1_pipe3[27])
         );
  DFFSX1 U1_pipe3_reg_25_ ( .D(n5065), .CK(clk), .SN(rst_n), .Q(n28943), .QN(
        U1_pipe3[25]) );
  DFFSX1 U1_pipe3_reg_21_ ( .D(n5061), .CK(clk), .SN(rst_n), .Q(n28840), .QN(
        U1_pipe3[21]) );
  DFFSX1 U1_pipe3_reg_15_ ( .D(n5055), .CK(clk), .SN(rst_n), .Q(n28846), .QN(
        U1_pipe3[15]) );
  DFFSX1 U1_pipe3_reg_14_ ( .D(n5054), .CK(clk), .SN(rst_n), .Q(n28847), .QN(
        U1_pipe3[14]) );
  DFFSX1 U1_pipe3_reg_13_ ( .D(n5053), .CK(clk), .SN(rst_n), .Q(n28848), .QN(
        U1_pipe3[13]) );
  DFFSX1 U1_pipe3_reg_12_ ( .D(n5052), .CK(clk), .SN(rst_n), .Q(n28849), .QN(
        U1_pipe3[12]) );
  DFFSX1 U1_pipe3_reg_11_ ( .D(n5051), .CK(clk), .SN(rst_n), .Q(n28850), .QN(
        U1_pipe3[11]) );
  DFFSX1 U1_pipe3_reg_10_ ( .D(n5050), .CK(clk), .SN(rst_n), .Q(n28851), .QN(
        U1_pipe3[10]) );
  DFFSX1 U1_pipe3_reg_9_ ( .D(n5049), .CK(clk), .SN(rst_n), .Q(n28733), .QN(
        U1_pipe3[9]) );
  DFFSX1 U1_pipe3_reg_8_ ( .D(n5048), .CK(clk), .SN(rst_n), .Q(n28852), .QN(
        U1_pipe3[8]) );
  DFFSX1 U1_pipe3_reg_7_ ( .D(n5047), .CK(clk), .SN(rst_n), .Q(n28853), .QN(
        U1_pipe3[7]) );
  DFFSX1 U1_pipe3_reg_6_ ( .D(n5046), .CK(clk), .SN(rst_n), .Q(n28734), .QN(
        U1_pipe3[6]) );
  DFFSX1 U1_pipe3_reg_5_ ( .D(n5045), .CK(clk), .SN(rst_n), .Q(n28854), .QN(
        U1_pipe3[5]) );
  DFFSX1 U1_pipe3_reg_4_ ( .D(n5044), .CK(clk), .SN(rst_n), .Q(n28855), .QN(
        U1_pipe3[4]) );
  DFFSX1 U1_pipe3_reg_3_ ( .D(n5043), .CK(clk), .SN(rst_n), .Q(n28735), .QN(
        U1_pipe3[3]) );
  DFFSX1 U1_pipe3_reg_2_ ( .D(n5042), .CK(clk), .SN(rst_n), .Q(n28736), .QN(
        U1_pipe3[2]) );
  DFFSX1 U1_pipe3_reg_1_ ( .D(n5041), .CK(clk), .SN(rst_n), .Q(n28901), .QN(
        U1_pipe3[1]) );
  DFFSX1 U1_pipe3_reg_0_ ( .D(n5040), .CK(clk), .SN(rst_n), .Q(n28909), .QN(
        U1_pipe3[0]) );
  DFFSX1 U1_pipe2_reg_21_ ( .D(n5033), .CK(clk), .SN(rst_n), .QN(U1_pipe2[21])
         );
  DFFSX1 U1_pipe2_reg_20_ ( .D(n5032), .CK(clk), .SN(rst_n), .QN(U1_pipe2[20])
         );
  DFFSX1 U1_pipe2_reg_19_ ( .D(n5031), .CK(clk), .SN(rst_n), .QN(U1_pipe2[19])
         );
  DFFSX1 U1_pipe2_reg_18_ ( .D(n5030), .CK(clk), .SN(rst_n), .QN(U1_pipe2[18])
         );
  DFFSX1 U1_pipe2_reg_17_ ( .D(n5029), .CK(clk), .SN(rst_n), .QN(U1_pipe2[17])
         );
  DFFSX1 U1_pipe2_reg_16_ ( .D(n5028), .CK(clk), .SN(rst_n), .QN(U1_pipe2[16])
         );
  DFFSX1 U1_pipe2_reg_15_ ( .D(n5027), .CK(clk), .SN(rst_n), .QN(U1_pipe2[15])
         );
  DFFSX1 U1_pipe2_reg_14_ ( .D(n5026), .CK(clk), .SN(rst_n), .QN(U1_pipe2[14])
         );
  DFFSX1 U1_pipe2_reg_13_ ( .D(n5025), .CK(clk), .SN(rst_n), .QN(U1_pipe2[13])
         );
  DFFSX1 U1_pipe2_reg_12_ ( .D(n5024), .CK(clk), .SN(rst_n), .QN(U1_pipe2[12])
         );
  DFFSX1 U1_pipe2_reg_11_ ( .D(n5023), .CK(clk), .SN(rst_n), .QN(U1_pipe2[11])
         );
  DFFSX1 U1_pipe2_reg_10_ ( .D(n5022), .CK(clk), .SN(rst_n), .QN(U1_pipe2[10])
         );
  DFFSX1 U1_pipe2_reg_9_ ( .D(n5021), .CK(clk), .SN(rst_n), .QN(U1_pipe2[9])
         );
  DFFSX1 U1_pipe2_reg_8_ ( .D(n5020), .CK(clk), .SN(rst_n), .QN(U1_pipe2[8])
         );
  DFFSX1 U1_pipe2_reg_7_ ( .D(n5019), .CK(clk), .SN(rst_n), .QN(U1_pipe2[7])
         );
  DFFSX1 U1_pipe2_reg_6_ ( .D(n5018), .CK(clk), .SN(rst_n), .QN(U1_pipe2[6])
         );
  DFFSX1 U1_pipe2_reg_5_ ( .D(n5017), .CK(clk), .SN(rst_n), .QN(U1_pipe2[5])
         );
  DFFSX1 U1_pipe2_reg_4_ ( .D(n5016), .CK(clk), .SN(rst_n), .QN(U1_pipe2[4])
         );
  DFFSX1 U1_pipe2_reg_3_ ( .D(n5015), .CK(clk), .SN(rst_n), .QN(U1_pipe2[3])
         );
  DFFSX1 U1_pipe2_reg_2_ ( .D(n5014), .CK(clk), .SN(rst_n), .QN(U1_pipe2[2])
         );
  DFFSX1 U1_pipe2_reg_1_ ( .D(n5013), .CK(clk), .SN(rst_n), .QN(U1_pipe2[1])
         );
  DFFSX1 U1_pipe2_reg_0_ ( .D(n5012), .CK(clk), .SN(rst_n), .QN(U1_pipe2[0])
         );
  DFFSX1 U1_pipe1_reg_26_ ( .D(n5010), .CK(clk), .SN(rst_n), .QN(U1_pipe1[26])
         );
  DFFSX1 U1_pipe1_reg_25_ ( .D(n5009), .CK(clk), .SN(rst_n), .QN(U1_pipe1[25])
         );
  DFFSX1 U1_pipe1_reg_24_ ( .D(n5008), .CK(clk), .SN(rst_n), .QN(U1_pipe1[24])
         );
  DFFSX1 U1_pipe0_reg_2_ ( .D(n5007), .CK(clk), .SN(rst_n), .QN(U1_pipe0[2])
         );
  DFFSX1 U1_pipe8_reg_25_ ( .D(n5006), .CK(clk), .SN(rst_n), .QN(U1_pipe8[25])
         );
  DFFSX1 U1_pipe8_reg_24_ ( .D(n5005), .CK(clk), .SN(rst_n), .QN(U1_pipe8[24])
         );
  DFFSX1 U1_pipe8_reg_23_ ( .D(n5004), .CK(clk), .SN(rst_n), .QN(U1_pipe8[23])
         );
  DFFSX1 U1_pipe8_reg_22_ ( .D(n5003), .CK(clk), .SN(rst_n), .QN(U1_pipe8[22])
         );
  DFFSX1 U1_pipe8_reg_21_ ( .D(n5002), .CK(clk), .SN(rst_n), .QN(U1_pipe8[21])
         );
  DFFSX1 U1_pipe8_reg_20_ ( .D(n5001), .CK(clk), .SN(rst_n), .QN(U1_pipe8[20])
         );
  DFFSX1 U1_pipe8_reg_19_ ( .D(n5000), .CK(clk), .SN(rst_n), .QN(U1_pipe8[19])
         );
  DFFSX1 U1_pipe8_reg_18_ ( .D(n4999), .CK(clk), .SN(rst_n), .QN(U1_pipe8[18])
         );
  DFFSX1 U1_pipe8_reg_17_ ( .D(n4998), .CK(clk), .SN(rst_n), .QN(U1_pipe8[17])
         );
  DFFSX1 U1_pipe8_reg_16_ ( .D(n4997), .CK(clk), .SN(rst_n), .QN(U1_pipe8[16])
         );
  DFFSX1 U1_pipe8_reg_15_ ( .D(n4996), .CK(clk), .SN(rst_n), .QN(U1_pipe8[15])
         );
  DFFSX1 U1_pipe8_reg_14_ ( .D(n4995), .CK(clk), .SN(rst_n), .QN(U1_pipe8[14])
         );
  DFFSX1 U1_pipe8_reg_13_ ( .D(n4994), .CK(clk), .SN(rst_n), .QN(U1_pipe8[13])
         );
  DFFSX1 U1_pipe8_reg_12_ ( .D(n4993), .CK(clk), .SN(rst_n), .QN(U1_pipe8[12])
         );
  DFFSX1 U1_pipe8_reg_11_ ( .D(n4992), .CK(clk), .SN(rst_n), .QN(U1_pipe8[11])
         );
  DFFSX1 U1_pipe8_reg_10_ ( .D(n4991), .CK(clk), .SN(rst_n), .QN(U1_pipe8[10])
         );
  DFFSX1 U1_pipe8_reg_9_ ( .D(n4990), .CK(clk), .SN(rst_n), .QN(U1_pipe8[9])
         );
  DFFSX1 U1_pipe8_reg_8_ ( .D(n4989), .CK(clk), .SN(rst_n), .QN(U1_pipe8[8])
         );
  DFFSX1 U1_pipe8_reg_7_ ( .D(n4988), .CK(clk), .SN(rst_n), .QN(U1_pipe8[7])
         );
  DFFSX1 U1_pipe8_reg_6_ ( .D(n4987), .CK(clk), .SN(rst_n), .QN(U1_pipe8[6])
         );
  DFFSX1 U1_pipe8_reg_5_ ( .D(n4986), .CK(clk), .SN(rst_n), .QN(U1_pipe8[5])
         );
  DFFSX1 U1_pipe8_reg_4_ ( .D(n4985), .CK(clk), .SN(rst_n), .QN(U1_pipe8[4])
         );
  DFFSX1 U1_pipe8_reg_3_ ( .D(n4984), .CK(clk), .SN(rst_n), .QN(U1_pipe8[3])
         );
  DFFSX1 U1_pipe8_reg_2_ ( .D(n4983), .CK(clk), .SN(rst_n), .QN(U1_pipe8[2])
         );
  DFFSX1 U1_pipe8_reg_1_ ( .D(n4982), .CK(clk), .SN(rst_n), .QN(U1_pipe8[1])
         );
  DFFSX1 U1_pipe8_reg_0_ ( .D(n4981), .CK(clk), .SN(rst_n), .QN(U1_pipe8[0])
         );
  DFFSX1 U1_pipe7_reg_26_ ( .D(n4979), .CK(clk), .SN(rst_n), .QN(U1_pipe7[26])
         );
  DFFSX1 U1_pipe7_reg_25_ ( .D(n4978), .CK(clk), .SN(rst_n), .QN(U1_pipe7[25])
         );
  DFFSX1 U1_pipe7_reg_24_ ( .D(n4977), .CK(clk), .SN(rst_n), .QN(U1_pipe7[24])
         );
  DFFSX1 U1_pipe7_reg_23_ ( .D(n4976), .CK(clk), .SN(rst_n), .QN(U1_pipe7[23])
         );
  DFFSX1 U1_pipe7_reg_22_ ( .D(n4975), .CK(clk), .SN(rst_n), .QN(U1_pipe7[22])
         );
  DFFSX1 U1_pipe7_reg_21_ ( .D(n4974), .CK(clk), .SN(rst_n), .QN(U1_pipe7[21])
         );
  DFFSX1 U1_pipe7_reg_20_ ( .D(n4973), .CK(clk), .SN(rst_n), .QN(U1_pipe7[20])
         );
  DFFSX1 U1_pipe7_reg_19_ ( .D(n4972), .CK(clk), .SN(rst_n), .QN(U1_pipe7[19])
         );
  DFFSX1 U1_pipe7_reg_18_ ( .D(n4971), .CK(clk), .SN(rst_n), .QN(U1_pipe7[18])
         );
  DFFSX1 U1_pipe7_reg_17_ ( .D(n4970), .CK(clk), .SN(rst_n), .QN(U1_pipe7[17])
         );
  DFFSX1 U1_pipe7_reg_16_ ( .D(n4969), .CK(clk), .SN(rst_n), .QN(U1_pipe7[16])
         );
  DFFSX1 U1_pipe7_reg_15_ ( .D(n4968), .CK(clk), .SN(rst_n), .QN(U1_pipe7[15])
         );
  DFFSX1 U1_pipe7_reg_14_ ( .D(n4967), .CK(clk), .SN(rst_n), .QN(U1_pipe7[14])
         );
  DFFSX1 U1_pipe7_reg_13_ ( .D(n4966), .CK(clk), .SN(rst_n), .QN(U1_pipe7[13])
         );
  DFFSX1 U1_pipe7_reg_12_ ( .D(n4965), .CK(clk), .SN(rst_n), .QN(U1_pipe7[12])
         );
  DFFSX1 U1_pipe7_reg_11_ ( .D(n4964), .CK(clk), .SN(rst_n), .QN(U1_pipe7[11])
         );
  DFFSX1 U1_pipe7_reg_10_ ( .D(n4963), .CK(clk), .SN(rst_n), .QN(U1_pipe7[10])
         );
  DFFSX1 U1_pipe7_reg_9_ ( .D(n4962), .CK(clk), .SN(rst_n), .QN(U1_pipe7[9])
         );
  DFFSX1 U1_pipe7_reg_8_ ( .D(n4961), .CK(clk), .SN(rst_n), .QN(U1_pipe7[8])
         );
  DFFSX1 U1_pipe7_reg_7_ ( .D(n4960), .CK(clk), .SN(rst_n), .QN(U1_pipe7[7])
         );
  DFFSX1 U1_pipe7_reg_6_ ( .D(n4959), .CK(clk), .SN(rst_n), .QN(U1_pipe7[6])
         );
  DFFSX1 U1_pipe7_reg_5_ ( .D(n4958), .CK(clk), .SN(rst_n), .QN(U1_pipe7[5])
         );
  DFFSX1 U1_pipe7_reg_4_ ( .D(n4957), .CK(clk), .SN(rst_n), .QN(U1_pipe7[4])
         );
  DFFSX1 U1_pipe7_reg_3_ ( .D(n4956), .CK(clk), .SN(rst_n), .QN(U1_pipe7[3])
         );
  DFFSX1 U1_pipe7_reg_2_ ( .D(n4955), .CK(clk), .SN(rst_n), .QN(U1_pipe7[2])
         );
  DFFSX1 U1_pipe7_reg_1_ ( .D(n4954), .CK(clk), .SN(rst_n), .QN(U1_pipe7[1])
         );
  DFFSX1 U1_pipe7_reg_0_ ( .D(n4953), .CK(clk), .SN(rst_n), .QN(U1_pipe7[0])
         );
  DFFSX1 U1_pipe6_reg_26_ ( .D(n4951), .CK(clk), .SN(rst_n), .QN(U1_pipe6[26])
         );
  DFFSX1 U1_pipe6_reg_25_ ( .D(n4950), .CK(clk), .SN(rst_n), .QN(U1_pipe6[25])
         );
  DFFSX1 U1_pipe6_reg_24_ ( .D(n4949), .CK(clk), .SN(rst_n), .QN(U1_pipe6[24])
         );
  DFFSX1 U1_pipe6_reg_23_ ( .D(n4948), .CK(clk), .SN(rst_n), .QN(U1_pipe6[23])
         );
  DFFSX1 U1_pipe6_reg_21_ ( .D(n4946), .CK(clk), .SN(rst_n), .QN(U1_pipe6[21])
         );
  DFFSX1 U1_pipe6_reg_20_ ( .D(n4945), .CK(clk), .SN(rst_n), .QN(U1_pipe6[20])
         );
  DFFSX1 U1_pipe6_reg_19_ ( .D(n4944), .CK(clk), .SN(rst_n), .QN(U1_pipe6[19])
         );
  DFFSX1 U1_pipe6_reg_18_ ( .D(n4943), .CK(clk), .SN(rst_n), .QN(U1_pipe6[18])
         );
  DFFSX1 U1_pipe6_reg_17_ ( .D(n4942), .CK(clk), .SN(rst_n), .QN(U1_pipe6[17])
         );
  DFFSX1 U1_pipe6_reg_16_ ( .D(n4941), .CK(clk), .SN(rst_n), .QN(U1_pipe6[16])
         );
  DFFSX1 U1_pipe6_reg_15_ ( .D(n4940), .CK(clk), .SN(rst_n), .QN(U1_pipe6[15])
         );
  DFFSX1 U1_pipe6_reg_14_ ( .D(n4939), .CK(clk), .SN(rst_n), .QN(U1_pipe6[14])
         );
  DFFSX1 U1_pipe6_reg_13_ ( .D(n4938), .CK(clk), .SN(rst_n), .QN(U1_pipe6[13])
         );
  DFFSX1 U1_pipe6_reg_12_ ( .D(n4937), .CK(clk), .SN(rst_n), .QN(U1_pipe6[12])
         );
  DFFSX1 U1_pipe6_reg_11_ ( .D(n4936), .CK(clk), .SN(rst_n), .QN(U1_pipe6[11])
         );
  DFFSX1 U1_pipe6_reg_10_ ( .D(n4935), .CK(clk), .SN(rst_n), .QN(U1_pipe6[10])
         );
  DFFSX1 U1_pipe6_reg_9_ ( .D(n4934), .CK(clk), .SN(rst_n), .QN(U1_pipe6[9])
         );
  DFFSX1 U1_pipe6_reg_8_ ( .D(n4933), .CK(clk), .SN(rst_n), .QN(U1_pipe6[8])
         );
  DFFSX1 U1_pipe6_reg_7_ ( .D(n4932), .CK(clk), .SN(rst_n), .QN(U1_pipe6[7])
         );
  DFFSX1 U1_pipe6_reg_6_ ( .D(n4931), .CK(clk), .SN(rst_n), .QN(U1_pipe6[6])
         );
  DFFSX1 U1_pipe6_reg_5_ ( .D(n4930), .CK(clk), .SN(rst_n), .QN(U1_pipe6[5])
         );
  DFFSX1 U1_pipe6_reg_4_ ( .D(n4929), .CK(clk), .SN(rst_n), .QN(U1_pipe6[4])
         );
  DFFSX1 U1_pipe6_reg_3_ ( .D(n4928), .CK(clk), .SN(rst_n), .QN(U1_pipe6[3])
         );
  DFFSX1 U1_pipe6_reg_2_ ( .D(n4927), .CK(clk), .SN(rst_n), .QN(U1_pipe6[2])
         );
  DFFSX1 U1_pipe6_reg_1_ ( .D(n4926), .CK(clk), .SN(rst_n), .Q(n28895), .QN(
        U1_pipe6[1]) );
  DFFSX1 U1_pipe6_reg_0_ ( .D(n4925), .CK(clk), .SN(rst_n), .QN(U1_pipe6[0])
         );
  DFFSX1 U1_pipe5_reg_27_ ( .D(n4924), .CK(clk), .SN(rst_n), .Q(n28694), .QN(
        U1_pipe5[27]) );
  DFFSX1 U1_pipe5_reg_26_ ( .D(n4923), .CK(clk), .SN(rst_n), .QN(U1_pipe5[26])
         );
  DFFSX1 U1_pipe5_reg_25_ ( .D(n4922), .CK(clk), .SN(rst_n), .QN(U1_pipe5[25])
         );
  DFFSX1 U1_pipe5_reg_24_ ( .D(n4921), .CK(clk), .SN(rst_n), .QN(U1_pipe5[24])
         );
  DFFSX1 U1_pipe5_reg_23_ ( .D(n4920), .CK(clk), .SN(rst_n), .QN(U1_pipe5[23])
         );
  DFFSX1 U1_pipe5_reg_22_ ( .D(n4919), .CK(clk), .SN(rst_n), .QN(U1_pipe5[22])
         );
  DFFSX1 U1_pipe5_reg_21_ ( .D(n4918), .CK(clk), .SN(rst_n), .QN(U1_pipe5[21])
         );
  DFFSX1 U1_pipe5_reg_20_ ( .D(n4917), .CK(clk), .SN(rst_n), .QN(U1_pipe5[20])
         );
  DFFSX1 U1_pipe5_reg_19_ ( .D(n4916), .CK(clk), .SN(rst_n), .QN(U1_pipe5[19])
         );
  DFFSX1 U1_pipe5_reg_18_ ( .D(n4915), .CK(clk), .SN(rst_n), .QN(U1_pipe5[18])
         );
  DFFSX1 U1_pipe5_reg_17_ ( .D(n4914), .CK(clk), .SN(rst_n), .QN(U1_pipe5[17])
         );
  DFFSX1 U1_pipe5_reg_16_ ( .D(n4913), .CK(clk), .SN(rst_n), .QN(U1_pipe5[16])
         );
  DFFSX1 U1_pipe5_reg_15_ ( .D(n4912), .CK(clk), .SN(rst_n), .QN(U1_pipe5[15])
         );
  DFFSX1 U1_pipe5_reg_14_ ( .D(n4911), .CK(clk), .SN(rst_n), .QN(U1_pipe5[14])
         );
  DFFSX1 U1_pipe5_reg_13_ ( .D(n4910), .CK(clk), .SN(rst_n), .QN(U1_pipe5[13])
         );
  DFFSX1 U1_pipe5_reg_12_ ( .D(n4909), .CK(clk), .SN(rst_n), .QN(U1_pipe5[12])
         );
  DFFSX1 U1_pipe5_reg_11_ ( .D(n4908), .CK(clk), .SN(rst_n), .QN(U1_pipe5[11])
         );
  DFFSX1 U1_pipe0_reg_1_ ( .D(n4907), .CK(clk), .SN(rst_n), .Q(n28892), .QN(
        U1_pipe0[1]) );
  DFFSX1 U1_pipe12_reg_12_ ( .D(n4906), .CK(clk), .SN(rst_n), .QN(
        U1_pipe12[12]) );
  DFFSX1 U1_pipe12_reg_11_ ( .D(n4905), .CK(clk), .SN(rst_n), .QN(
        U1_pipe12[11]) );
  DFFSX1 U1_pipe12_reg_10_ ( .D(n4904), .CK(clk), .SN(rst_n), .QN(
        U1_pipe12[10]) );
  DFFSX1 U1_pipe12_reg_9_ ( .D(n4903), .CK(clk), .SN(rst_n), .QN(U1_pipe12[9])
         );
  DFFSX1 U1_pipe12_reg_8_ ( .D(n4902), .CK(clk), .SN(rst_n), .QN(U1_pipe12[8])
         );
  DFFSX1 U1_pipe12_reg_7_ ( .D(n4901), .CK(clk), .SN(rst_n), .QN(U1_pipe12[7])
         );
  DFFSX1 U1_pipe12_reg_6_ ( .D(n4900), .CK(clk), .SN(rst_n), .QN(U1_pipe12[6])
         );
  DFFSX1 U1_pipe12_reg_5_ ( .D(n4899), .CK(clk), .SN(rst_n), .QN(U1_pipe12[5])
         );
  DFFSX1 U1_pipe12_reg_4_ ( .D(n4898), .CK(clk), .SN(rst_n), .QN(U1_pipe12[4])
         );
  DFFSX1 U1_pipe12_reg_3_ ( .D(n4897), .CK(clk), .SN(rst_n), .QN(U1_pipe12[3])
         );
  DFFSX1 U1_pipe12_reg_2_ ( .D(n4896), .CK(clk), .SN(rst_n), .QN(U1_pipe12[2])
         );
  DFFSX1 U1_pipe12_reg_1_ ( .D(n4895), .CK(clk), .SN(rst_n), .QN(U1_pipe12[1])
         );
  DFFSX1 U1_pipe12_reg_0_ ( .D(n4894), .CK(clk), .SN(rst_n), .QN(U1_pipe12[0])
         );
  DFFSX1 U1_pipe11_reg_27_ ( .D(n4893), .CK(clk), .SN(rst_n), .Q(n28695), .QN(
        U1_pipe11[27]) );
  DFFSX1 U1_pipe11_reg_26_ ( .D(n4892), .CK(clk), .SN(rst_n), .QN(
        U1_pipe11[26]) );
  DFFSX1 U1_pipe11_reg_25_ ( .D(n4891), .CK(clk), .SN(rst_n), .QN(
        U1_pipe11[25]) );
  DFFSX1 U1_pipe11_reg_24_ ( .D(n4890), .CK(clk), .SN(rst_n), .QN(
        U1_pipe11[24]) );
  DFFSX1 U1_pipe11_reg_23_ ( .D(n4889), .CK(clk), .SN(rst_n), .QN(
        U1_pipe11[23]) );
  DFFSX1 U1_pipe11_reg_22_ ( .D(n4888), .CK(clk), .SN(rst_n), .QN(
        U1_pipe11[22]) );
  DFFSX1 U1_pipe11_reg_21_ ( .D(n4887), .CK(clk), .SN(rst_n), .QN(
        U1_pipe11[21]) );
  DFFSX1 U1_pipe11_reg_20_ ( .D(n4886), .CK(clk), .SN(rst_n), .QN(
        U1_pipe11[20]) );
  DFFSX1 U1_pipe11_reg_19_ ( .D(n4885), .CK(clk), .SN(rst_n), .QN(
        U1_pipe11[19]) );
  DFFSX1 U1_pipe11_reg_18_ ( .D(n4884), .CK(clk), .SN(rst_n), .QN(
        U1_pipe11[18]) );
  DFFSX1 U1_pipe11_reg_17_ ( .D(n4883), .CK(clk), .SN(rst_n), .QN(
        U1_pipe11[17]) );
  DFFSX1 U1_pipe11_reg_16_ ( .D(n4882), .CK(clk), .SN(rst_n), .QN(
        U1_pipe11[16]) );
  DFFSX1 U1_pipe11_reg_15_ ( .D(n4881), .CK(clk), .SN(rst_n), .QN(
        U1_pipe11[15]) );
  DFFSX1 U1_pipe11_reg_14_ ( .D(n4880), .CK(clk), .SN(rst_n), .QN(
        U1_pipe11[14]) );
  DFFSX1 U1_pipe11_reg_13_ ( .D(n4879), .CK(clk), .SN(rst_n), .QN(
        U1_pipe11[13]) );
  DFFSX1 U1_pipe11_reg_12_ ( .D(n4878), .CK(clk), .SN(rst_n), .QN(
        U1_pipe11[12]) );
  DFFSX1 U1_pipe11_reg_11_ ( .D(n4877), .CK(clk), .SN(rst_n), .QN(
        U1_pipe11[11]) );
  DFFSX1 U1_pipe11_reg_10_ ( .D(n4876), .CK(clk), .SN(rst_n), .QN(
        U1_pipe11[10]) );
  DFFSX1 U1_pipe11_reg_9_ ( .D(n4875), .CK(clk), .SN(rst_n), .QN(U1_pipe11[9])
         );
  DFFSX1 U1_pipe11_reg_8_ ( .D(n4874), .CK(clk), .SN(rst_n), .QN(U1_pipe11[8])
         );
  DFFSX1 U1_pipe11_reg_7_ ( .D(n4873), .CK(clk), .SN(rst_n), .QN(U1_pipe11[7])
         );
  DFFSX1 U1_pipe11_reg_6_ ( .D(n4872), .CK(clk), .SN(rst_n), .QN(U1_pipe11[6])
         );
  DFFSX1 U1_pipe11_reg_5_ ( .D(n4871), .CK(clk), .SN(rst_n), .QN(U1_pipe11[5])
         );
  DFFSX1 U1_pipe11_reg_4_ ( .D(n4870), .CK(clk), .SN(rst_n), .QN(U1_pipe11[4])
         );
  DFFSX1 U1_pipe11_reg_3_ ( .D(n4869), .CK(clk), .SN(rst_n), .QN(U1_pipe11[3])
         );
  DFFSX1 U1_pipe11_reg_2_ ( .D(n4868), .CK(clk), .SN(rst_n), .QN(U1_pipe11[2])
         );
  DFFSX1 U1_pipe11_reg_1_ ( .D(n4867), .CK(clk), .SN(rst_n), .QN(U1_pipe11[1])
         );
  DFFSX1 U1_pipe11_reg_0_ ( .D(n4866), .CK(clk), .SN(rst_n), .QN(U1_pipe11[0])
         );
  DFFSX1 U1_pipe10_reg_20_ ( .D(n4858), .CK(clk), .SN(rst_n), .QN(
        U1_pipe10[20]) );
  DFFSX1 U1_pipe10_reg_19_ ( .D(n4857), .CK(clk), .SN(rst_n), .QN(
        U1_pipe10[19]) );
  DFFSX1 U1_pipe10_reg_18_ ( .D(n4856), .CK(clk), .SN(rst_n), .QN(
        U1_pipe10[18]) );
  DFFSX1 U1_pipe10_reg_17_ ( .D(n4855), .CK(clk), .SN(rst_n), .QN(
        U1_pipe10[17]) );
  DFFSX1 U1_pipe10_reg_16_ ( .D(n4854), .CK(clk), .SN(rst_n), .QN(
        U1_pipe10[16]) );
  DFFSX1 U1_pipe10_reg_15_ ( .D(n4853), .CK(clk), .SN(rst_n), .QN(
        U1_pipe10[15]) );
  DFFSX1 U1_pipe10_reg_14_ ( .D(n4852), .CK(clk), .SN(rst_n), .QN(
        U1_pipe10[14]) );
  DFFSX1 U1_pipe10_reg_13_ ( .D(n4851), .CK(clk), .SN(rst_n), .QN(
        U1_pipe10[13]) );
  DFFSX1 U1_pipe10_reg_12_ ( .D(n4850), .CK(clk), .SN(rst_n), .QN(
        U1_pipe10[12]) );
  DFFSX1 U1_pipe10_reg_11_ ( .D(n4849), .CK(clk), .SN(rst_n), .QN(
        U1_pipe10[11]) );
  DFFSX1 U1_pipe10_reg_10_ ( .D(n4848), .CK(clk), .SN(rst_n), .QN(
        U1_pipe10[10]) );
  DFFSX1 U1_pipe10_reg_9_ ( .D(n4847), .CK(clk), .SN(rst_n), .QN(U1_pipe10[9])
         );
  DFFSX1 U1_pipe10_reg_8_ ( .D(n4846), .CK(clk), .SN(rst_n), .QN(U1_pipe10[8])
         );
  DFFSX1 U1_pipe10_reg_7_ ( .D(n4845), .CK(clk), .SN(rst_n), .QN(U1_pipe10[7])
         );
  DFFSX1 U1_pipe10_reg_6_ ( .D(n4844), .CK(clk), .SN(rst_n), .QN(U1_pipe10[6])
         );
  DFFSX1 U1_pipe10_reg_5_ ( .D(n4843), .CK(clk), .SN(rst_n), .QN(U1_pipe10[5])
         );
  DFFSX1 U1_pipe10_reg_4_ ( .D(n4842), .CK(clk), .SN(rst_n), .QN(U1_pipe10[4])
         );
  DFFSX1 U1_pipe10_reg_3_ ( .D(n4841), .CK(clk), .SN(rst_n), .QN(U1_pipe10[3])
         );
  DFFSX1 U1_pipe10_reg_2_ ( .D(n4840), .CK(clk), .SN(rst_n), .QN(U1_pipe10[2])
         );
  DFFSX1 U1_pipe10_reg_1_ ( .D(n4839), .CK(clk), .SN(rst_n), .Q(n28894), .QN(
        U1_pipe10[1]) );
  DFFSX1 U1_pipe10_reg_0_ ( .D(n4838), .CK(clk), .SN(rst_n), .QN(U1_pipe10[0])
         );
  DFFSX1 U1_pipe9_reg_27_ ( .D(n4837), .CK(clk), .SN(rst_n), .QN(U1_pipe9[27])
         );
  DFFSX1 U1_pipe9_reg_24_ ( .D(n4834), .CK(clk), .SN(rst_n), .Q(n28940), .QN(
        U1_pipe9[24]) );
  DFFSX1 U1_pipe9_reg_23_ ( .D(n4833), .CK(clk), .SN(rst_n), .Q(n28941), .QN(
        U1_pipe9[23]) );
  DFFSX1 U1_pipe9_reg_22_ ( .D(n4832), .CK(clk), .SN(rst_n), .Q(n28942), .QN(
        U1_pipe9[22]) );
  DFFSX1 U1_pipe9_reg_21_ ( .D(n4831), .CK(clk), .SN(rst_n), .Q(n28824), .QN(
        U1_pipe9[21]) );
  DFFSX1 U1_pipe9_reg_19_ ( .D(n4829), .CK(clk), .SN(rst_n), .Q(n28826), .QN(
        U1_pipe9[19]) );
  DFFSX1 U1_pipe9_reg_18_ ( .D(n4828), .CK(clk), .SN(rst_n), .Q(n28827), .QN(
        U1_pipe9[18]) );
  DFFSX1 U1_pipe9_reg_17_ ( .D(n4827), .CK(clk), .SN(rst_n), .Q(n28828), .QN(
        U1_pipe9[17]) );
  DFFSX1 U1_pipe9_reg_16_ ( .D(n4826), .CK(clk), .SN(rst_n), .Q(n28829), .QN(
        U1_pipe9[16]) );
  DFFSX1 U1_pipe9_reg_15_ ( .D(n4825), .CK(clk), .SN(rst_n), .Q(n28830), .QN(
        U1_pipe9[15]) );
  DFFSX1 U1_pipe9_reg_14_ ( .D(n4824), .CK(clk), .SN(rst_n), .Q(n28831), .QN(
        U1_pipe9[14]) );
  DFFSX1 U1_pipe9_reg_13_ ( .D(n4823), .CK(clk), .SN(rst_n), .Q(n28832), .QN(
        U1_pipe9[13]) );
  DFFSX1 U1_pipe9_reg_12_ ( .D(n4822), .CK(clk), .SN(rst_n), .Q(n28833), .QN(
        U1_pipe9[12]) );
  DFFSX1 U1_pipe9_reg_11_ ( .D(n4821), .CK(clk), .SN(rst_n), .Q(n28834), .QN(
        U1_pipe9[11]) );
  DFFSX1 U1_pipe9_reg_10_ ( .D(n4820), .CK(clk), .SN(rst_n), .Q(n28835), .QN(
        U1_pipe9[10]) );
  DFFSX1 U1_pipe9_reg_9_ ( .D(n4819), .CK(clk), .SN(rst_n), .Q(n28729), .QN(
        U1_pipe9[9]) );
  DFFSX1 U1_pipe9_reg_8_ ( .D(n4818), .CK(clk), .SN(rst_n), .Q(n28836), .QN(
        U1_pipe9[8]) );
  DFFSX1 U1_pipe9_reg_7_ ( .D(n4817), .CK(clk), .SN(rst_n), .Q(n28837), .QN(
        U1_pipe9[7]) );
  DFFSX1 U1_pipe9_reg_6_ ( .D(n4816), .CK(clk), .SN(rst_n), .Q(n28730), .QN(
        U1_pipe9[6]) );
  DFFSX1 U1_pipe9_reg_5_ ( .D(n4815), .CK(clk), .SN(rst_n), .Q(n28838), .QN(
        U1_pipe9[5]) );
  DFFSX1 U1_pipe9_reg_4_ ( .D(n4814), .CK(clk), .SN(rst_n), .Q(n28839), .QN(
        U1_pipe9[4]) );
  DFFSX1 U1_pipe9_reg_3_ ( .D(n4813), .CK(clk), .SN(rst_n), .Q(n28731), .QN(
        U1_pipe9[3]) );
  DFFSX1 U1_pipe9_reg_2_ ( .D(n4812), .CK(clk), .SN(rst_n), .Q(n28732), .QN(
        U1_pipe9[2]) );
  DFFSX1 U1_pipe9_reg_1_ ( .D(n4811), .CK(clk), .SN(rst_n), .Q(n28900), .QN(
        U1_pipe9[1]) );
  DFFSX1 U1_pipe9_reg_0_ ( .D(n4810), .CK(clk), .SN(rst_n), .Q(n28908), .QN(
        U1_pipe9[0]) );
  DFFSX1 U1_pipe8_reg_26_ ( .D(n4808), .CK(clk), .SN(rst_n), .QN(U1_pipe8[26])
         );
  DFFSX1 U1_pipe0_reg_0_ ( .D(n4807), .CK(clk), .SN(rst_n), .QN(U1_pipe0[0])
         );
  DFFSX1 U1_pipe15_reg_27_ ( .D(n4806), .CK(clk), .SN(rst_n), .QN(
        U1_pipe15[27]) );
  DFFSX1 U1_pipe15_reg_24_ ( .D(n4803), .CK(clk), .SN(rst_n), .Q(n28952), .QN(
        U1_pipe15[24]) );
  DFFSX1 U1_pipe15_reg_23_ ( .D(n4802), .CK(clk), .SN(rst_n), .Q(n28953), .QN(
        U1_pipe15[23]) );
  DFFSX1 U1_pipe15_reg_22_ ( .D(n4801), .CK(clk), .SN(rst_n), .Q(n28954), .QN(
        U1_pipe15[22]) );
  DFFSX1 U1_pipe15_reg_21_ ( .D(n4800), .CK(clk), .SN(rst_n), .Q(n28872), .QN(
        U1_pipe15[21]) );
  DFFSX1 U1_pipe15_reg_19_ ( .D(n4798), .CK(clk), .SN(rst_n), .Q(n28874), .QN(
        U1_pipe15[19]) );
  DFFSX1 U1_pipe15_reg_18_ ( .D(n4797), .CK(clk), .SN(rst_n), .Q(n28875), .QN(
        U1_pipe15[18]) );
  DFFSX1 U1_pipe15_reg_17_ ( .D(n4796), .CK(clk), .SN(rst_n), .Q(n28876), .QN(
        U1_pipe15[17]) );
  DFFSX1 U1_pipe15_reg_16_ ( .D(n4795), .CK(clk), .SN(rst_n), .Q(n28877), .QN(
        U1_pipe15[16]) );
  DFFSX1 U1_pipe15_reg_15_ ( .D(n4794), .CK(clk), .SN(rst_n), .Q(n28878), .QN(
        U1_pipe15[15]) );
  DFFSX1 U1_pipe15_reg_14_ ( .D(n4793), .CK(clk), .SN(rst_n), .Q(n28879), .QN(
        U1_pipe15[14]) );
  DFFSX1 U1_pipe15_reg_13_ ( .D(n4792), .CK(clk), .SN(rst_n), .Q(n28880), .QN(
        U1_pipe15[13]) );
  DFFSX1 U1_pipe15_reg_12_ ( .D(n4791), .CK(clk), .SN(rst_n), .Q(n28881), .QN(
        U1_pipe15[12]) );
  DFFSX1 U1_pipe15_reg_11_ ( .D(n4790), .CK(clk), .SN(rst_n), .Q(n28882), .QN(
        U1_pipe15[11]) );
  DFFSX1 U1_pipe15_reg_10_ ( .D(n4789), .CK(clk), .SN(rst_n), .Q(n28883), .QN(
        U1_pipe15[10]) );
  DFFSX1 U1_pipe15_reg_9_ ( .D(n4788), .CK(clk), .SN(rst_n), .Q(n28741), .QN(
        U1_pipe15[9]) );
  DFFSX1 U1_pipe15_reg_8_ ( .D(n4787), .CK(clk), .SN(rst_n), .Q(n28884), .QN(
        U1_pipe15[8]) );
  DFFSX1 U1_pipe15_reg_7_ ( .D(n4786), .CK(clk), .SN(rst_n), .Q(n28885), .QN(
        U1_pipe15[7]) );
  DFFSX1 U1_pipe15_reg_6_ ( .D(n4785), .CK(clk), .SN(rst_n), .Q(n28742), .QN(
        U1_pipe15[6]) );
  DFFSX1 U1_pipe15_reg_5_ ( .D(n4784), .CK(clk), .SN(rst_n), .Q(n28886), .QN(
        U1_pipe15[5]) );
  DFFSX1 U1_pipe15_reg_4_ ( .D(n4783), .CK(clk), .SN(rst_n), .Q(n28887), .QN(
        U1_pipe15[4]) );
  DFFSX1 U1_pipe15_reg_3_ ( .D(n4782), .CK(clk), .SN(rst_n), .Q(n28743), .QN(
        U1_pipe15[3]) );
  DFFSX1 U1_pipe15_reg_2_ ( .D(n4781), .CK(clk), .SN(rst_n), .Q(n28744), .QN(
        U1_pipe15[2]) );
  DFFSX1 U1_pipe15_reg_1_ ( .D(n4780), .CK(clk), .SN(rst_n), .Q(n28903), .QN(
        U1_pipe15[1]) );
  DFFSX1 U1_pipe15_reg_0_ ( .D(n4779), .CK(clk), .SN(rst_n), .Q(n28911), .QN(
        U1_pipe15[0]) );
  DFFSX1 U1_pipe14_reg_24_ ( .D(n4775), .CK(clk), .SN(rst_n), .QN(
        U1_pipe14[24]) );
  DFFSX1 U1_pipe14_reg_21_ ( .D(n4772), .CK(clk), .SN(rst_n), .QN(
        U1_pipe14[21]) );
  DFFSX1 U1_pipe14_reg_20_ ( .D(n4771), .CK(clk), .SN(rst_n), .QN(
        U1_pipe14[20]) );
  DFFSX1 U1_pipe14_reg_19_ ( .D(n4770), .CK(clk), .SN(rst_n), .QN(
        U1_pipe14[19]) );
  DFFSX1 U1_pipe14_reg_18_ ( .D(n4769), .CK(clk), .SN(rst_n), .QN(
        U1_pipe14[18]) );
  DFFSX1 U1_pipe14_reg_17_ ( .D(n4768), .CK(clk), .SN(rst_n), .QN(
        U1_pipe14[17]) );
  DFFSX1 U1_pipe14_reg_16_ ( .D(n4767), .CK(clk), .SN(rst_n), .QN(
        U1_pipe14[16]) );
  DFFSX1 U1_pipe14_reg_15_ ( .D(n4766), .CK(clk), .SN(rst_n), .QN(
        U1_pipe14[15]) );
  DFFSX1 U1_pipe14_reg_14_ ( .D(n4765), .CK(clk), .SN(rst_n), .QN(
        U1_pipe14[14]) );
  DFFSX1 U1_pipe14_reg_13_ ( .D(n4764), .CK(clk), .SN(rst_n), .QN(
        U1_pipe14[13]) );
  DFFSX1 U1_pipe14_reg_12_ ( .D(n4763), .CK(clk), .SN(rst_n), .QN(
        U1_pipe14[12]) );
  DFFSX1 U1_pipe14_reg_11_ ( .D(n4762), .CK(clk), .SN(rst_n), .QN(
        U1_pipe14[11]) );
  DFFSX1 U1_pipe14_reg_10_ ( .D(n4761), .CK(clk), .SN(rst_n), .QN(
        U1_pipe14[10]) );
  DFFSX1 U1_pipe14_reg_9_ ( .D(n4760), .CK(clk), .SN(rst_n), .QN(U1_pipe14[9])
         );
  DFFSX1 U1_pipe14_reg_8_ ( .D(n4759), .CK(clk), .SN(rst_n), .QN(U1_pipe14[8])
         );
  DFFSX1 U1_pipe14_reg_7_ ( .D(n4758), .CK(clk), .SN(rst_n), .QN(U1_pipe14[7])
         );
  DFFSX1 U1_pipe14_reg_6_ ( .D(n4757), .CK(clk), .SN(rst_n), .QN(U1_pipe14[6])
         );
  DFFSX1 U1_pipe14_reg_5_ ( .D(n4756), .CK(clk), .SN(rst_n), .QN(U1_pipe14[5])
         );
  DFFSX1 U1_pipe14_reg_4_ ( .D(n4755), .CK(clk), .SN(rst_n), .QN(U1_pipe14[4])
         );
  DFFSX1 U1_pipe14_reg_3_ ( .D(n4754), .CK(clk), .SN(rst_n), .QN(U1_pipe14[3])
         );
  DFFSX1 U1_pipe14_reg_2_ ( .D(n4753), .CK(clk), .SN(rst_n), .QN(U1_pipe14[2])
         );
  DFFSX1 U1_pipe14_reg_1_ ( .D(n4752), .CK(clk), .SN(rst_n), .QN(U1_pipe14[1])
         );
  DFFSX1 U1_pipe14_reg_0_ ( .D(n4751), .CK(clk), .SN(rst_n), .QN(U1_pipe14[0])
         );
  DFFSX1 U1_pipe13_reg_27_ ( .D(n4750), .CK(clk), .SN(rst_n), .QN(
        U1_pipe13[27]) );
  DFFSX1 U1_pipe13_reg_25_ ( .D(n4748), .CK(clk), .SN(rst_n), .Q(n28947), .QN(
        U1_pipe13[25]) );
  DFFSX1 U1_pipe13_reg_21_ ( .D(n4744), .CK(clk), .SN(rst_n), .Q(n28856), .QN(
        U1_pipe13[21]) );
  DFFSX1 U1_pipe13_reg_20_ ( .D(n4743), .CK(clk), .SN(rst_n), .Q(n28857), .QN(
        U1_pipe13[20]) );
  DFFSX1 U1_pipe13_reg_19_ ( .D(n4742), .CK(clk), .SN(rst_n), .Q(n28858), .QN(
        U1_pipe13[19]) );
  DFFSX1 U1_pipe13_reg_18_ ( .D(n4741), .CK(clk), .SN(rst_n), .Q(n28859), .QN(
        U1_pipe13[18]) );
  DFFSX1 U1_pipe13_reg_17_ ( .D(n4740), .CK(clk), .SN(rst_n), .Q(n28860), .QN(
        U1_pipe13[17]) );
  DFFSX1 U1_pipe13_reg_16_ ( .D(n4739), .CK(clk), .SN(rst_n), .Q(n28861), .QN(
        U1_pipe13[16]) );
  DFFSX1 U1_pipe13_reg_15_ ( .D(n4738), .CK(clk), .SN(rst_n), .Q(n28862), .QN(
        U1_pipe13[15]) );
  DFFSX1 U1_pipe13_reg_14_ ( .D(n4737), .CK(clk), .SN(rst_n), .Q(n28863), .QN(
        U1_pipe13[14]) );
  DFFSX1 U1_pipe13_reg_13_ ( .D(n4736), .CK(clk), .SN(rst_n), .Q(n28864), .QN(
        U1_pipe13[13]) );
  DFFSX1 U1_pipe13_reg_12_ ( .D(n4735), .CK(clk), .SN(rst_n), .Q(n28865), .QN(
        U1_pipe13[12]) );
  DFFSX1 U1_pipe13_reg_11_ ( .D(n4734), .CK(clk), .SN(rst_n), .Q(n28866), .QN(
        U1_pipe13[11]) );
  DFFSX1 U1_pipe13_reg_10_ ( .D(n4733), .CK(clk), .SN(rst_n), .Q(n28867), .QN(
        U1_pipe13[10]) );
  DFFSX1 U1_pipe13_reg_9_ ( .D(n4732), .CK(clk), .SN(rst_n), .Q(n28737), .QN(
        U1_pipe13[9]) );
  DFFSX1 U1_pipe13_reg_8_ ( .D(n4731), .CK(clk), .SN(rst_n), .Q(n28868), .QN(
        U1_pipe13[8]) );
  DFFSX1 U1_pipe13_reg_7_ ( .D(n4730), .CK(clk), .SN(rst_n), .Q(n28869), .QN(
        U1_pipe13[7]) );
  DFFSX1 U1_pipe13_reg_6_ ( .D(n4729), .CK(clk), .SN(rst_n), .Q(n28738), .QN(
        U1_pipe13[6]) );
  DFFSX1 U1_pipe13_reg_5_ ( .D(n4728), .CK(clk), .SN(rst_n), .Q(n28870), .QN(
        U1_pipe13[5]) );
  DFFSX1 U1_pipe13_reg_4_ ( .D(n4727), .CK(clk), .SN(rst_n), .Q(n28871), .QN(
        U1_pipe13[4]) );
  DFFSX1 U1_pipe13_reg_3_ ( .D(n4726), .CK(clk), .SN(rst_n), .Q(n28739), .QN(
        U1_pipe13[3]) );
  DFFSX1 U1_pipe13_reg_2_ ( .D(n4725), .CK(clk), .SN(rst_n), .Q(n28740), .QN(
        U1_pipe13[2]) );
  DFFSX1 U1_pipe13_reg_1_ ( .D(n4724), .CK(clk), .SN(rst_n), .Q(n28902), .QN(
        U1_pipe13[1]) );
  DFFSX1 U1_pipe13_reg_0_ ( .D(n4723), .CK(clk), .SN(rst_n), .Q(n28910), .QN(
        U1_pipe13[0]) );
  DFFSX1 U1_pipe12_reg_26_ ( .D(n4721), .CK(clk), .SN(rst_n), .QN(
        U1_pipe12[26]) );
  DFFSX1 U1_pipe12_reg_25_ ( .D(n4720), .CK(clk), .SN(rst_n), .QN(
        U1_pipe12[25]) );
  DFFSX1 U1_pipe12_reg_24_ ( .D(n4719), .CK(clk), .SN(rst_n), .QN(
        U1_pipe12[24]) );
  DFFSX1 U1_pipe12_reg_23_ ( .D(n4718), .CK(clk), .SN(rst_n), .QN(
        U1_pipe12[23]) );
  DFFSX1 U1_pipe12_reg_22_ ( .D(n4717), .CK(clk), .SN(rst_n), .QN(
        U1_pipe12[22]) );
  DFFSX1 U1_pipe12_reg_21_ ( .D(n4716), .CK(clk), .SN(rst_n), .QN(
        U1_pipe12[21]) );
  DFFSX1 U1_pipe12_reg_20_ ( .D(n4715), .CK(clk), .SN(rst_n), .QN(
        U1_pipe12[20]) );
  DFFSX1 U1_pipe12_reg_19_ ( .D(n4714), .CK(clk), .SN(rst_n), .QN(
        U1_pipe12[19]) );
  DFFSX1 U1_pipe12_reg_18_ ( .D(n4713), .CK(clk), .SN(rst_n), .QN(
        U1_pipe12[18]) );
  DFFSX1 U1_pipe12_reg_17_ ( .D(n4712), .CK(clk), .SN(rst_n), .QN(
        U1_pipe12[17]) );
  DFFSX1 U1_pipe12_reg_16_ ( .D(n4711), .CK(clk), .SN(rst_n), .QN(
        U1_pipe12[16]) );
  DFFSX1 U1_pipe12_reg_15_ ( .D(n4710), .CK(clk), .SN(rst_n), .QN(
        U1_pipe12[15]) );
  DFFSX1 U1_pipe12_reg_14_ ( .D(n4709), .CK(clk), .SN(rst_n), .QN(
        U1_pipe12[14]) );
  DFFSX1 U1_pipe12_reg_13_ ( .D(n4708), .CK(clk), .SN(rst_n), .QN(
        U1_pipe12[13]) );
  DFFSX1 U0_pipe12_reg_13_ ( .D(n4707), .CK(clk), .SN(rst_n), .QN(
        U0_pipe12[13]) );
  DFFSX1 U0_pipe12_reg_14_ ( .D(n4706), .CK(clk), .SN(rst_n), .QN(
        U0_pipe12[14]) );
  DFFSX1 U0_pipe12_reg_15_ ( .D(n4705), .CK(clk), .SN(rst_n), .QN(
        U0_pipe12[15]) );
  DFFSX1 U0_pipe12_reg_16_ ( .D(n4704), .CK(clk), .SN(rst_n), .QN(
        U0_pipe12[16]) );
  DFFSX1 U0_pipe12_reg_17_ ( .D(n4703), .CK(clk), .SN(rst_n), .QN(
        U0_pipe12[17]) );
  DFFSX1 U0_pipe12_reg_18_ ( .D(n4702), .CK(clk), .SN(rst_n), .QN(
        U0_pipe12[18]) );
  DFFSX1 U0_pipe12_reg_19_ ( .D(n4701), .CK(clk), .SN(rst_n), .QN(
        U0_pipe12[19]) );
  DFFSX1 U0_pipe12_reg_20_ ( .D(n4700), .CK(clk), .SN(rst_n), .QN(
        U0_pipe12[20]) );
  DFFSX1 U0_pipe12_reg_21_ ( .D(n4699), .CK(clk), .SN(rst_n), .QN(
        U0_pipe12[21]) );
  DFFSX1 U0_pipe12_reg_22_ ( .D(n4698), .CK(clk), .SN(rst_n), .QN(
        U0_pipe12[22]) );
  DFFSX1 U0_pipe12_reg_23_ ( .D(n4697), .CK(clk), .SN(rst_n), .QN(
        U0_pipe12[23]) );
  DFFSX1 U0_pipe12_reg_24_ ( .D(n4696), .CK(clk), .SN(rst_n), .QN(
        U0_pipe12[24]) );
  DFFSX1 U0_pipe12_reg_25_ ( .D(n4695), .CK(clk), .SN(rst_n), .QN(
        U0_pipe12[25]) );
  DFFSX1 U0_pipe12_reg_26_ ( .D(n4694), .CK(clk), .SN(rst_n), .QN(
        U0_pipe12[26]) );
  DFFSX1 U0_pipe13_reg_0_ ( .D(n4692), .CK(clk), .SN(rst_n), .Q(n28906), .QN(
        U0_pipe13[0]) );
  DFFSX1 U0_pipe13_reg_1_ ( .D(n4691), .CK(clk), .SN(rst_n), .Q(n28898), .QN(
        U0_pipe13[1]) );
  DFFSX1 U0_pipe13_reg_2_ ( .D(n4690), .CK(clk), .SN(rst_n), .Q(n28745), .QN(
        U0_pipe13[2]) );
  DFFSX1 U0_pipe13_reg_3_ ( .D(n4689), .CK(clk), .SN(rst_n), .Q(n28724), .QN(
        U0_pipe13[3]) );
  DFFSX1 U0_pipe13_reg_4_ ( .D(n4688), .CK(clk), .SN(rst_n), .Q(n28807), .QN(
        U0_pipe13[4]) );
  DFFSX1 U0_pipe13_reg_5_ ( .D(n4687), .CK(clk), .SN(rst_n), .Q(n28806), .QN(
        U0_pipe13[5]) );
  DFFSX1 U0_pipe13_reg_6_ ( .D(n4686), .CK(clk), .SN(rst_n), .Q(n28723), .QN(
        U0_pipe13[6]) );
  DFFSX1 U0_pipe13_reg_7_ ( .D(n4685), .CK(clk), .SN(rst_n), .Q(n28805), .QN(
        U0_pipe13[7]) );
  DFFSX1 U0_pipe13_reg_8_ ( .D(n4684), .CK(clk), .SN(rst_n), .Q(n28804), .QN(
        U0_pipe13[8]) );
  DFFSX1 U0_pipe13_reg_9_ ( .D(n4683), .CK(clk), .SN(rst_n), .Q(n28722), .QN(
        U0_pipe13[9]) );
  DFFSX1 U0_pipe13_reg_10_ ( .D(n4682), .CK(clk), .SN(rst_n), .Q(n28803), .QN(
        U0_pipe13[10]) );
  DFFSX1 U0_pipe13_reg_11_ ( .D(n4681), .CK(clk), .SN(rst_n), .Q(n28802), .QN(
        U0_pipe13[11]) );
  DFFSX1 U0_pipe13_reg_12_ ( .D(n4680), .CK(clk), .SN(rst_n), .Q(n28801), .QN(
        U0_pipe13[12]) );
  DFFSX1 U0_pipe13_reg_13_ ( .D(n4679), .CK(clk), .SN(rst_n), .Q(n28800), .QN(
        U0_pipe13[13]) );
  DFFSX1 U0_pipe13_reg_14_ ( .D(n4678), .CK(clk), .SN(rst_n), .Q(n28799), .QN(
        U0_pipe13[14]) );
  DFFSX1 U0_pipe13_reg_15_ ( .D(n4677), .CK(clk), .SN(rst_n), .Q(n28798), .QN(
        U0_pipe13[15]) );
  DFFSX1 U0_pipe13_reg_16_ ( .D(n4676), .CK(clk), .SN(rst_n), .Q(n28797), .QN(
        U0_pipe13[16]) );
  DFFSX1 U0_pipe13_reg_17_ ( .D(n4675), .CK(clk), .SN(rst_n), .Q(n28796), .QN(
        U0_pipe13[17]) );
  DFFSX1 U0_pipe13_reg_19_ ( .D(n4673), .CK(clk), .SN(rst_n), .Q(n28794), .QN(
        U0_pipe13[19]) );
  DFFSX1 U0_pipe13_reg_21_ ( .D(n4671), .CK(clk), .SN(rst_n), .Q(n28792), .QN(
        U0_pipe13[21]) );
  DFFSX1 U0_pipe13_reg_25_ ( .D(n4667), .CK(clk), .SN(rst_n), .Q(n28931), .QN(
        U0_pipe13[25]) );
  DFFSX1 U0_pipe13_reg_27_ ( .D(n4665), .CK(clk), .SN(rst_n), .QN(
        U0_pipe13[27]) );
  DFFSX1 U0_pipe14_reg_0_ ( .D(n4664), .CK(clk), .SN(rst_n), .QN(U0_pipe14[0])
         );
  DFFSX1 U0_pipe14_reg_1_ ( .D(n4663), .CK(clk), .SN(rst_n), .QN(U0_pipe14[1])
         );
  DFFSX1 U0_pipe14_reg_2_ ( .D(n4662), .CK(clk), .SN(rst_n), .QN(U0_pipe14[2])
         );
  DFFSX1 U0_pipe14_reg_3_ ( .D(n4661), .CK(clk), .SN(rst_n), .QN(U0_pipe14[3])
         );
  DFFSX1 U0_pipe14_reg_4_ ( .D(n4660), .CK(clk), .SN(rst_n), .QN(U0_pipe14[4])
         );
  DFFSX1 U0_pipe14_reg_5_ ( .D(n4659), .CK(clk), .SN(rst_n), .QN(U0_pipe14[5])
         );
  DFFSX1 U0_pipe14_reg_6_ ( .D(n4658), .CK(clk), .SN(rst_n), .QN(U0_pipe14[6])
         );
  DFFSX1 U0_pipe14_reg_7_ ( .D(n4657), .CK(clk), .SN(rst_n), .QN(U0_pipe14[7])
         );
  DFFSX1 U0_pipe14_reg_8_ ( .D(n4656), .CK(clk), .SN(rst_n), .QN(U0_pipe14[8])
         );
  DFFSX1 U0_pipe14_reg_9_ ( .D(n4655), .CK(clk), .SN(rst_n), .QN(U0_pipe14[9])
         );
  DFFSX1 U0_pipe14_reg_10_ ( .D(n4654), .CK(clk), .SN(rst_n), .QN(
        U0_pipe14[10]) );
  DFFSX1 U0_pipe14_reg_11_ ( .D(n4653), .CK(clk), .SN(rst_n), .QN(
        U0_pipe14[11]) );
  DFFSX1 U0_pipe14_reg_12_ ( .D(n4652), .CK(clk), .SN(rst_n), .QN(
        U0_pipe14[12]) );
  DFFSX1 U0_pipe14_reg_13_ ( .D(n4651), .CK(clk), .SN(rst_n), .QN(
        U0_pipe14[13]) );
  DFFSX1 U0_pipe14_reg_14_ ( .D(n4650), .CK(clk), .SN(rst_n), .QN(
        U0_pipe14[14]) );
  DFFSX1 U0_pipe14_reg_15_ ( .D(n4649), .CK(clk), .SN(rst_n), .QN(
        U0_pipe14[15]) );
  DFFSX1 U0_pipe14_reg_16_ ( .D(n4648), .CK(clk), .SN(rst_n), .QN(
        U0_pipe14[16]) );
  DFFSX1 U0_pipe14_reg_17_ ( .D(n4647), .CK(clk), .SN(rst_n), .QN(
        U0_pipe14[17]) );
  DFFSX1 U0_pipe14_reg_18_ ( .D(n4646), .CK(clk), .SN(rst_n), .QN(
        U0_pipe14[18]) );
  DFFSX1 U0_pipe14_reg_19_ ( .D(n4645), .CK(clk), .SN(rst_n), .QN(
        U0_pipe14[19]) );
  DFFSX1 U0_pipe14_reg_20_ ( .D(n4644), .CK(clk), .SN(rst_n), .QN(
        U0_pipe14[20]) );
  DFFSX1 U0_pipe14_reg_21_ ( .D(n4643), .CK(clk), .SN(rst_n), .QN(
        U0_pipe14[21]) );
  DFFSX1 U0_pipe14_reg_22_ ( .D(n4642), .CK(clk), .SN(rst_n), .QN(
        U0_pipe14[22]) );
  DFFSX1 U0_pipe14_reg_23_ ( .D(n4641), .CK(clk), .SN(rst_n), .QN(
        U0_pipe14[23]) );
  DFFSX1 U0_pipe14_reg_24_ ( .D(n4640), .CK(clk), .SN(rst_n), .QN(
        U0_pipe14[24]) );
  DFFSX1 U0_pipe14_reg_25_ ( .D(n4639), .CK(clk), .SN(rst_n), .QN(
        U0_pipe14[25]) );
  DFFSX1 U0_pipe14_reg_26_ ( .D(n4638), .CK(clk), .SN(rst_n), .QN(
        U0_pipe14[26]) );
  DFFSX1 U0_pipe15_reg_0_ ( .D(n4636), .CK(clk), .SN(rst_n), .Q(n28907), .QN(
        U0_pipe15[0]) );
  DFFSX1 U0_pipe15_reg_1_ ( .D(n4635), .CK(clk), .SN(rst_n), .Q(n28899), .QN(
        U0_pipe15[1]) );
  DFFSX1 U0_pipe15_reg_2_ ( .D(n4634), .CK(clk), .SN(rst_n), .Q(n28728), .QN(
        U0_pipe15[2]) );
  DFFSX1 U0_pipe15_reg_3_ ( .D(n4633), .CK(clk), .SN(rst_n), .Q(n28727), .QN(
        U0_pipe15[3]) );
  DFFSX1 U0_pipe15_reg_4_ ( .D(n4632), .CK(clk), .SN(rst_n), .Q(n28823), .QN(
        U0_pipe15[4]) );
  DFFSX1 U0_pipe15_reg_5_ ( .D(n4631), .CK(clk), .SN(rst_n), .Q(n28822), .QN(
        U0_pipe15[5]) );
  DFFSX1 U0_pipe15_reg_6_ ( .D(n4630), .CK(clk), .SN(rst_n), .Q(n28726), .QN(
        U0_pipe15[6]) );
  DFFSX1 U0_pipe15_reg_7_ ( .D(n4629), .CK(clk), .SN(rst_n), .Q(n28821), .QN(
        U0_pipe15[7]) );
  DFFSX1 U0_pipe15_reg_8_ ( .D(n4628), .CK(clk), .SN(rst_n), .Q(n28820), .QN(
        U0_pipe15[8]) );
  DFFSX1 U0_pipe15_reg_9_ ( .D(n4627), .CK(clk), .SN(rst_n), .Q(n28725), .QN(
        U0_pipe15[9]) );
  DFFSX1 U0_pipe15_reg_10_ ( .D(n4626), .CK(clk), .SN(rst_n), .Q(n28819), .QN(
        U0_pipe15[10]) );
  DFFSX1 U0_pipe15_reg_11_ ( .D(n4625), .CK(clk), .SN(rst_n), .Q(n28818), .QN(
        U0_pipe15[11]) );
  DFFSX1 U0_pipe15_reg_12_ ( .D(n4624), .CK(clk), .SN(rst_n), .Q(n28817), .QN(
        U0_pipe15[12]) );
  DFFSX1 U0_pipe15_reg_13_ ( .D(n4623), .CK(clk), .SN(rst_n), .Q(n28816), .QN(
        U0_pipe15[13]) );
  DFFSX1 U0_pipe15_reg_14_ ( .D(n4622), .CK(clk), .SN(rst_n), .Q(n28815), .QN(
        U0_pipe15[14]) );
  DFFSX1 U0_pipe15_reg_15_ ( .D(n4621), .CK(clk), .SN(rst_n), .Q(n28814), .QN(
        U0_pipe15[15]) );
  DFFSX1 U0_pipe15_reg_16_ ( .D(n4620), .CK(clk), .SN(rst_n), .Q(n28813), .QN(
        U0_pipe15[16]) );
  DFFSX1 U0_pipe15_reg_17_ ( .D(n4619), .CK(clk), .SN(rst_n), .Q(n28812), .QN(
        U0_pipe15[17]) );
  DFFSX1 U0_pipe15_reg_18_ ( .D(n4618), .CK(clk), .SN(rst_n), .Q(n28811), .QN(
        U0_pipe15[18]) );
  DFFSX1 U0_pipe15_reg_19_ ( .D(n4617), .CK(clk), .SN(rst_n), .Q(n28810), .QN(
        U0_pipe15[19]) );
  DFFSX1 U0_pipe15_reg_21_ ( .D(n4615), .CK(clk), .SN(rst_n), .Q(n28808), .QN(
        U0_pipe15[21]) );
  DFFSX1 U0_pipe15_reg_24_ ( .D(n4612), .CK(clk), .SN(rst_n), .Q(n28936), .QN(
        U0_pipe15[24]) );
  DFFSX1 U0_pipe15_reg_27_ ( .D(n4609), .CK(clk), .SN(rst_n), .QN(
        U0_pipe15[27]) );
  DFFSX1 U0_pipe0_reg_0_ ( .D(n4608), .CK(clk), .SN(rst_n), .QN(U0_pipe0[0])
         );
  DFFSX1 U0_pipe8_reg_26_ ( .D(n4607), .CK(clk), .SN(rst_n), .QN(U0_pipe8[26])
         );
  DFFSX1 U0_pipe9_reg_0_ ( .D(n4605), .CK(clk), .SN(rst_n), .Q(n28904), .QN(
        U0_pipe9[0]) );
  DFFSX1 U0_pipe9_reg_1_ ( .D(n4604), .CK(clk), .SN(rst_n), .Q(n28896), .QN(
        U0_pipe9[1]) );
  DFFSX1 U0_pipe9_reg_2_ ( .D(n4603), .CK(clk), .SN(rst_n), .Q(n28717), .QN(
        U0_pipe9[2]) );
  DFFSX1 U0_pipe9_reg_3_ ( .D(n4602), .CK(clk), .SN(rst_n), .Q(n28716), .QN(
        U0_pipe9[3]) );
  DFFSX1 U0_pipe9_reg_4_ ( .D(n4601), .CK(clk), .SN(rst_n), .Q(n28775), .QN(
        U0_pipe9[4]) );
  DFFSX1 U0_pipe9_reg_5_ ( .D(n4600), .CK(clk), .SN(rst_n), .Q(n28774), .QN(
        U0_pipe9[5]) );
  DFFSX1 U0_pipe9_reg_6_ ( .D(n4599), .CK(clk), .SN(rst_n), .Q(n28715), .QN(
        U0_pipe9[6]) );
  DFFSX1 U0_pipe9_reg_7_ ( .D(n4598), .CK(clk), .SN(rst_n), .Q(n28773), .QN(
        U0_pipe9[7]) );
  DFFSX1 U0_pipe9_reg_8_ ( .D(n4597), .CK(clk), .SN(rst_n), .Q(n28772), .QN(
        U0_pipe9[8]) );
  DFFSX1 U0_pipe9_reg_9_ ( .D(n4596), .CK(clk), .SN(rst_n), .Q(n28714), .QN(
        U0_pipe9[9]) );
  DFFSX1 U0_pipe9_reg_10_ ( .D(n4595), .CK(clk), .SN(rst_n), .Q(n28771), .QN(
        U0_pipe9[10]) );
  DFFSX1 U0_pipe9_reg_11_ ( .D(n4594), .CK(clk), .SN(rst_n), .Q(n28770), .QN(
        U0_pipe9[11]) );
  DFFSX1 U0_pipe9_reg_12_ ( .D(n4593), .CK(clk), .SN(rst_n), .Q(n28769), .QN(
        U0_pipe9[12]) );
  DFFSX1 U0_pipe9_reg_13_ ( .D(n4592), .CK(clk), .SN(rst_n), .Q(n28768), .QN(
        U0_pipe9[13]) );
  DFFSX1 U0_pipe9_reg_14_ ( .D(n4591), .CK(clk), .SN(rst_n), .Q(n28767), .QN(
        U0_pipe9[14]) );
  DFFSX1 U0_pipe9_reg_15_ ( .D(n4590), .CK(clk), .SN(rst_n), .Q(n28766), .QN(
        U0_pipe9[15]) );
  DFFSX1 U0_pipe9_reg_16_ ( .D(n4589), .CK(clk), .SN(rst_n), .Q(n28765), .QN(
        U0_pipe9[16]) );
  DFFSX1 U0_pipe9_reg_17_ ( .D(n4588), .CK(clk), .SN(rst_n), .Q(n28764), .QN(
        U0_pipe9[17]) );
  DFFSX1 U0_pipe9_reg_18_ ( .D(n4587), .CK(clk), .SN(rst_n), .Q(n28763), .QN(
        U0_pipe9[18]) );
  DFFSX1 U0_pipe9_reg_19_ ( .D(n4586), .CK(clk), .SN(rst_n), .Q(n28762), .QN(
        U0_pipe9[19]) );
  DFFSX1 U0_pipe9_reg_20_ ( .D(n4585), .CK(clk), .SN(rst_n), .Q(n28761), .QN(
        U0_pipe9[20]) );
  DFFSX1 U0_pipe9_reg_21_ ( .D(n4584), .CK(clk), .SN(rst_n), .Q(n28760), .QN(
        U0_pipe9[21]) );
  DFFSX1 U0_pipe9_reg_22_ ( .D(n4583), .CK(clk), .SN(rst_n), .Q(n28926), .QN(
        U0_pipe9[22]) );
  DFFSX1 U0_pipe9_reg_23_ ( .D(n4582), .CK(clk), .SN(rst_n), .Q(n28925), .QN(
        U0_pipe9[23]) );
  DFFSX1 U0_pipe9_reg_24_ ( .D(n4581), .CK(clk), .SN(rst_n), .Q(n28924), .QN(
        U0_pipe9[24]) );
  DFFSX1 U0_pipe9_reg_25_ ( .D(n4580), .CK(clk), .SN(rst_n), .Q(n28923), .QN(
        U0_pipe9[25]) );
  DFFSX1 U0_pipe9_reg_27_ ( .D(n4578), .CK(clk), .SN(rst_n), .QN(U0_pipe9[27])
         );
  DFFSX1 U0_pipe10_reg_0_ ( .D(n4577), .CK(clk), .SN(rst_n), .QN(U0_pipe10[0])
         );
  DFFSX1 U0_pipe10_reg_1_ ( .D(n4576), .CK(clk), .SN(rst_n), .Q(n28890), .QN(
        U0_pipe10[1]) );
  DFFSX1 U0_pipe10_reg_2_ ( .D(n4575), .CK(clk), .SN(rst_n), .QN(U0_pipe10[2])
         );
  DFFSX1 U0_pipe10_reg_3_ ( .D(n4574), .CK(clk), .SN(rst_n), .QN(U0_pipe10[3])
         );
  DFFSX1 U0_pipe10_reg_4_ ( .D(n4573), .CK(clk), .SN(rst_n), .QN(U0_pipe10[4])
         );
  DFFSX1 U0_pipe10_reg_5_ ( .D(n4572), .CK(clk), .SN(rst_n), .QN(U0_pipe10[5])
         );
  DFFSX1 U0_pipe10_reg_6_ ( .D(n4571), .CK(clk), .SN(rst_n), .QN(U0_pipe10[6])
         );
  DFFSX1 U0_pipe10_reg_7_ ( .D(n4570), .CK(clk), .SN(rst_n), .QN(U0_pipe10[7])
         );
  DFFSX1 U0_pipe10_reg_8_ ( .D(n4569), .CK(clk), .SN(rst_n), .QN(U0_pipe10[8])
         );
  DFFSX1 U0_pipe10_reg_9_ ( .D(n4568), .CK(clk), .SN(rst_n), .QN(U0_pipe10[9])
         );
  DFFSX1 U0_pipe10_reg_10_ ( .D(n4567), .CK(clk), .SN(rst_n), .QN(
        U0_pipe10[10]) );
  DFFSX1 U0_pipe10_reg_11_ ( .D(n4566), .CK(clk), .SN(rst_n), .QN(
        U0_pipe10[11]) );
  DFFSX1 U0_pipe10_reg_12_ ( .D(n4565), .CK(clk), .SN(rst_n), .QN(
        U0_pipe10[12]) );
  DFFSX1 U0_pipe10_reg_13_ ( .D(n4564), .CK(clk), .SN(rst_n), .QN(
        U0_pipe10[13]) );
  DFFSX1 U0_pipe10_reg_14_ ( .D(n4563), .CK(clk), .SN(rst_n), .QN(
        U0_pipe10[14]) );
  DFFSX1 U0_pipe10_reg_15_ ( .D(n4562), .CK(clk), .SN(rst_n), .QN(
        U0_pipe10[15]) );
  DFFSX1 U0_pipe10_reg_16_ ( .D(n4561), .CK(clk), .SN(rst_n), .QN(
        U0_pipe10[16]) );
  DFFSX1 U0_pipe10_reg_17_ ( .D(n4560), .CK(clk), .SN(rst_n), .QN(
        U0_pipe10[17]) );
  DFFSX1 U0_pipe10_reg_18_ ( .D(n4559), .CK(clk), .SN(rst_n), .QN(
        U0_pipe10[18]) );
  DFFSX1 U0_pipe10_reg_19_ ( .D(n4558), .CK(clk), .SN(rst_n), .QN(
        U0_pipe10[19]) );
  DFFSX1 U0_pipe10_reg_20_ ( .D(n4557), .CK(clk), .SN(rst_n), .QN(
        U0_pipe10[20]) );
  DFFSX1 U0_pipe10_reg_21_ ( .D(n4556), .CK(clk), .SN(rst_n), .QN(
        U0_pipe10[21]) );
  DFFSX1 U0_pipe10_reg_22_ ( .D(n4555), .CK(clk), .SN(rst_n), .QN(
        U0_pipe10[22]) );
  DFFSX1 U0_pipe10_reg_23_ ( .D(n4554), .CK(clk), .SN(rst_n), .QN(
        U0_pipe10[23]) );
  DFFSX1 U0_pipe10_reg_24_ ( .D(n4553), .CK(clk), .SN(rst_n), .QN(
        U0_pipe10[24]) );
  DFFSX1 U0_pipe10_reg_25_ ( .D(n4552), .CK(clk), .SN(rst_n), .QN(
        U0_pipe10[25]) );
  DFFSX1 U0_pipe10_reg_26_ ( .D(n4551), .CK(clk), .SN(rst_n), .QN(
        U0_pipe10[26]) );
  DFFSX1 U0_pipe11_reg_0_ ( .D(n4549), .CK(clk), .SN(rst_n), .QN(U0_pipe11[0])
         );
  DFFSX1 U0_pipe11_reg_1_ ( .D(n4548), .CK(clk), .SN(rst_n), .QN(U0_pipe11[1])
         );
  DFFSX1 U0_pipe11_reg_2_ ( .D(n4547), .CK(clk), .SN(rst_n), .QN(U0_pipe11[2])
         );
  DFFSX1 U0_pipe11_reg_3_ ( .D(n4546), .CK(clk), .SN(rst_n), .QN(U0_pipe11[3])
         );
  DFFSX1 U0_pipe11_reg_4_ ( .D(n4545), .CK(clk), .SN(rst_n), .QN(U0_pipe11[4])
         );
  DFFSX1 U0_pipe11_reg_5_ ( .D(n4544), .CK(clk), .SN(rst_n), .QN(U0_pipe11[5])
         );
  DFFSX1 U0_pipe11_reg_6_ ( .D(n4543), .CK(clk), .SN(rst_n), .QN(U0_pipe11[6])
         );
  DFFSX1 U0_pipe11_reg_7_ ( .D(n4542), .CK(clk), .SN(rst_n), .QN(U0_pipe11[7])
         );
  DFFSX1 U0_pipe11_reg_8_ ( .D(n4541), .CK(clk), .SN(rst_n), .QN(U0_pipe11[8])
         );
  DFFSX1 U0_pipe11_reg_9_ ( .D(n4540), .CK(clk), .SN(rst_n), .QN(U0_pipe11[9])
         );
  DFFSX1 U0_pipe11_reg_10_ ( .D(n4539), .CK(clk), .SN(rst_n), .QN(
        U0_pipe11[10]) );
  DFFSX1 U0_pipe11_reg_11_ ( .D(n4538), .CK(clk), .SN(rst_n), .QN(
        U0_pipe11[11]) );
  DFFSX1 U0_pipe11_reg_12_ ( .D(n4537), .CK(clk), .SN(rst_n), .QN(
        U0_pipe11[12]) );
  DFFSX1 U0_pipe11_reg_13_ ( .D(n4536), .CK(clk), .SN(rst_n), .QN(
        U0_pipe11[13]) );
  DFFSX1 U0_pipe11_reg_14_ ( .D(n4535), .CK(clk), .SN(rst_n), .QN(
        U0_pipe11[14]) );
  DFFSX1 U0_pipe11_reg_15_ ( .D(n4534), .CK(clk), .SN(rst_n), .QN(
        U0_pipe11[15]) );
  DFFSX1 U0_pipe11_reg_16_ ( .D(n4533), .CK(clk), .SN(rst_n), .QN(
        U0_pipe11[16]) );
  DFFSX1 U0_pipe11_reg_17_ ( .D(n4532), .CK(clk), .SN(rst_n), .QN(
        U0_pipe11[17]) );
  DFFSX1 U0_pipe11_reg_18_ ( .D(n4531), .CK(clk), .SN(rst_n), .QN(
        U0_pipe11[18]) );
  DFFSX1 U0_pipe11_reg_19_ ( .D(n4530), .CK(clk), .SN(rst_n), .QN(
        U0_pipe11[19]) );
  DFFSX1 U0_pipe11_reg_20_ ( .D(n4529), .CK(clk), .SN(rst_n), .QN(
        U0_pipe11[20]) );
  DFFSX1 U0_pipe11_reg_21_ ( .D(n4528), .CK(clk), .SN(rst_n), .QN(
        U0_pipe11[21]) );
  DFFSX1 U0_pipe11_reg_22_ ( .D(n4527), .CK(clk), .SN(rst_n), .QN(
        U0_pipe11[22]) );
  DFFSX1 U0_pipe11_reg_23_ ( .D(n4526), .CK(clk), .SN(rst_n), .QN(
        U0_pipe11[23]) );
  DFFSX1 U0_pipe11_reg_24_ ( .D(n4525), .CK(clk), .SN(rst_n), .QN(
        U0_pipe11[24]) );
  DFFSX1 U0_pipe11_reg_25_ ( .D(n4524), .CK(clk), .SN(rst_n), .QN(
        U0_pipe11[25]) );
  DFFSX1 U0_pipe11_reg_26_ ( .D(n4523), .CK(clk), .SN(rst_n), .QN(
        U0_pipe11[26]) );
  DFFSX1 U0_pipe12_reg_0_ ( .D(n4521), .CK(clk), .SN(rst_n), .QN(U0_pipe12[0])
         );
  DFFSX1 U0_pipe12_reg_1_ ( .D(n4520), .CK(clk), .SN(rst_n), .QN(U0_pipe12[1])
         );
  DFFSX1 U0_pipe12_reg_2_ ( .D(n4519), .CK(clk), .SN(rst_n), .QN(U0_pipe12[2])
         );
  DFFSX1 U0_pipe12_reg_3_ ( .D(n4518), .CK(clk), .SN(rst_n), .QN(U0_pipe12[3])
         );
  DFFSX1 U0_pipe12_reg_4_ ( .D(n4517), .CK(clk), .SN(rst_n), .QN(U0_pipe12[4])
         );
  DFFSX1 U0_pipe12_reg_5_ ( .D(n4516), .CK(clk), .SN(rst_n), .QN(U0_pipe12[5])
         );
  DFFSX1 U0_pipe12_reg_6_ ( .D(n4515), .CK(clk), .SN(rst_n), .QN(U0_pipe12[6])
         );
  DFFSX1 U0_pipe12_reg_7_ ( .D(n4514), .CK(clk), .SN(rst_n), .QN(U0_pipe12[7])
         );
  DFFSX1 U0_pipe12_reg_8_ ( .D(n4513), .CK(clk), .SN(rst_n), .QN(U0_pipe12[8])
         );
  DFFSX1 U0_pipe12_reg_9_ ( .D(n4512), .CK(clk), .SN(rst_n), .QN(U0_pipe12[9])
         );
  DFFSX1 U0_pipe12_reg_10_ ( .D(n4511), .CK(clk), .SN(rst_n), .QN(
        U0_pipe12[10]) );
  DFFSX1 U0_pipe12_reg_11_ ( .D(n4510), .CK(clk), .SN(rst_n), .QN(
        U0_pipe12[11]) );
  DFFSX1 U0_pipe12_reg_12_ ( .D(n4509), .CK(clk), .SN(rst_n), .QN(
        U0_pipe12[12]) );
  DFFSX1 U0_pipe0_reg_1_ ( .D(n4508), .CK(clk), .SN(rst_n), .Q(n28888), .QN(
        U0_pipe0[1]) );
  DFFSX1 U0_pipe5_reg_11_ ( .D(n4507), .CK(clk), .SN(rst_n), .QN(U0_pipe5[11])
         );
  DFFSX1 U0_pipe5_reg_12_ ( .D(n4506), .CK(clk), .SN(rst_n), .QN(U0_pipe5[12])
         );
  DFFSX1 U0_pipe5_reg_13_ ( .D(n4505), .CK(clk), .SN(rst_n), .QN(U0_pipe5[13])
         );
  DFFSX1 U0_pipe5_reg_14_ ( .D(n4504), .CK(clk), .SN(rst_n), .QN(U0_pipe5[14])
         );
  DFFSX1 U0_pipe5_reg_15_ ( .D(n4503), .CK(clk), .SN(rst_n), .QN(U0_pipe5[15])
         );
  DFFSX1 U0_pipe5_reg_16_ ( .D(n4502), .CK(clk), .SN(rst_n), .QN(U0_pipe5[16])
         );
  DFFSX1 U0_pipe5_reg_17_ ( .D(n4501), .CK(clk), .SN(rst_n), .QN(U0_pipe5[17])
         );
  DFFSX1 U0_pipe5_reg_18_ ( .D(n4500), .CK(clk), .SN(rst_n), .QN(U0_pipe5[18])
         );
  DFFSX1 U0_pipe5_reg_19_ ( .D(n4499), .CK(clk), .SN(rst_n), .QN(U0_pipe5[19])
         );
  DFFSX1 U0_pipe5_reg_20_ ( .D(n4498), .CK(clk), .SN(rst_n), .QN(U0_pipe5[20])
         );
  DFFSX1 U0_pipe5_reg_21_ ( .D(n4497), .CK(clk), .SN(rst_n), .QN(U0_pipe5[21])
         );
  DFFSX1 U0_pipe5_reg_22_ ( .D(n4496), .CK(clk), .SN(rst_n), .QN(U0_pipe5[22])
         );
  DFFSX1 U0_pipe5_reg_23_ ( .D(n4495), .CK(clk), .SN(rst_n), .QN(U0_pipe5[23])
         );
  DFFSX1 U0_pipe5_reg_24_ ( .D(n4494), .CK(clk), .SN(rst_n), .QN(U0_pipe5[24])
         );
  DFFSX1 U0_pipe5_reg_25_ ( .D(n4493), .CK(clk), .SN(rst_n), .QN(U0_pipe5[25])
         );
  DFFSX1 U0_pipe5_reg_26_ ( .D(n4492), .CK(clk), .SN(rst_n), .QN(U0_pipe5[26])
         );
  DFFSX1 U0_pipe6_reg_0_ ( .D(n4490), .CK(clk), .SN(rst_n), .QN(U0_pipe6[0])
         );
  DFFSX1 U0_pipe6_reg_1_ ( .D(n4489), .CK(clk), .SN(rst_n), .Q(n28891), .QN(
        U0_pipe6[1]) );
  DFFSX1 U0_pipe6_reg_2_ ( .D(n4488), .CK(clk), .SN(rst_n), .QN(U0_pipe6[2])
         );
  DFFSX1 U0_pipe6_reg_3_ ( .D(n4487), .CK(clk), .SN(rst_n), .QN(U0_pipe6[3])
         );
  DFFSX1 U0_pipe6_reg_4_ ( .D(n4486), .CK(clk), .SN(rst_n), .QN(U0_pipe6[4])
         );
  DFFSX1 U0_pipe6_reg_5_ ( .D(n4485), .CK(clk), .SN(rst_n), .QN(U0_pipe6[5])
         );
  DFFSX1 U0_pipe6_reg_6_ ( .D(n4484), .CK(clk), .SN(rst_n), .QN(U0_pipe6[6])
         );
  DFFSX1 U0_pipe6_reg_7_ ( .D(n4483), .CK(clk), .SN(rst_n), .QN(U0_pipe6[7])
         );
  DFFSX1 U0_pipe6_reg_8_ ( .D(n4482), .CK(clk), .SN(rst_n), .QN(U0_pipe6[8])
         );
  DFFSX1 U0_pipe6_reg_9_ ( .D(n4481), .CK(clk), .SN(rst_n), .QN(U0_pipe6[9])
         );
  DFFSX1 U0_pipe6_reg_10_ ( .D(n4480), .CK(clk), .SN(rst_n), .QN(U0_pipe6[10])
         );
  DFFSX1 U0_pipe6_reg_11_ ( .D(n4479), .CK(clk), .SN(rst_n), .QN(U0_pipe6[11])
         );
  DFFSX1 U0_pipe6_reg_12_ ( .D(n4478), .CK(clk), .SN(rst_n), .QN(U0_pipe6[12])
         );
  DFFSX1 U0_pipe6_reg_13_ ( .D(n4477), .CK(clk), .SN(rst_n), .QN(U0_pipe6[13])
         );
  DFFSX1 U0_pipe6_reg_14_ ( .D(n4476), .CK(clk), .SN(rst_n), .QN(U0_pipe6[14])
         );
  DFFSX1 U0_pipe6_reg_15_ ( .D(n4475), .CK(clk), .SN(rst_n), .QN(U0_pipe6[15])
         );
  DFFSX1 U0_pipe6_reg_16_ ( .D(n4474), .CK(clk), .SN(rst_n), .QN(U0_pipe6[16])
         );
  DFFSX1 U0_pipe6_reg_17_ ( .D(n4473), .CK(clk), .SN(rst_n), .QN(U0_pipe6[17])
         );
  DFFSX1 U0_pipe6_reg_18_ ( .D(n4472), .CK(clk), .SN(rst_n), .QN(U0_pipe6[18])
         );
  DFFSX1 U0_pipe6_reg_19_ ( .D(n4471), .CK(clk), .SN(rst_n), .QN(U0_pipe6[19])
         );
  DFFSX1 U0_pipe6_reg_20_ ( .D(n4470), .CK(clk), .SN(rst_n), .QN(U0_pipe6[20])
         );
  DFFSX1 U0_pipe6_reg_21_ ( .D(n4469), .CK(clk), .SN(rst_n), .QN(U0_pipe6[21])
         );
  DFFSX1 U0_pipe6_reg_22_ ( .D(n4468), .CK(clk), .SN(rst_n), .QN(U0_pipe6[22])
         );
  DFFSX1 U0_pipe6_reg_23_ ( .D(n4467), .CK(clk), .SN(rst_n), .QN(U0_pipe6[23])
         );
  DFFSX1 U0_pipe6_reg_24_ ( .D(n4466), .CK(clk), .SN(rst_n), .QN(U0_pipe6[24])
         );
  DFFSX1 U0_pipe6_reg_25_ ( .D(n4465), .CK(clk), .SN(rst_n), .QN(U0_pipe6[25])
         );
  DFFSX1 U0_pipe6_reg_26_ ( .D(n4464), .CK(clk), .SN(rst_n), .QN(U0_pipe6[26])
         );
  DFFSX1 U0_pipe6_reg_27_ ( .D(n4463), .CK(clk), .SN(rst_n), .Q(n28996), .QN(
        U0_pipe6[27]) );
  DFFSX1 U0_pipe7_reg_0_ ( .D(n4462), .CK(clk), .SN(rst_n), .QN(U0_pipe7[0])
         );
  DFFSX1 U0_pipe7_reg_1_ ( .D(n4461), .CK(clk), .SN(rst_n), .QN(U0_pipe7[1])
         );
  DFFSX1 U0_pipe7_reg_2_ ( .D(n4460), .CK(clk), .SN(rst_n), .QN(U0_pipe7[2])
         );
  DFFSX1 U0_pipe7_reg_3_ ( .D(n4459), .CK(clk), .SN(rst_n), .QN(U0_pipe7[3])
         );
  DFFSX1 U0_pipe7_reg_4_ ( .D(n4458), .CK(clk), .SN(rst_n), .QN(U0_pipe7[4])
         );
  DFFSX1 U0_pipe7_reg_5_ ( .D(n4457), .CK(clk), .SN(rst_n), .QN(U0_pipe7[5])
         );
  DFFSX1 U0_pipe7_reg_6_ ( .D(n4456), .CK(clk), .SN(rst_n), .QN(U0_pipe7[6])
         );
  DFFSX1 U0_pipe7_reg_7_ ( .D(n4455), .CK(clk), .SN(rst_n), .QN(U0_pipe7[7])
         );
  DFFSX1 U0_pipe7_reg_8_ ( .D(n4454), .CK(clk), .SN(rst_n), .QN(U0_pipe7[8])
         );
  DFFSX1 U0_pipe7_reg_9_ ( .D(n4453), .CK(clk), .SN(rst_n), .QN(U0_pipe7[9])
         );
  DFFSX1 U0_pipe7_reg_10_ ( .D(n4452), .CK(clk), .SN(rst_n), .QN(U0_pipe7[10])
         );
  DFFSX1 U0_pipe7_reg_11_ ( .D(n4451), .CK(clk), .SN(rst_n), .QN(U0_pipe7[11])
         );
  DFFSX1 U0_pipe7_reg_12_ ( .D(n4450), .CK(clk), .SN(rst_n), .QN(U0_pipe7[12])
         );
  DFFSX1 U0_pipe7_reg_13_ ( .D(n4449), .CK(clk), .SN(rst_n), .QN(U0_pipe7[13])
         );
  DFFSX1 U0_pipe7_reg_14_ ( .D(n4448), .CK(clk), .SN(rst_n), .QN(U0_pipe7[14])
         );
  DFFSX1 U0_pipe7_reg_15_ ( .D(n4447), .CK(clk), .SN(rst_n), .QN(U0_pipe7[15])
         );
  DFFSX1 U0_pipe7_reg_16_ ( .D(n4446), .CK(clk), .SN(rst_n), .QN(U0_pipe7[16])
         );
  DFFSX1 U0_pipe7_reg_17_ ( .D(n4445), .CK(clk), .SN(rst_n), .QN(U0_pipe7[17])
         );
  DFFSX1 U0_pipe7_reg_18_ ( .D(n4444), .CK(clk), .SN(rst_n), .QN(U0_pipe7[18])
         );
  DFFSX1 U0_pipe7_reg_19_ ( .D(n4443), .CK(clk), .SN(rst_n), .QN(U0_pipe7[19])
         );
  DFFSX1 U0_pipe7_reg_20_ ( .D(n4442), .CK(clk), .SN(rst_n), .QN(U0_pipe7[20])
         );
  DFFSX1 U0_pipe7_reg_21_ ( .D(n4441), .CK(clk), .SN(rst_n), .QN(U0_pipe7[21])
         );
  DFFSX1 U0_pipe7_reg_22_ ( .D(n4440), .CK(clk), .SN(rst_n), .QN(U0_pipe7[22])
         );
  DFFSX1 U0_pipe7_reg_23_ ( .D(n4439), .CK(clk), .SN(rst_n), .QN(U0_pipe7[23])
         );
  DFFSX1 U0_pipe7_reg_24_ ( .D(n4438), .CK(clk), .SN(rst_n), .QN(U0_pipe7[24])
         );
  DFFSX1 U0_pipe7_reg_25_ ( .D(n4437), .CK(clk), .SN(rst_n), .QN(U0_pipe7[25])
         );
  DFFSX1 U0_pipe7_reg_26_ ( .D(n4436), .CK(clk), .SN(rst_n), .QN(U0_pipe7[26])
         );
  DFFSX1 U0_pipe8_reg_0_ ( .D(n4434), .CK(clk), .SN(rst_n), .QN(U0_pipe8[0])
         );
  DFFSX1 U0_pipe8_reg_1_ ( .D(n4433), .CK(clk), .SN(rst_n), .QN(U0_pipe8[1])
         );
  DFFSX1 U0_pipe8_reg_2_ ( .D(n4432), .CK(clk), .SN(rst_n), .QN(U0_pipe8[2])
         );
  DFFSX1 U0_pipe8_reg_3_ ( .D(n4431), .CK(clk), .SN(rst_n), .QN(U0_pipe8[3])
         );
  DFFSX1 U0_pipe8_reg_4_ ( .D(n4430), .CK(clk), .SN(rst_n), .QN(U0_pipe8[4])
         );
  DFFSX1 U0_pipe8_reg_5_ ( .D(n4429), .CK(clk), .SN(rst_n), .QN(U0_pipe8[5])
         );
  DFFSX1 U0_pipe8_reg_6_ ( .D(n4428), .CK(clk), .SN(rst_n), .QN(U0_pipe8[6])
         );
  DFFSX1 U0_pipe8_reg_7_ ( .D(n4427), .CK(clk), .SN(rst_n), .QN(U0_pipe8[7])
         );
  DFFSX1 U0_pipe8_reg_8_ ( .D(n4426), .CK(clk), .SN(rst_n), .QN(U0_pipe8[8])
         );
  DFFSX1 U0_pipe8_reg_9_ ( .D(n4425), .CK(clk), .SN(rst_n), .QN(U0_pipe8[9])
         );
  DFFSX1 U0_pipe8_reg_10_ ( .D(n4424), .CK(clk), .SN(rst_n), .QN(U0_pipe8[10])
         );
  DFFSX1 U0_pipe8_reg_11_ ( .D(n4423), .CK(clk), .SN(rst_n), .QN(U0_pipe8[11])
         );
  DFFSX1 U0_pipe8_reg_12_ ( .D(n4422), .CK(clk), .SN(rst_n), .QN(U0_pipe8[12])
         );
  DFFSX1 U0_pipe8_reg_13_ ( .D(n4421), .CK(clk), .SN(rst_n), .QN(U0_pipe8[13])
         );
  DFFSX1 U0_pipe8_reg_14_ ( .D(n4420), .CK(clk), .SN(rst_n), .QN(U0_pipe8[14])
         );
  DFFSX1 U0_pipe8_reg_15_ ( .D(n4419), .CK(clk), .SN(rst_n), .QN(U0_pipe8[15])
         );
  DFFSX1 U0_pipe8_reg_16_ ( .D(n4418), .CK(clk), .SN(rst_n), .QN(U0_pipe8[16])
         );
  DFFSX1 U0_pipe8_reg_17_ ( .D(n4417), .CK(clk), .SN(rst_n), .QN(U0_pipe8[17])
         );
  DFFSX1 U0_pipe8_reg_18_ ( .D(n4416), .CK(clk), .SN(rst_n), .QN(U0_pipe8[18])
         );
  DFFSX1 U0_pipe8_reg_19_ ( .D(n4415), .CK(clk), .SN(rst_n), .QN(U0_pipe8[19])
         );
  DFFSX1 U0_pipe8_reg_20_ ( .D(n4414), .CK(clk), .SN(rst_n), .QN(U0_pipe8[20])
         );
  DFFSX1 U0_pipe8_reg_21_ ( .D(n4413), .CK(clk), .SN(rst_n), .QN(U0_pipe8[21])
         );
  DFFSX1 U0_pipe8_reg_22_ ( .D(n4412), .CK(clk), .SN(rst_n), .QN(U0_pipe8[22])
         );
  DFFSX1 U0_pipe8_reg_23_ ( .D(n4411), .CK(clk), .SN(rst_n), .QN(U0_pipe8[23])
         );
  DFFSX1 U0_pipe8_reg_24_ ( .D(n4410), .CK(clk), .SN(rst_n), .QN(U0_pipe8[24])
         );
  DFFSX1 U0_pipe8_reg_25_ ( .D(n4409), .CK(clk), .SN(rst_n), .QN(U0_pipe8[25])
         );
  DFFSX1 U0_pipe0_reg_2_ ( .D(n4408), .CK(clk), .SN(rst_n), .QN(U0_pipe0[2])
         );
  DFFSX1 U0_pipe1_reg_24_ ( .D(n4407), .CK(clk), .SN(rst_n), .QN(U0_pipe1[24])
         );
  DFFSX1 U0_pipe1_reg_25_ ( .D(n4406), .CK(clk), .SN(rst_n), .QN(U0_pipe1[25])
         );
  DFFSX1 U0_pipe1_reg_26_ ( .D(n4405), .CK(clk), .SN(rst_n), .QN(U0_pipe1[26])
         );
  DFFSX1 U0_pipe2_reg_0_ ( .D(n4403), .CK(clk), .SN(rst_n), .QN(U0_pipe2[0])
         );
  DFFSX1 U0_pipe2_reg_1_ ( .D(n4402), .CK(clk), .SN(rst_n), .QN(U0_pipe2[1])
         );
  DFFSX1 U0_pipe2_reg_2_ ( .D(n4401), .CK(clk), .SN(rst_n), .QN(U0_pipe2[2])
         );
  DFFSX1 U0_pipe2_reg_3_ ( .D(n4400), .CK(clk), .SN(rst_n), .QN(U0_pipe2[3])
         );
  DFFSX1 U0_pipe2_reg_4_ ( .D(n4399), .CK(clk), .SN(rst_n), .QN(U0_pipe2[4])
         );
  DFFSX1 U0_pipe2_reg_5_ ( .D(n4398), .CK(clk), .SN(rst_n), .QN(U0_pipe2[5])
         );
  DFFSX1 U0_pipe2_reg_6_ ( .D(n4397), .CK(clk), .SN(rst_n), .QN(U0_pipe2[6])
         );
  DFFSX1 U0_pipe2_reg_7_ ( .D(n4396), .CK(clk), .SN(rst_n), .QN(U0_pipe2[7])
         );
  DFFSX1 U0_pipe2_reg_8_ ( .D(n4395), .CK(clk), .SN(rst_n), .QN(U0_pipe2[8])
         );
  DFFSX1 U0_pipe2_reg_9_ ( .D(n4394), .CK(clk), .SN(rst_n), .QN(U0_pipe2[9])
         );
  DFFSX1 U0_pipe2_reg_10_ ( .D(n4393), .CK(clk), .SN(rst_n), .QN(U0_pipe2[10])
         );
  DFFSX1 U0_pipe2_reg_11_ ( .D(n4392), .CK(clk), .SN(rst_n), .QN(U0_pipe2[11])
         );
  DFFSX1 U0_pipe2_reg_12_ ( .D(n4391), .CK(clk), .SN(rst_n), .QN(U0_pipe2[12])
         );
  DFFSX1 U0_pipe2_reg_13_ ( .D(n4390), .CK(clk), .SN(rst_n), .QN(U0_pipe2[13])
         );
  DFFSX1 U0_pipe2_reg_14_ ( .D(n4389), .CK(clk), .SN(rst_n), .QN(U0_pipe2[14])
         );
  DFFSX1 U0_pipe2_reg_15_ ( .D(n4388), .CK(clk), .SN(rst_n), .QN(U0_pipe2[15])
         );
  DFFSX1 U0_pipe2_reg_16_ ( .D(n4387), .CK(clk), .SN(rst_n), .QN(U0_pipe2[16])
         );
  DFFSX1 U0_pipe2_reg_17_ ( .D(n4386), .CK(clk), .SN(rst_n), .QN(U0_pipe2[17])
         );
  DFFSX1 U0_pipe2_reg_18_ ( .D(n4385), .CK(clk), .SN(rst_n), .QN(U0_pipe2[18])
         );
  DFFSX1 U0_pipe2_reg_19_ ( .D(n4384), .CK(clk), .SN(rst_n), .QN(U0_pipe2[19])
         );
  DFFSX1 U0_pipe2_reg_20_ ( .D(n4383), .CK(clk), .SN(rst_n), .QN(U0_pipe2[20])
         );
  DFFSX1 U0_pipe2_reg_21_ ( .D(n4382), .CK(clk), .SN(rst_n), .QN(U0_pipe2[21])
         );
  DFFSX1 U0_pipe2_reg_22_ ( .D(n4381), .CK(clk), .SN(rst_n), .QN(U0_pipe2[22])
         );
  DFFSX1 U0_pipe2_reg_23_ ( .D(n4380), .CK(clk), .SN(rst_n), .QN(U0_pipe2[23])
         );
  DFFSX1 U0_pipe2_reg_24_ ( .D(n4379), .CK(clk), .SN(rst_n), .QN(U0_pipe2[24])
         );
  DFFSX1 U0_pipe2_reg_25_ ( .D(n4378), .CK(clk), .SN(rst_n), .QN(U0_pipe2[25])
         );
  DFFSX1 U0_pipe2_reg_26_ ( .D(n4377), .CK(clk), .SN(rst_n), .QN(U0_pipe2[26])
         );
  DFFSX1 U0_pipe3_reg_0_ ( .D(n4375), .CK(clk), .SN(rst_n), .Q(n28905), .QN(
        U0_pipe3[0]) );
  DFFSX1 U0_pipe3_reg_1_ ( .D(n4374), .CK(clk), .SN(rst_n), .Q(n28897), .QN(
        U0_pipe3[1]) );
  DFFSX1 U0_pipe3_reg_2_ ( .D(n4373), .CK(clk), .SN(rst_n), .Q(n28721), .QN(
        U0_pipe3[2]) );
  DFFSX1 U0_pipe3_reg_3_ ( .D(n4372), .CK(clk), .SN(rst_n), .Q(n28720), .QN(
        U0_pipe3[3]) );
  DFFSX1 U0_pipe3_reg_4_ ( .D(n4371), .CK(clk), .SN(rst_n), .Q(n28791), .QN(
        U0_pipe3[4]) );
  DFFSX1 U0_pipe3_reg_5_ ( .D(n4370), .CK(clk), .SN(rst_n), .Q(n28790), .QN(
        U0_pipe3[5]) );
  DFFSX1 U0_pipe3_reg_6_ ( .D(n4369), .CK(clk), .SN(rst_n), .Q(n28719), .QN(
        U0_pipe3[6]) );
  DFFSX1 U0_pipe3_reg_7_ ( .D(n4368), .CK(clk), .SN(rst_n), .Q(n28789), .QN(
        U0_pipe3[7]) );
  DFFSX1 U0_pipe3_reg_8_ ( .D(n4367), .CK(clk), .SN(rst_n), .Q(n28788), .QN(
        U0_pipe3[8]) );
  DFFSX1 U0_pipe3_reg_9_ ( .D(n4366), .CK(clk), .SN(rst_n), .Q(n28718), .QN(
        U0_pipe3[9]) );
  DFFSX1 U0_pipe3_reg_10_ ( .D(n4365), .CK(clk), .SN(rst_n), .Q(n28787), .QN(
        U0_pipe3[10]) );
  DFFSX1 U0_pipe3_reg_11_ ( .D(n4364), .CK(clk), .SN(rst_n), .Q(n28786), .QN(
        U0_pipe3[11]) );
  DFFSX1 U0_pipe3_reg_12_ ( .D(n4363), .CK(clk), .SN(rst_n), .Q(n28785), .QN(
        U0_pipe3[12]) );
  DFFSX1 U0_pipe3_reg_13_ ( .D(n4362), .CK(clk), .SN(rst_n), .Q(n28784), .QN(
        U0_pipe3[13]) );
  DFFSX1 U0_pipe3_reg_14_ ( .D(n4361), .CK(clk), .SN(rst_n), .Q(n28783), .QN(
        U0_pipe3[14]) );
  DFFSX1 U0_pipe3_reg_15_ ( .D(n4360), .CK(clk), .SN(rst_n), .Q(n28782), .QN(
        U0_pipe3[15]) );
  DFFSX1 U0_pipe3_reg_19_ ( .D(n4356), .CK(clk), .SN(rst_n), .Q(n28778), .QN(
        U0_pipe3[19]) );
  DFFSX1 U0_pipe3_reg_21_ ( .D(n4354), .CK(clk), .SN(rst_n), .Q(n28776), .QN(
        U0_pipe3[21]) );
  DFFSX1 U0_pipe3_reg_26_ ( .D(n4349), .CK(clk), .SN(rst_n), .Q(n29000), .QN(
        U0_pipe3[26]) );
  DFFSX1 U0_pipe3_reg_27_ ( .D(n4348), .CK(clk), .SN(rst_n), .QN(U0_pipe3[27])
         );
  DFFSX1 U0_pipe4_reg_0_ ( .D(n4347), .CK(clk), .SN(rst_n), .QN(U0_pipe4[0])
         );
  DFFSX1 U0_pipe4_reg_1_ ( .D(n4346), .CK(clk), .SN(rst_n), .Q(n28889), .QN(
        U0_pipe4[1]) );
  DFFSX1 U0_pipe4_reg_2_ ( .D(n4345), .CK(clk), .SN(rst_n), .QN(U0_pipe4[2])
         );
  DFFSX1 U0_pipe4_reg_3_ ( .D(n4344), .CK(clk), .SN(rst_n), .QN(U0_pipe4[3])
         );
  DFFSX1 U0_pipe4_reg_4_ ( .D(n4343), .CK(clk), .SN(rst_n), .QN(U0_pipe4[4])
         );
  DFFSX1 U0_pipe4_reg_5_ ( .D(n4342), .CK(clk), .SN(rst_n), .QN(U0_pipe4[5])
         );
  DFFSX1 U0_pipe4_reg_6_ ( .D(n4341), .CK(clk), .SN(rst_n), .QN(U0_pipe4[6])
         );
  DFFSX1 U0_pipe4_reg_7_ ( .D(n4340), .CK(clk), .SN(rst_n), .QN(U0_pipe4[7])
         );
  DFFSX1 U0_pipe4_reg_8_ ( .D(n4339), .CK(clk), .SN(rst_n), .QN(U0_pipe4[8])
         );
  DFFSX1 U0_pipe4_reg_9_ ( .D(n4338), .CK(clk), .SN(rst_n), .QN(U0_pipe4[9])
         );
  DFFSX1 U0_pipe4_reg_10_ ( .D(n4337), .CK(clk), .SN(rst_n), .QN(U0_pipe4[10])
         );
  DFFSX1 U0_pipe4_reg_11_ ( .D(n4336), .CK(clk), .SN(rst_n), .QN(U0_pipe4[11])
         );
  DFFSX1 U0_pipe4_reg_12_ ( .D(n4335), .CK(clk), .SN(rst_n), .QN(U0_pipe4[12])
         );
  DFFSX1 U0_pipe4_reg_13_ ( .D(n4334), .CK(clk), .SN(rst_n), .QN(U0_pipe4[13])
         );
  DFFSX1 U0_pipe4_reg_14_ ( .D(n4333), .CK(clk), .SN(rst_n), .QN(U0_pipe4[14])
         );
  DFFSX1 U0_pipe4_reg_15_ ( .D(n4332), .CK(clk), .SN(rst_n), .QN(U0_pipe4[15])
         );
  DFFSX1 U0_pipe4_reg_16_ ( .D(n4331), .CK(clk), .SN(rst_n), .QN(U0_pipe4[16])
         );
  DFFSX1 U0_pipe4_reg_17_ ( .D(n4330), .CK(clk), .SN(rst_n), .QN(U0_pipe4[17])
         );
  DFFSX1 U0_pipe4_reg_18_ ( .D(n4329), .CK(clk), .SN(rst_n), .QN(U0_pipe4[18])
         );
  DFFSX1 U0_pipe4_reg_19_ ( .D(n4328), .CK(clk), .SN(rst_n), .QN(U0_pipe4[19])
         );
  DFFSX1 U0_pipe4_reg_20_ ( .D(n4327), .CK(clk), .SN(rst_n), .QN(U0_pipe4[20])
         );
  DFFSX1 U0_pipe4_reg_21_ ( .D(n4326), .CK(clk), .SN(rst_n), .QN(U0_pipe4[21])
         );
  DFFSX1 U0_pipe4_reg_22_ ( .D(n4325), .CK(clk), .SN(rst_n), .QN(U0_pipe4[22])
         );
  DFFSX1 U0_pipe4_reg_23_ ( .D(n4324), .CK(clk), .SN(rst_n), .QN(U0_pipe4[23])
         );
  DFFSX1 U0_pipe4_reg_24_ ( .D(n4323), .CK(clk), .SN(rst_n), .QN(U0_pipe4[24])
         );
  DFFSX1 U0_pipe4_reg_25_ ( .D(n4322), .CK(clk), .SN(rst_n), .QN(U0_pipe4[25])
         );
  DFFSX1 U0_pipe4_reg_26_ ( .D(n4321), .CK(clk), .SN(rst_n), .QN(U0_pipe4[26])
         );
  DFFSX1 U0_pipe5_reg_0_ ( .D(n4319), .CK(clk), .SN(rst_n), .QN(U0_pipe5[0])
         );
  DFFSX1 U0_pipe5_reg_1_ ( .D(n4318), .CK(clk), .SN(rst_n), .QN(U0_pipe5[1])
         );
  DFFSX1 U0_pipe5_reg_2_ ( .D(n4317), .CK(clk), .SN(rst_n), .QN(U0_pipe5[2])
         );
  DFFSX1 U0_pipe5_reg_3_ ( .D(n4316), .CK(clk), .SN(rst_n), .QN(U0_pipe5[3])
         );
  DFFSX1 U0_pipe5_reg_4_ ( .D(n4315), .CK(clk), .SN(rst_n), .QN(U0_pipe5[4])
         );
  DFFSX1 U0_pipe5_reg_5_ ( .D(n4314), .CK(clk), .SN(rst_n), .QN(U0_pipe5[5])
         );
  DFFSX1 U0_pipe5_reg_6_ ( .D(n4313), .CK(clk), .SN(rst_n), .QN(U0_pipe5[6])
         );
  DFFSX1 U0_pipe5_reg_7_ ( .D(n4312), .CK(clk), .SN(rst_n), .QN(U0_pipe5[7])
         );
  DFFSX1 U0_pipe5_reg_8_ ( .D(n4311), .CK(clk), .SN(rst_n), .QN(U0_pipe5[8])
         );
  DFFSX1 U0_pipe5_reg_9_ ( .D(n4310), .CK(clk), .SN(rst_n), .QN(U0_pipe5[9])
         );
  DFFSX1 U0_pipe5_reg_10_ ( .D(n4309), .CK(clk), .SN(rst_n), .QN(U0_pipe5[10])
         );
  DFFSX1 U0_pipe0_reg_3_ ( .D(n4308), .CK(clk), .SN(rst_n), .QN(U0_pipe0[3])
         );
  DFFSX1 U0_pipe0_reg_5_ ( .D(n4307), .CK(clk), .SN(rst_n), .QN(U0_pipe0[5])
         );
  DFFSX1 U0_pipe0_reg_6_ ( .D(n4306), .CK(clk), .SN(rst_n), .QN(U0_pipe0[6])
         );
  DFFSX1 U0_pipe0_reg_7_ ( .D(n4305), .CK(clk), .SN(rst_n), .QN(U0_pipe0[7])
         );
  DFFSX1 U0_pipe0_reg_8_ ( .D(n4304), .CK(clk), .SN(rst_n), .QN(U0_pipe0[8])
         );
  DFFSX1 U0_pipe0_reg_9_ ( .D(n4303), .CK(clk), .SN(rst_n), .QN(U0_pipe0[9])
         );
  DFFSX1 U0_pipe0_reg_10_ ( .D(n4302), .CK(clk), .SN(rst_n), .QN(U0_pipe0[10])
         );
  DFFSX1 U0_pipe0_reg_11_ ( .D(n4301), .CK(clk), .SN(rst_n), .QN(U0_pipe0[11])
         );
  DFFSX1 U0_pipe0_reg_12_ ( .D(n4300), .CK(clk), .SN(rst_n), .QN(U0_pipe0[12])
         );
  DFFSX1 U0_pipe0_reg_13_ ( .D(n4299), .CK(clk), .SN(rst_n), .QN(U0_pipe0[13])
         );
  DFFSX1 U0_pipe0_reg_14_ ( .D(n4298), .CK(clk), .SN(rst_n), .QN(U0_pipe0[14])
         );
  DFFSX1 U0_pipe0_reg_15_ ( .D(n4297), .CK(clk), .SN(rst_n), .QN(U0_pipe0[15])
         );
  DFFSX1 U0_pipe0_reg_16_ ( .D(n4296), .CK(clk), .SN(rst_n), .QN(U0_pipe0[16])
         );
  DFFSX1 U0_pipe0_reg_17_ ( .D(n4295), .CK(clk), .SN(rst_n), .QN(U0_pipe0[17])
         );
  DFFSX1 U0_pipe0_reg_18_ ( .D(n4294), .CK(clk), .SN(rst_n), .QN(U0_pipe0[18])
         );
  DFFSX1 U0_pipe0_reg_19_ ( .D(n4293), .CK(clk), .SN(rst_n), .QN(U0_pipe0[19])
         );
  DFFSX1 U0_pipe0_reg_20_ ( .D(n4292), .CK(clk), .SN(rst_n), .QN(U0_pipe0[20])
         );
  DFFSX1 U0_pipe0_reg_21_ ( .D(n4291), .CK(clk), .SN(rst_n), .QN(U0_pipe0[21])
         );
  DFFSX1 U0_pipe0_reg_22_ ( .D(n4290), .CK(clk), .SN(rst_n), .QN(U0_pipe0[22])
         );
  DFFSX1 U0_pipe0_reg_23_ ( .D(n4289), .CK(clk), .SN(rst_n), .QN(U0_pipe0[23])
         );
  DFFSX1 U0_pipe0_reg_24_ ( .D(n4288), .CK(clk), .SN(rst_n), .QN(U0_pipe0[24])
         );
  DFFSX1 U0_pipe0_reg_25_ ( .D(n4287), .CK(clk), .SN(rst_n), .QN(U0_pipe0[25])
         );
  DFFSX1 U0_pipe0_reg_26_ ( .D(n4286), .CK(clk), .SN(rst_n), .QN(U0_pipe0[26])
         );
  DFFSX1 U0_pipe1_reg_0_ ( .D(n4284), .CK(clk), .SN(rst_n), .QN(U0_pipe1[0])
         );
  DFFSX1 U0_pipe1_reg_1_ ( .D(n4283), .CK(clk), .SN(rst_n), .QN(U0_pipe1[1])
         );
  DFFSX1 U0_pipe1_reg_2_ ( .D(n4282), .CK(clk), .SN(rst_n), .QN(U0_pipe1[2])
         );
  DFFSX1 U0_pipe1_reg_3_ ( .D(n4281), .CK(clk), .SN(rst_n), .QN(U0_pipe1[3])
         );
  DFFSX1 U0_pipe1_reg_4_ ( .D(n4280), .CK(clk), .SN(rst_n), .QN(U0_pipe1[4])
         );
  DFFSX1 U0_pipe1_reg_5_ ( .D(n4279), .CK(clk), .SN(rst_n), .QN(U0_pipe1[5])
         );
  DFFSX1 U0_pipe1_reg_6_ ( .D(n4278), .CK(clk), .SN(rst_n), .QN(U0_pipe1[6])
         );
  DFFSX1 U0_pipe1_reg_7_ ( .D(n4277), .CK(clk), .SN(rst_n), .QN(U0_pipe1[7])
         );
  DFFSX1 U0_pipe1_reg_8_ ( .D(n4276), .CK(clk), .SN(rst_n), .QN(U0_pipe1[8])
         );
  DFFSX1 U0_pipe1_reg_9_ ( .D(n4275), .CK(clk), .SN(rst_n), .QN(U0_pipe1[9])
         );
  DFFSX1 U0_pipe1_reg_10_ ( .D(n4274), .CK(clk), .SN(rst_n), .QN(U0_pipe1[10])
         );
  DFFSX1 U0_pipe1_reg_11_ ( .D(n4273), .CK(clk), .SN(rst_n), .QN(U0_pipe1[11])
         );
  DFFSX1 U0_pipe1_reg_12_ ( .D(n4272), .CK(clk), .SN(rst_n), .QN(U0_pipe1[12])
         );
  DFFSX1 U0_pipe1_reg_13_ ( .D(n4271), .CK(clk), .SN(rst_n), .QN(U0_pipe1[13])
         );
  DFFSX1 U0_pipe1_reg_14_ ( .D(n4270), .CK(clk), .SN(rst_n), .QN(U0_pipe1[14])
         );
  DFFSX1 U0_pipe1_reg_15_ ( .D(n4269), .CK(clk), .SN(rst_n), .QN(U0_pipe1[15])
         );
  DFFSX1 U0_pipe1_reg_16_ ( .D(n4268), .CK(clk), .SN(rst_n), .QN(U0_pipe1[16])
         );
  DFFSX1 U0_pipe1_reg_17_ ( .D(n4267), .CK(clk), .SN(rst_n), .QN(U0_pipe1[17])
         );
  DFFSX1 U0_pipe1_reg_18_ ( .D(n4266), .CK(clk), .SN(rst_n), .QN(U0_pipe1[18])
         );
  DFFSX1 U0_pipe1_reg_19_ ( .D(n4265), .CK(clk), .SN(rst_n), .QN(U0_pipe1[19])
         );
  DFFSX1 U0_pipe1_reg_20_ ( .D(n4264), .CK(clk), .SN(rst_n), .QN(U0_pipe1[20])
         );
  DFFSX1 U0_pipe1_reg_21_ ( .D(n4263), .CK(clk), .SN(rst_n), .QN(U0_pipe1[21])
         );
  DFFSX1 U0_pipe1_reg_22_ ( .D(n4262), .CK(clk), .SN(rst_n), .QN(U0_pipe1[22])
         );
  DFFSX1 U0_pipe1_reg_23_ ( .D(n4261), .CK(clk), .SN(rst_n), .QN(U0_pipe1[23])
         );
  DFFSX1 U0_pipe0_reg_4_ ( .D(n4260), .CK(clk), .SN(rst_n), .QN(U0_pipe0[4])
         );
  DFFSX1 U2_pipe0_reg_1_ ( .D(n4259), .CK(clk), .SN(rst_n), .QN(U2_pipe0[1])
         );
  DFFSX1 U2_Q0_reg_27_ ( .D(n4258), .CK(clk), .SN(rst_n), .QN(CQ0[27]) );
  DFFSX1 U2_pipe0_reg_4_ ( .D(n4257), .CK(clk), .SN(rst_n), .QN(U2_pipe0[4])
         );
  DFFSX1 U2_Q0_reg_30_ ( .D(n4256), .CK(clk), .SN(rst_n), .QN(CQ0[30]) );
  DFFSX1 U2_pipe0_reg_3_ ( .D(n4255), .CK(clk), .SN(rst_n), .QN(U2_pipe0[3])
         );
  DFFSX1 U2_Q0_reg_29_ ( .D(n4254), .CK(clk), .SN(rst_n), .QN(CQ0[29]) );
  DFFSX1 U2_pipe0_reg_2_ ( .D(n4253), .CK(clk), .SN(rst_n), .QN(U2_pipe0[2])
         );
  DFFSX1 U2_Q0_reg_28_ ( .D(n4252), .CK(clk), .SN(rst_n), .QN(CQ0[28]) );
  DFFSX1 U2_pipe0_reg_0_ ( .D(n4251), .CK(clk), .SN(rst_n), .QN(U2_pipe0[0])
         );
  DFFSX1 U2_Q0_reg_26_ ( .D(n4250), .CK(clk), .SN(rst_n), .QN(CQ0[26]) );
  DFFSX1 U2_pipe3_reg_25_ ( .D(n4249), .CK(clk), .SN(rst_n), .QN(U2_pipe3[25])
         );
  DFFSX1 U2_Q1_reg_25_ ( .D(n4248), .CK(clk), .SN(rst_n), .Q(n28969), .QN(
        CQ1[25]) );
  DFFSX1 U2_pipe3_reg_24_ ( .D(n4247), .CK(clk), .SN(rst_n), .QN(U2_pipe3[24])
         );
  DFFSX1 U2_Q1_reg_24_ ( .D(n4246), .CK(clk), .SN(rst_n), .Q(n28968), .QN(
        CQ1[24]) );
  DFFSX1 U2_pipe3_reg_23_ ( .D(n4245), .CK(clk), .SN(rst_n), .QN(U2_pipe3[23])
         );
  DFFSX1 U2_Q1_reg_23_ ( .D(n4244), .CK(clk), .SN(rst_n), .Q(n28967), .QN(
        CQ1[23]) );
  DFFSX1 U2_pipe3_reg_22_ ( .D(n4243), .CK(clk), .SN(rst_n), .QN(U2_pipe3[22])
         );
  DFFSX1 U2_Q1_reg_22_ ( .D(n4242), .CK(clk), .SN(rst_n), .Q(n28966), .QN(
        CQ1[22]) );
  DFFSX1 U2_pipe3_reg_21_ ( .D(n4241), .CK(clk), .SN(rst_n), .QN(U2_pipe3[21])
         );
  DFFSX1 U2_Q1_reg_21_ ( .D(n4240), .CK(clk), .SN(rst_n), .Q(n28965), .QN(
        CQ1[21]) );
  DFFSX1 U2_pipe3_reg_20_ ( .D(n4239), .CK(clk), .SN(rst_n), .QN(U2_pipe3[20])
         );
  DFFSX1 U2_Q1_reg_20_ ( .D(n4238), .CK(clk), .SN(rst_n), .Q(n28964), .QN(
        CQ1[20]) );
  DFFSX1 U2_pipe3_reg_19_ ( .D(n4237), .CK(clk), .SN(rst_n), .QN(U2_pipe3[19])
         );
  DFFSX1 U2_Q1_reg_19_ ( .D(n4236), .CK(clk), .SN(rst_n), .Q(n28963), .QN(
        CQ1[19]) );
  DFFSX1 U2_pipe3_reg_18_ ( .D(n4235), .CK(clk), .SN(rst_n), .QN(U2_pipe3[18])
         );
  DFFSX1 U2_Q1_reg_18_ ( .D(n4234), .CK(clk), .SN(rst_n), .Q(n28962), .QN(
        CQ1[18]) );
  DFFSX1 U2_pipe3_reg_17_ ( .D(n4233), .CK(clk), .SN(rst_n), .QN(U2_pipe3[17])
         );
  DFFSX1 U2_Q1_reg_17_ ( .D(n4232), .CK(clk), .SN(rst_n), .Q(n28961), .QN(
        CQ1[17]) );
  DFFSX1 U2_pipe3_reg_16_ ( .D(n4231), .CK(clk), .SN(rst_n), .QN(U2_pipe3[16])
         );
  DFFSX1 U2_Q1_reg_16_ ( .D(n4230), .CK(clk), .SN(rst_n), .Q(n28960), .QN(
        CQ1[16]) );
  DFFSX1 U2_pipe3_reg_15_ ( .D(n4229), .CK(clk), .SN(rst_n), .QN(U2_pipe3[15])
         );
  DFFSX1 U2_Q1_reg_15_ ( .D(n4228), .CK(clk), .SN(rst_n), .Q(n28959), .QN(
        CQ1[15]) );
  DFFSX1 U2_pipe3_reg_14_ ( .D(n4227), .CK(clk), .SN(rst_n), .QN(U2_pipe3[14])
         );
  DFFSX1 U2_Q1_reg_14_ ( .D(n4226), .CK(clk), .SN(rst_n), .Q(n28958), .QN(
        CQ1[14]) );
  DFFSX1 U2_pipe3_reg_13_ ( .D(n4225), .CK(clk), .SN(rst_n), .QN(U2_pipe3[13])
         );
  DFFSX1 U2_Q1_reg_13_ ( .D(n4224), .CK(clk), .SN(rst_n), .Q(n28957), .QN(
        CQ1[13]) );
  DFFSX1 U2_pipe3_reg_12_ ( .D(n4223), .CK(clk), .SN(rst_n), .QN(U2_pipe3[12])
         );
  DFFSX1 U2_Q1_reg_12_ ( .D(n4222), .CK(clk), .SN(rst_n), .Q(n28956), .QN(
        CQ1[12]) );
  DFFSX1 U2_pipe3_reg_11_ ( .D(n4221), .CK(clk), .SN(rst_n), .QN(U2_pipe3[11])
         );
  DFFSX1 U2_Q1_reg_11_ ( .D(n4220), .CK(clk), .SN(rst_n), .Q(n28955), .QN(
        CQ1[11]) );
  DFFSX1 U2_pipe3_reg_10_ ( .D(n4219), .CK(clk), .SN(rst_n), .QN(U2_pipe3[10])
         );
  DFFSX1 U2_Q1_reg_10_ ( .D(n4218), .CK(clk), .SN(rst_n), .QN(CQ1[10]) );
  DFFSX1 U2_pipe3_reg_9_ ( .D(n4217), .CK(clk), .SN(rst_n), .QN(U2_pipe3[9])
         );
  DFFSX1 U2_Q1_reg_9_ ( .D(n4216), .CK(clk), .SN(rst_n), .QN(CQ1[9]) );
  DFFSX1 U2_pipe3_reg_8_ ( .D(n4215), .CK(clk), .SN(rst_n), .QN(U2_pipe3[8])
         );
  DFFSX1 U2_Q1_reg_8_ ( .D(n4214), .CK(clk), .SN(rst_n), .QN(CQ1[8]) );
  DFFSX1 U2_pipe3_reg_7_ ( .D(n4213), .CK(clk), .SN(rst_n), .QN(U2_pipe3[7])
         );
  DFFSX1 U2_Q1_reg_7_ ( .D(n4212), .CK(clk), .SN(rst_n), .QN(CQ1[7]) );
  DFFSX1 U2_pipe3_reg_6_ ( .D(n4211), .CK(clk), .SN(rst_n), .QN(U2_pipe3[6])
         );
  DFFSX1 U2_Q1_reg_6_ ( .D(n4210), .CK(clk), .SN(rst_n), .QN(CQ1[6]) );
  DFFSX1 U2_pipe3_reg_5_ ( .D(n4209), .CK(clk), .SN(rst_n), .QN(U2_pipe3[5])
         );
  DFFSX1 U2_Q1_reg_5_ ( .D(n4208), .CK(clk), .SN(rst_n), .QN(CQ1[5]) );
  DFFSX1 U2_pipe3_reg_4_ ( .D(n4207), .CK(clk), .SN(rst_n), .QN(U2_pipe3[4])
         );
  DFFSX1 U2_Q1_reg_4_ ( .D(n4206), .CK(clk), .SN(rst_n), .QN(CQ1[4]) );
  DFFSX1 U2_pipe3_reg_3_ ( .D(n4205), .CK(clk), .SN(rst_n), .QN(U2_pipe3[3])
         );
  DFFSX1 U2_Q1_reg_3_ ( .D(n4204), .CK(clk), .SN(rst_n), .QN(CQ1[3]) );
  DFFSX1 U2_pipe3_reg_2_ ( .D(n4203), .CK(clk), .SN(rst_n), .QN(U2_pipe3[2])
         );
  DFFSX1 U2_Q1_reg_2_ ( .D(n4202), .CK(clk), .SN(rst_n), .QN(CQ1[2]) );
  DFFSX1 U2_pipe3_reg_1_ ( .D(n4201), .CK(clk), .SN(rst_n), .QN(U2_pipe3[1])
         );
  DFFSX1 U2_Q1_reg_1_ ( .D(n4200), .CK(clk), .SN(rst_n), .QN(CQ1[1]) );
  DFFSX1 U2_pipe3_reg_0_ ( .D(n4199), .CK(clk), .SN(rst_n), .QN(U2_pipe3[0])
         );
  DFFSX1 U2_Q1_reg_0_ ( .D(n4198), .CK(clk), .SN(rst_n), .QN(CQ1[0]) );
  DFFSX1 U2_pipe2_reg_25_ ( .D(n4197), .CK(clk), .SN(rst_n), .QN(U2_pipe2[25])
         );
  DFFSX1 U2_Q1_reg_51_ ( .D(n4196), .CK(clk), .SN(rst_n), .Q(n28984), .QN(
        CQ1[51]) );
  DFFSX1 U2_pipe2_reg_24_ ( .D(n4195), .CK(clk), .SN(rst_n), .QN(U2_pipe2[24])
         );
  DFFSX1 U2_Q1_reg_50_ ( .D(n4194), .CK(clk), .SN(rst_n), .Q(n28983), .QN(
        CQ1[50]) );
  DFFSX1 U2_pipe2_reg_23_ ( .D(n4193), .CK(clk), .SN(rst_n), .QN(U2_pipe2[23])
         );
  DFFSX1 U2_Q1_reg_49_ ( .D(n4192), .CK(clk), .SN(rst_n), .Q(n28982), .QN(
        CQ1[49]) );
  DFFSX1 U2_pipe2_reg_22_ ( .D(n4191), .CK(clk), .SN(rst_n), .QN(U2_pipe2[22])
         );
  DFFSX1 U2_Q1_reg_48_ ( .D(n4190), .CK(clk), .SN(rst_n), .Q(n28981), .QN(
        CQ1[48]) );
  DFFSX1 U2_pipe2_reg_21_ ( .D(n4189), .CK(clk), .SN(rst_n), .QN(U2_pipe2[21])
         );
  DFFSX1 U2_Q1_reg_47_ ( .D(n4188), .CK(clk), .SN(rst_n), .Q(n28980), .QN(
        CQ1[47]) );
  DFFSX1 U2_pipe2_reg_20_ ( .D(n4187), .CK(clk), .SN(rst_n), .QN(U2_pipe2[20])
         );
  DFFSX1 U2_Q1_reg_46_ ( .D(n4186), .CK(clk), .SN(rst_n), .Q(n28979), .QN(
        CQ1[46]) );
  DFFSX1 U2_pipe2_reg_19_ ( .D(n4185), .CK(clk), .SN(rst_n), .QN(U2_pipe2[19])
         );
  DFFSX1 U2_Q1_reg_45_ ( .D(n4184), .CK(clk), .SN(rst_n), .Q(n28978), .QN(
        CQ1[45]) );
  DFFSX1 U2_pipe2_reg_18_ ( .D(n4183), .CK(clk), .SN(rst_n), .QN(U2_pipe2[18])
         );
  DFFSX1 U2_Q1_reg_44_ ( .D(n4182), .CK(clk), .SN(rst_n), .Q(n28977), .QN(
        CQ1[44]) );
  DFFSX1 U2_pipe2_reg_17_ ( .D(n4181), .CK(clk), .SN(rst_n), .QN(U2_pipe2[17])
         );
  DFFSX1 U2_Q1_reg_43_ ( .D(n4180), .CK(clk), .SN(rst_n), .Q(n28976), .QN(
        CQ1[43]) );
  DFFSX1 U2_pipe2_reg_16_ ( .D(n4179), .CK(clk), .SN(rst_n), .QN(U2_pipe2[16])
         );
  DFFSX1 U2_Q1_reg_42_ ( .D(n4178), .CK(clk), .SN(rst_n), .Q(n28975), .QN(
        CQ1[42]) );
  DFFSX1 U2_pipe2_reg_15_ ( .D(n4177), .CK(clk), .SN(rst_n), .QN(U2_pipe2[15])
         );
  DFFSX1 U2_Q1_reg_41_ ( .D(n4176), .CK(clk), .SN(rst_n), .Q(n28974), .QN(
        CQ1[41]) );
  DFFSX1 U2_pipe2_reg_14_ ( .D(n4175), .CK(clk), .SN(rst_n), .QN(U2_pipe2[14])
         );
  DFFSX1 U2_Q1_reg_40_ ( .D(n4174), .CK(clk), .SN(rst_n), .Q(n28973), .QN(
        CQ1[40]) );
  DFFSX1 U2_pipe2_reg_13_ ( .D(n4173), .CK(clk), .SN(rst_n), .QN(U2_pipe2[13])
         );
  DFFSX1 U2_Q1_reg_39_ ( .D(n4172), .CK(clk), .SN(rst_n), .Q(n28972), .QN(
        CQ1[39]) );
  DFFSX1 U2_pipe2_reg_12_ ( .D(n4171), .CK(clk), .SN(rst_n), .QN(U2_pipe2[12])
         );
  DFFSX1 U2_Q1_reg_38_ ( .D(n4170), .CK(clk), .SN(rst_n), .Q(n28971), .QN(
        CQ1[38]) );
  DFFSX1 U2_pipe2_reg_11_ ( .D(n4169), .CK(clk), .SN(rst_n), .QN(U2_pipe2[11])
         );
  DFFSX1 U2_Q1_reg_37_ ( .D(n4168), .CK(clk), .SN(rst_n), .Q(n28970), .QN(
        CQ1[37]) );
  DFFSX1 U2_pipe2_reg_10_ ( .D(n4167), .CK(clk), .SN(rst_n), .QN(U2_pipe2[10])
         );
  DFFSX1 U2_Q1_reg_36_ ( .D(n4166), .CK(clk), .SN(rst_n), .QN(CQ1[36]) );
  DFFSX1 U2_pipe2_reg_9_ ( .D(n4165), .CK(clk), .SN(rst_n), .QN(U2_pipe2[9])
         );
  DFFSX1 U2_Q1_reg_35_ ( .D(n4164), .CK(clk), .SN(rst_n), .QN(CQ1[35]) );
  DFFSX1 U2_pipe2_reg_8_ ( .D(n4163), .CK(clk), .SN(rst_n), .QN(U2_pipe2[8])
         );
  DFFSX1 U2_Q1_reg_34_ ( .D(n4162), .CK(clk), .SN(rst_n), .QN(CQ1[34]) );
  DFFSX1 U2_pipe2_reg_7_ ( .D(n4161), .CK(clk), .SN(rst_n), .QN(U2_pipe2[7])
         );
  DFFSX1 U2_Q1_reg_33_ ( .D(n4160), .CK(clk), .SN(rst_n), .QN(CQ1[33]) );
  DFFSX1 U2_pipe2_reg_6_ ( .D(n4159), .CK(clk), .SN(rst_n), .QN(U2_pipe2[6])
         );
  DFFSX1 U2_Q1_reg_32_ ( .D(n4158), .CK(clk), .SN(rst_n), .QN(CQ1[32]) );
  DFFSX1 U2_pipe2_reg_5_ ( .D(n4157), .CK(clk), .SN(rst_n), .QN(U2_pipe2[5])
         );
  DFFSX1 U2_Q1_reg_31_ ( .D(n4156), .CK(clk), .SN(rst_n), .QN(CQ1[31]) );
  DFFSX1 U2_pipe2_reg_4_ ( .D(n4155), .CK(clk), .SN(rst_n), .QN(U2_pipe2[4])
         );
  DFFSX1 U2_Q1_reg_30_ ( .D(n4154), .CK(clk), .SN(rst_n), .QN(CQ1[30]) );
  DFFSX1 U2_pipe2_reg_3_ ( .D(n4153), .CK(clk), .SN(rst_n), .QN(U2_pipe2[3])
         );
  DFFSX1 U2_Q1_reg_29_ ( .D(n4152), .CK(clk), .SN(rst_n), .QN(CQ1[29]) );
  DFFSX1 U2_pipe2_reg_2_ ( .D(n4151), .CK(clk), .SN(rst_n), .QN(U2_pipe2[2])
         );
  DFFSX1 U2_Q1_reg_28_ ( .D(n4150), .CK(clk), .SN(rst_n), .QN(CQ1[28]) );
  DFFSX1 U2_pipe2_reg_1_ ( .D(n4149), .CK(clk), .SN(rst_n), .QN(U2_pipe2[1])
         );
  DFFSX1 U2_Q1_reg_27_ ( .D(n4148), .CK(clk), .SN(rst_n), .QN(CQ1[27]) );
  DFFSX1 U2_pipe2_reg_0_ ( .D(n4147), .CK(clk), .SN(rst_n), .QN(U2_pipe2[0])
         );
  DFFSX1 U2_Q1_reg_26_ ( .D(n4146), .CK(clk), .SN(rst_n), .QN(CQ1[26]) );
  DFFSX1 U2_pipe1_reg_25_ ( .D(n4145), .CK(clk), .SN(rst_n), .QN(U2_pipe1[25])
         );
  DFFSX1 U2_Q0_reg_25_ ( .D(n4144), .CK(clk), .SN(rst_n), .QN(CQ0[25]) );
  DFFSX1 U2_pipe1_reg_24_ ( .D(n4143), .CK(clk), .SN(rst_n), .QN(U2_pipe1[24])
         );
  DFFSX1 U2_Q0_reg_24_ ( .D(n4142), .CK(clk), .SN(rst_n), .QN(CQ0[24]) );
  DFFSX1 U2_pipe1_reg_23_ ( .D(n4141), .CK(clk), .SN(rst_n), .QN(U2_pipe1[23])
         );
  DFFSX1 U2_Q0_reg_23_ ( .D(n4140), .CK(clk), .SN(rst_n), .QN(CQ0[23]) );
  DFFSX1 U2_pipe1_reg_22_ ( .D(n4139), .CK(clk), .SN(rst_n), .QN(U2_pipe1[22])
         );
  DFFSX1 U2_Q0_reg_22_ ( .D(n4138), .CK(clk), .SN(rst_n), .QN(CQ0[22]) );
  DFFSX1 U2_pipe1_reg_21_ ( .D(n4137), .CK(clk), .SN(rst_n), .QN(U2_pipe1[21])
         );
  DFFSX1 U2_Q0_reg_21_ ( .D(n4136), .CK(clk), .SN(rst_n), .QN(CQ0[21]) );
  DFFSX1 U2_pipe1_reg_20_ ( .D(n4135), .CK(clk), .SN(rst_n), .QN(U2_pipe1[20])
         );
  DFFSX1 U2_Q0_reg_20_ ( .D(n4134), .CK(clk), .SN(rst_n), .QN(CQ0[20]) );
  DFFSX1 U2_pipe1_reg_19_ ( .D(n4133), .CK(clk), .SN(rst_n), .QN(U2_pipe1[19])
         );
  DFFSX1 U2_Q0_reg_19_ ( .D(n4132), .CK(clk), .SN(rst_n), .QN(CQ0[19]) );
  DFFSX1 U2_pipe1_reg_18_ ( .D(n4131), .CK(clk), .SN(rst_n), .QN(U2_pipe1[18])
         );
  DFFSX1 U2_Q0_reg_18_ ( .D(n4130), .CK(clk), .SN(rst_n), .QN(CQ0[18]) );
  DFFSX1 U2_pipe1_reg_17_ ( .D(n4129), .CK(clk), .SN(rst_n), .QN(U2_pipe1[17])
         );
  DFFSX1 U2_Q0_reg_17_ ( .D(n4128), .CK(clk), .SN(rst_n), .QN(CQ0[17]) );
  DFFSX1 U2_pipe1_reg_16_ ( .D(n4127), .CK(clk), .SN(rst_n), .QN(U2_pipe1[16])
         );
  DFFSX1 U2_Q0_reg_16_ ( .D(n4126), .CK(clk), .SN(rst_n), .QN(CQ0[16]) );
  DFFSX1 U2_pipe1_reg_15_ ( .D(n4125), .CK(clk), .SN(rst_n), .QN(U2_pipe1[15])
         );
  DFFSX1 U2_Q0_reg_15_ ( .D(n4124), .CK(clk), .SN(rst_n), .QN(CQ0[15]) );
  DFFSX1 U2_pipe1_reg_14_ ( .D(n4123), .CK(clk), .SN(rst_n), .QN(U2_pipe1[14])
         );
  DFFSX1 U2_Q0_reg_14_ ( .D(n4122), .CK(clk), .SN(rst_n), .QN(CQ0[14]) );
  DFFSX1 U2_pipe1_reg_13_ ( .D(n4121), .CK(clk), .SN(rst_n), .QN(U2_pipe1[13])
         );
  DFFSX1 U2_Q0_reg_13_ ( .D(n4120), .CK(clk), .SN(rst_n), .QN(CQ0[13]) );
  DFFSX1 U2_pipe1_reg_12_ ( .D(n4119), .CK(clk), .SN(rst_n), .QN(U2_pipe1[12])
         );
  DFFSX1 U2_Q0_reg_12_ ( .D(n4118), .CK(clk), .SN(rst_n), .QN(CQ0[12]) );
  DFFSX1 U2_pipe1_reg_11_ ( .D(n4117), .CK(clk), .SN(rst_n), .QN(U2_pipe1[11])
         );
  DFFSX1 U2_Q0_reg_11_ ( .D(n4116), .CK(clk), .SN(rst_n), .QN(CQ0[11]) );
  DFFSX1 U2_pipe1_reg_10_ ( .D(n4115), .CK(clk), .SN(rst_n), .QN(U2_pipe1[10])
         );
  DFFSX1 U2_Q0_reg_10_ ( .D(n4114), .CK(clk), .SN(rst_n), .QN(CQ0[10]) );
  DFFSX1 U2_pipe1_reg_9_ ( .D(n4113), .CK(clk), .SN(rst_n), .QN(U2_pipe1[9])
         );
  DFFSX1 U2_Q0_reg_9_ ( .D(n4112), .CK(clk), .SN(rst_n), .QN(CQ0[9]) );
  DFFSX1 U2_pipe1_reg_8_ ( .D(n4111), .CK(clk), .SN(rst_n), .QN(U2_pipe1[8])
         );
  DFFSX1 U2_Q0_reg_8_ ( .D(n4110), .CK(clk), .SN(rst_n), .QN(CQ0[8]) );
  DFFSX1 U2_pipe1_reg_7_ ( .D(n4109), .CK(clk), .SN(rst_n), .QN(U2_pipe1[7])
         );
  DFFSX1 U2_Q0_reg_7_ ( .D(n4108), .CK(clk), .SN(rst_n), .QN(CQ0[7]) );
  DFFSX1 U2_pipe1_reg_6_ ( .D(n4107), .CK(clk), .SN(rst_n), .QN(U2_pipe1[6])
         );
  DFFSX1 U2_Q0_reg_6_ ( .D(n4106), .CK(clk), .SN(rst_n), .QN(CQ0[6]) );
  DFFSX1 U2_pipe1_reg_5_ ( .D(n4105), .CK(clk), .SN(rst_n), .QN(U2_pipe1[5])
         );
  DFFSX1 U2_Q0_reg_5_ ( .D(n4104), .CK(clk), .SN(rst_n), .QN(CQ0[5]) );
  DFFSX1 U2_pipe1_reg_4_ ( .D(n4103), .CK(clk), .SN(rst_n), .QN(U2_pipe1[4])
         );
  DFFSX1 U2_Q0_reg_4_ ( .D(n4102), .CK(clk), .SN(rst_n), .QN(CQ0[4]) );
  DFFSX1 U2_pipe1_reg_3_ ( .D(n4101), .CK(clk), .SN(rst_n), .QN(U2_pipe1[3])
         );
  DFFSX1 U2_Q0_reg_3_ ( .D(n4100), .CK(clk), .SN(rst_n), .QN(CQ0[3]) );
  DFFSX1 U2_pipe1_reg_2_ ( .D(n4099), .CK(clk), .SN(rst_n), .QN(U2_pipe1[2])
         );
  DFFSX1 U2_Q0_reg_2_ ( .D(n4098), .CK(clk), .SN(rst_n), .QN(CQ0[2]) );
  DFFSX1 U2_pipe1_reg_1_ ( .D(n4097), .CK(clk), .SN(rst_n), .QN(U2_pipe1[1])
         );
  DFFSX1 U2_Q0_reg_1_ ( .D(n4096), .CK(clk), .SN(rst_n), .QN(CQ0[1]) );
  DFFSX1 U2_pipe1_reg_0_ ( .D(n4095), .CK(clk), .SN(rst_n), .QN(U2_pipe1[0])
         );
  DFFSX1 U2_Q0_reg_0_ ( .D(n4094), .CK(clk), .SN(rst_n), .QN(CQ0[0]) );
  DFFSX1 U2_pipe0_reg_25_ ( .D(n4093), .CK(clk), .SN(rst_n), .QN(U2_pipe0[25])
         );
  DFFSX1 U2_Q0_reg_51_ ( .D(n4092), .CK(clk), .SN(rst_n), .QN(CQ0[51]) );
  DFFSX1 U2_pipe0_reg_24_ ( .D(n4091), .CK(clk), .SN(rst_n), .QN(U2_pipe0[24])
         );
  DFFSX1 U2_Q0_reg_50_ ( .D(n4090), .CK(clk), .SN(rst_n), .QN(CQ0[50]) );
  DFFSX1 U2_pipe0_reg_23_ ( .D(n4089), .CK(clk), .SN(rst_n), .QN(U2_pipe0[23])
         );
  DFFSX1 U2_Q0_reg_49_ ( .D(n4088), .CK(clk), .SN(rst_n), .QN(CQ0[49]) );
  DFFSX1 U2_pipe0_reg_22_ ( .D(n4087), .CK(clk), .SN(rst_n), .QN(U2_pipe0[22])
         );
  DFFSX1 U2_Q0_reg_48_ ( .D(n4086), .CK(clk), .SN(rst_n), .QN(CQ0[48]) );
  DFFSX1 U2_pipe0_reg_21_ ( .D(n4085), .CK(clk), .SN(rst_n), .QN(U2_pipe0[21])
         );
  DFFSX1 U2_Q0_reg_47_ ( .D(n4084), .CK(clk), .SN(rst_n), .QN(CQ0[47]) );
  DFFSX1 U2_pipe0_reg_20_ ( .D(n4083), .CK(clk), .SN(rst_n), .QN(U2_pipe0[20])
         );
  DFFSX1 U2_Q0_reg_46_ ( .D(n4082), .CK(clk), .SN(rst_n), .QN(CQ0[46]) );
  DFFSX1 U2_pipe0_reg_19_ ( .D(n4081), .CK(clk), .SN(rst_n), .QN(U2_pipe0[19])
         );
  DFFSX1 U2_Q0_reg_45_ ( .D(n4080), .CK(clk), .SN(rst_n), .QN(CQ0[45]) );
  DFFSX1 U2_pipe0_reg_18_ ( .D(n4079), .CK(clk), .SN(rst_n), .QN(U2_pipe0[18])
         );
  DFFSX1 U2_Q0_reg_44_ ( .D(n4078), .CK(clk), .SN(rst_n), .QN(CQ0[44]) );
  DFFSX1 U2_pipe0_reg_17_ ( .D(n4077), .CK(clk), .SN(rst_n), .QN(U2_pipe0[17])
         );
  DFFSX1 U2_Q0_reg_43_ ( .D(n4076), .CK(clk), .SN(rst_n), .QN(CQ0[43]) );
  DFFSX1 U2_pipe0_reg_16_ ( .D(n4075), .CK(clk), .SN(rst_n), .QN(U2_pipe0[16])
         );
  DFFSX1 U2_Q0_reg_42_ ( .D(n4074), .CK(clk), .SN(rst_n), .QN(CQ0[42]) );
  DFFSX1 U2_pipe0_reg_15_ ( .D(n4073), .CK(clk), .SN(rst_n), .QN(U2_pipe0[15])
         );
  DFFSX1 U2_Q0_reg_41_ ( .D(n4072), .CK(clk), .SN(rst_n), .QN(CQ0[41]) );
  DFFSX1 U2_pipe0_reg_14_ ( .D(n4071), .CK(clk), .SN(rst_n), .QN(U2_pipe0[14])
         );
  DFFSX1 U2_Q0_reg_40_ ( .D(n4070), .CK(clk), .SN(rst_n), .QN(CQ0[40]) );
  DFFSX1 U2_pipe0_reg_13_ ( .D(n4069), .CK(clk), .SN(rst_n), .QN(U2_pipe0[13])
         );
  DFFSX1 U2_Q0_reg_39_ ( .D(n4068), .CK(clk), .SN(rst_n), .QN(CQ0[39]) );
  DFFSX1 U2_pipe0_reg_12_ ( .D(n4067), .CK(clk), .SN(rst_n), .QN(U2_pipe0[12])
         );
  DFFSX1 U2_Q0_reg_38_ ( .D(n4066), .CK(clk), .SN(rst_n), .QN(CQ0[38]) );
  DFFSX1 U2_pipe0_reg_11_ ( .D(n4065), .CK(clk), .SN(rst_n), .QN(U2_pipe0[11])
         );
  DFFSX1 U2_Q0_reg_37_ ( .D(n4064), .CK(clk), .SN(rst_n), .QN(CQ0[37]) );
  DFFSX1 U2_pipe0_reg_10_ ( .D(n4063), .CK(clk), .SN(rst_n), .QN(U2_pipe0[10])
         );
  DFFSX1 U2_Q0_reg_36_ ( .D(n4062), .CK(clk), .SN(rst_n), .QN(CQ0[36]) );
  DFFSX1 U2_pipe0_reg_9_ ( .D(n4061), .CK(clk), .SN(rst_n), .QN(U2_pipe0[9])
         );
  DFFSX1 U2_Q0_reg_35_ ( .D(n4060), .CK(clk), .SN(rst_n), .QN(CQ0[35]) );
  DFFSX1 U2_pipe0_reg_8_ ( .D(n4059), .CK(clk), .SN(rst_n), .QN(U2_pipe0[8])
         );
  DFFSX1 U2_Q0_reg_34_ ( .D(n4058), .CK(clk), .SN(rst_n), .QN(CQ0[34]) );
  DFFSX1 U2_pipe0_reg_7_ ( .D(n4057), .CK(clk), .SN(rst_n), .QN(U2_pipe0[7])
         );
  DFFSX1 U2_Q0_reg_33_ ( .D(n4056), .CK(clk), .SN(rst_n), .QN(CQ0[33]) );
  DFFSX1 U2_pipe0_reg_6_ ( .D(n4055), .CK(clk), .SN(rst_n), .QN(U2_pipe0[6])
         );
  DFFSX1 U2_Q0_reg_32_ ( .D(n4054), .CK(clk), .SN(rst_n), .QN(CQ0[32]) );
  DFFSX1 U2_pipe0_reg_5_ ( .D(n4053), .CK(clk), .SN(rst_n), .QN(U2_pipe0[5])
         );
  DFFSX1 U2_Q0_reg_31_ ( .D(n4052), .CK(clk), .SN(rst_n), .QN(CQ0[31]) );
  DFFSX1 U1_Q0_r_reg_2_ ( .D(n4051), .CK(clk), .SN(rst_n), .QN(Q4[30]) );
  DFFSX1 U1_Q0_r_reg_25_ ( .D(n4050), .CK(clk), .SN(rst_n), .QN(Q4[53]) );
  DFFSX1 U1_Q0_r_reg_24_ ( .D(n4049), .CK(clk), .SN(rst_n), .QN(Q4[52]) );
  DFFSX1 U1_Q0_r_reg_23_ ( .D(n4048), .CK(clk), .SN(rst_n), .QN(Q4[51]) );
  DFFSX1 U1_Q0_r_reg_22_ ( .D(n4047), .CK(clk), .SN(rst_n), .QN(Q4[50]) );
  DFFSX1 U1_Q0_r_reg_21_ ( .D(n4046), .CK(clk), .SN(rst_n), .QN(Q4[49]) );
  DFFSX1 U1_Q0_r_reg_20_ ( .D(n4045), .CK(clk), .SN(rst_n), .QN(Q4[48]) );
  DFFSX1 U1_Q0_r_reg_19_ ( .D(n4044), .CK(clk), .SN(rst_n), .QN(Q4[47]) );
  DFFSX1 U1_Q0_r_reg_18_ ( .D(n4043), .CK(clk), .SN(rst_n), .QN(Q4[46]) );
  DFFSX1 U1_Q0_r_reg_17_ ( .D(n4042), .CK(clk), .SN(rst_n), .QN(Q4[45]) );
  DFFSX1 U1_Q0_r_reg_16_ ( .D(n4041), .CK(clk), .SN(rst_n), .QN(Q4[44]) );
  DFFSX1 U1_Q0_r_reg_15_ ( .D(n4040), .CK(clk), .SN(rst_n), .QN(Q4[43]) );
  DFFSX1 U1_Q0_r_reg_14_ ( .D(n4039), .CK(clk), .SN(rst_n), .QN(Q4[42]) );
  DFFSX1 U1_Q0_r_reg_13_ ( .D(n4038), .CK(clk), .SN(rst_n), .QN(Q4[41]) );
  DFFSX1 U1_Q0_r_reg_12_ ( .D(n4037), .CK(clk), .SN(rst_n), .QN(Q4[40]) );
  DFFSX1 U1_Q0_r_reg_11_ ( .D(n4036), .CK(clk), .SN(rst_n), .QN(Q4[39]) );
  DFFSX1 U1_Q0_r_reg_10_ ( .D(n4035), .CK(clk), .SN(rst_n), .QN(Q4[38]) );
  DFFSX1 U1_Q0_r_reg_9_ ( .D(n4034), .CK(clk), .SN(rst_n), .QN(Q4[37]) );
  DFFSX1 U1_Q0_r_reg_8_ ( .D(n4033), .CK(clk), .SN(rst_n), .QN(Q4[36]) );
  DFFSX1 U1_Q0_r_reg_7_ ( .D(n4032), .CK(clk), .SN(rst_n), .QN(Q4[35]) );
  DFFSX1 U1_Q0_r_reg_6_ ( .D(n4031), .CK(clk), .SN(rst_n), .QN(Q4[34]) );
  DFFSX1 U1_Q0_r_reg_5_ ( .D(n4030), .CK(clk), .SN(rst_n), .QN(Q4[33]) );
  DFFSX1 U1_Q0_r_reg_4_ ( .D(n4029), .CK(clk), .SN(rst_n), .QN(Q4[32]) );
  DFFSX1 U1_Q0_r_reg_3_ ( .D(n4028), .CK(clk), .SN(rst_n), .QN(Q4[31]) );
  DFFSX1 U1_Q0_r_reg_1_ ( .D(n4027), .CK(clk), .SN(rst_n), .QN(Q4[29]) );
  DFFSX1 U1_Q2_r_reg_12_ ( .D(n4026), .CK(clk), .SN(rst_n), .QN(Q6[40]) );
  DFFSX1 U1_Q2_r_reg_11_ ( .D(n4025), .CK(clk), .SN(rst_n), .QN(Q6[39]) );
  DFFSX1 U1_Q2_r_reg_10_ ( .D(n4024), .CK(clk), .SN(rst_n), .QN(Q6[38]) );
  DFFSX1 U1_Q2_r_reg_9_ ( .D(n4023), .CK(clk), .SN(rst_n), .QN(Q6[37]) );
  DFFSX1 U1_Q2_r_reg_8_ ( .D(n4022), .CK(clk), .SN(rst_n), .QN(Q6[36]) );
  DFFSX1 U1_Q2_r_reg_7_ ( .D(n4021), .CK(clk), .SN(rst_n), .QN(Q6[35]) );
  DFFSX1 U1_Q2_r_reg_6_ ( .D(n4020), .CK(clk), .SN(rst_n), .QN(Q6[34]) );
  DFFSX1 U1_Q2_r_reg_5_ ( .D(n4019), .CK(clk), .SN(rst_n), .QN(Q6[33]) );
  DFFSX1 U1_Q2_r_reg_4_ ( .D(n4018), .CK(clk), .SN(rst_n), .QN(Q6[32]) );
  DFFSX1 U1_Q2_r_reg_3_ ( .D(n4017), .CK(clk), .SN(rst_n), .QN(Q6[31]) );
  DFFSX1 U1_Q2_r_reg_2_ ( .D(n4016), .CK(clk), .SN(rst_n), .QN(Q6[30]) );
  DFFSX1 U1_Q2_r_reg_1_ ( .D(n4015), .CK(clk), .SN(rst_n), .QN(Q6[29]) );
  DFFSX1 U1_Q2_r_reg_0_ ( .D(n4014), .CK(clk), .SN(rst_n), .QN(Q6[28]) );
  DFFSX1 U1_Q1_i_reg_25_ ( .D(n4013), .CK(clk), .SN(rst_n), .QN(Q5[25]) );
  DFFSX1 U1_Q1_i_reg_24_ ( .D(n4012), .CK(clk), .SN(rst_n), .QN(Q5[24]) );
  DFFSX1 U1_Q1_i_reg_23_ ( .D(n4011), .CK(clk), .SN(rst_n), .QN(Q5[23]) );
  DFFSX1 U1_Q1_i_reg_22_ ( .D(n4010), .CK(clk), .SN(rst_n), .QN(Q5[22]) );
  DFFSX1 U1_Q1_i_reg_21_ ( .D(n4009), .CK(clk), .SN(rst_n), .QN(Q5[21]) );
  DFFSX1 U1_Q1_i_reg_20_ ( .D(n4008), .CK(clk), .SN(rst_n), .QN(Q5[20]) );
  DFFSX1 U1_Q1_i_reg_19_ ( .D(n4007), .CK(clk), .SN(rst_n), .QN(Q5[19]) );
  DFFSX1 U1_Q1_i_reg_18_ ( .D(n4006), .CK(clk), .SN(rst_n), .QN(Q5[18]) );
  DFFSX1 U1_Q1_i_reg_17_ ( .D(n4005), .CK(clk), .SN(rst_n), .QN(Q5[17]) );
  DFFSX1 U1_Q1_i_reg_16_ ( .D(n4004), .CK(clk), .SN(rst_n), .QN(Q5[16]) );
  DFFSX1 U1_Q1_i_reg_15_ ( .D(n4003), .CK(clk), .SN(rst_n), .QN(Q5[15]) );
  DFFSX1 U1_Q1_i_reg_14_ ( .D(n4002), .CK(clk), .SN(rst_n), .QN(Q5[14]) );
  DFFSX1 U1_Q1_i_reg_13_ ( .D(n4001), .CK(clk), .SN(rst_n), .QN(Q5[13]) );
  DFFSX1 U1_Q1_i_reg_12_ ( .D(n4000), .CK(clk), .SN(rst_n), .QN(Q5[12]) );
  DFFSX1 U1_Q1_i_reg_11_ ( .D(n3999), .CK(clk), .SN(rst_n), .QN(Q5[11]) );
  DFFSX1 U1_Q1_i_reg_10_ ( .D(n3998), .CK(clk), .SN(rst_n), .QN(Q5[10]) );
  DFFSX1 U1_Q1_i_reg_9_ ( .D(n3997), .CK(clk), .SN(rst_n), .QN(Q5[9]) );
  DFFSX1 U1_Q1_i_reg_8_ ( .D(n3996), .CK(clk), .SN(rst_n), .QN(Q5[8]) );
  DFFSX1 U1_Q1_i_reg_7_ ( .D(n3995), .CK(clk), .SN(rst_n), .QN(Q5[7]) );
  DFFSX1 U1_Q1_i_reg_6_ ( .D(n3994), .CK(clk), .SN(rst_n), .QN(Q5[6]) );
  DFFSX1 U1_Q1_i_reg_5_ ( .D(n3993), .CK(clk), .SN(rst_n), .QN(Q5[5]) );
  DFFSX1 U1_Q1_i_reg_4_ ( .D(n3992), .CK(clk), .SN(rst_n), .QN(Q5[4]) );
  DFFSX1 U1_Q1_i_reg_3_ ( .D(n3991), .CK(clk), .SN(rst_n), .QN(Q5[3]) );
  DFFSX1 U1_Q1_i_reg_2_ ( .D(n3990), .CK(clk), .SN(rst_n), .QN(Q5[2]) );
  DFFSX1 U1_Q1_i_reg_1_ ( .D(n3989), .CK(clk), .SN(rst_n), .QN(Q5[1]) );
  DFFSX1 U1_Q1_i_reg_0_ ( .D(n3988), .CK(clk), .SN(rst_n), .QN(Q5[0]) );
  DFFSX1 U1_Q1_r_reg_25_ ( .D(n3987), .CK(clk), .SN(rst_n), .QN(Q5[53]) );
  DFFSX1 U1_Q1_r_reg_24_ ( .D(n3986), .CK(clk), .SN(rst_n), .QN(Q5[52]) );
  DFFSX1 U1_Q1_r_reg_23_ ( .D(n3985), .CK(clk), .SN(rst_n), .QN(Q5[51]) );
  DFFSX1 U1_Q1_r_reg_22_ ( .D(n3984), .CK(clk), .SN(rst_n), .QN(Q5[50]) );
  DFFSX1 U1_Q1_r_reg_21_ ( .D(n3983), .CK(clk), .SN(rst_n), .QN(Q5[49]) );
  DFFSX1 U1_Q1_r_reg_20_ ( .D(n3982), .CK(clk), .SN(rst_n), .QN(Q5[48]) );
  DFFSX1 U1_Q1_r_reg_19_ ( .D(n3981), .CK(clk), .SN(rst_n), .QN(Q5[47]) );
  DFFSX1 U1_Q1_r_reg_18_ ( .D(n3980), .CK(clk), .SN(rst_n), .QN(Q5[46]) );
  DFFSX1 U1_Q1_r_reg_17_ ( .D(n3979), .CK(clk), .SN(rst_n), .QN(Q5[45]) );
  DFFSX1 U1_Q1_r_reg_16_ ( .D(n3978), .CK(clk), .SN(rst_n), .QN(Q5[44]) );
  DFFSX1 U1_Q1_r_reg_15_ ( .D(n3977), .CK(clk), .SN(rst_n), .QN(Q5[43]) );
  DFFSX1 U1_Q1_r_reg_14_ ( .D(n3976), .CK(clk), .SN(rst_n), .QN(Q5[42]) );
  DFFSX1 U1_Q1_r_reg_13_ ( .D(n3975), .CK(clk), .SN(rst_n), .QN(Q5[41]) );
  DFFSX1 U1_Q1_r_reg_12_ ( .D(n3974), .CK(clk), .SN(rst_n), .QN(Q5[40]) );
  DFFSX1 U1_Q1_r_reg_11_ ( .D(n3973), .CK(clk), .SN(rst_n), .QN(Q5[39]) );
  DFFSX1 U1_Q1_r_reg_10_ ( .D(n3972), .CK(clk), .SN(rst_n), .QN(Q5[38]) );
  DFFSX1 U1_Q1_r_reg_9_ ( .D(n3971), .CK(clk), .SN(rst_n), .QN(Q5[37]) );
  DFFSX1 U1_Q1_r_reg_8_ ( .D(n3970), .CK(clk), .SN(rst_n), .QN(Q5[36]) );
  DFFSX1 U1_Q1_r_reg_7_ ( .D(n3969), .CK(clk), .SN(rst_n), .QN(Q5[35]) );
  DFFSX1 U1_Q1_r_reg_6_ ( .D(n3968), .CK(clk), .SN(rst_n), .QN(Q5[34]) );
  DFFSX1 U1_Q1_r_reg_5_ ( .D(n3967), .CK(clk), .SN(rst_n), .QN(Q5[33]) );
  DFFSX1 U1_Q1_r_reg_4_ ( .D(n3966), .CK(clk), .SN(rst_n), .QN(Q5[32]) );
  DFFSX1 U1_Q1_r_reg_3_ ( .D(n3965), .CK(clk), .SN(rst_n), .QN(Q5[31]) );
  DFFSX1 U1_Q1_r_reg_2_ ( .D(n3964), .CK(clk), .SN(rst_n), .QN(Q5[30]) );
  DFFSX1 U1_Q1_r_reg_1_ ( .D(n3963), .CK(clk), .SN(rst_n), .QN(Q5[29]) );
  DFFSX1 U1_Q1_r_reg_0_ ( .D(n3962), .CK(clk), .SN(rst_n), .QN(Q5[28]) );
  DFFSX1 U1_Q0_i_reg_25_ ( .D(n3961), .CK(clk), .SN(rst_n), .QN(Q4[25]) );
  DFFSX1 U1_Q0_i_reg_24_ ( .D(n3960), .CK(clk), .SN(rst_n), .QN(Q4[24]) );
  DFFSX1 U1_Q0_i_reg_23_ ( .D(n3959), .CK(clk), .SN(rst_n), .QN(Q4[23]) );
  DFFSX1 U1_Q0_i_reg_22_ ( .D(n3958), .CK(clk), .SN(rst_n), .QN(Q4[22]) );
  DFFSX1 U1_Q0_i_reg_21_ ( .D(n3957), .CK(clk), .SN(rst_n), .QN(Q4[21]) );
  DFFSX1 U1_Q0_i_reg_20_ ( .D(n3956), .CK(clk), .SN(rst_n), .QN(Q4[20]) );
  DFFSX1 U1_Q0_i_reg_19_ ( .D(n3955), .CK(clk), .SN(rst_n), .QN(Q4[19]) );
  DFFSX1 U1_Q0_i_reg_18_ ( .D(n3954), .CK(clk), .SN(rst_n), .QN(Q4[18]) );
  DFFSX1 U1_Q0_i_reg_17_ ( .D(n3953), .CK(clk), .SN(rst_n), .QN(Q4[17]) );
  DFFSX1 U1_Q0_i_reg_16_ ( .D(n3952), .CK(clk), .SN(rst_n), .QN(Q4[16]) );
  DFFSX1 U1_Q0_i_reg_15_ ( .D(n3951), .CK(clk), .SN(rst_n), .QN(Q4[15]) );
  DFFSX1 U1_Q0_i_reg_14_ ( .D(n3950), .CK(clk), .SN(rst_n), .QN(Q4[14]) );
  DFFSX1 U1_Q0_i_reg_13_ ( .D(n3949), .CK(clk), .SN(rst_n), .QN(Q4[13]) );
  DFFSX1 U1_Q0_i_reg_12_ ( .D(n3948), .CK(clk), .SN(rst_n), .QN(Q4[12]) );
  DFFSX1 U1_Q0_i_reg_11_ ( .D(n3947), .CK(clk), .SN(rst_n), .QN(Q4[11]) );
  DFFSX1 U1_Q0_i_reg_10_ ( .D(n3946), .CK(clk), .SN(rst_n), .QN(Q4[10]) );
  DFFSX1 U1_Q0_i_reg_9_ ( .D(n3945), .CK(clk), .SN(rst_n), .QN(Q4[9]) );
  DFFSX1 U1_Q0_i_reg_8_ ( .D(n3944), .CK(clk), .SN(rst_n), .QN(Q4[8]) );
  DFFSX1 U1_Q0_i_reg_7_ ( .D(n3943), .CK(clk), .SN(rst_n), .QN(Q4[7]) );
  DFFSX1 U1_Q0_i_reg_6_ ( .D(n3942), .CK(clk), .SN(rst_n), .QN(Q4[6]) );
  DFFSX1 U1_Q0_i_reg_5_ ( .D(n3941), .CK(clk), .SN(rst_n), .QN(Q4[5]) );
  DFFSX1 U1_Q0_i_reg_4_ ( .D(n3940), .CK(clk), .SN(rst_n), .QN(Q4[4]) );
  DFFSX1 U1_Q0_i_reg_3_ ( .D(n3939), .CK(clk), .SN(rst_n), .QN(Q4[3]) );
  DFFSX1 U1_Q0_i_reg_2_ ( .D(n3938), .CK(clk), .SN(rst_n), .QN(Q4[2]) );
  DFFSX1 U1_Q0_i_reg_1_ ( .D(n3937), .CK(clk), .SN(rst_n), .QN(Q4[1]) );
  DFFSX1 U1_Q0_i_reg_0_ ( .D(n3936), .CK(clk), .SN(rst_n), .QN(Q4[0]) );
  DFFSX1 U1_Q0_r_reg_0_ ( .D(n3935), .CK(clk), .SN(rst_n), .QN(Q4[28]) );
  DFFSX1 U1_Q3_i_reg_25_ ( .D(n3934), .CK(clk), .SN(rst_n), .QN(Q7[25]) );
  DFFSX1 U1_Q3_i_reg_24_ ( .D(n3933), .CK(clk), .SN(rst_n), .QN(Q7[24]) );
  DFFSX1 U1_Q3_i_reg_23_ ( .D(n3932), .CK(clk), .SN(rst_n), .QN(Q7[23]) );
  DFFSX1 U1_Q3_i_reg_22_ ( .D(n3931), .CK(clk), .SN(rst_n), .QN(Q7[22]) );
  DFFSX1 U1_Q3_i_reg_21_ ( .D(n3930), .CK(clk), .SN(rst_n), .QN(Q7[21]) );
  DFFSX1 U1_Q3_i_reg_20_ ( .D(n3929), .CK(clk), .SN(rst_n), .QN(Q7[20]) );
  DFFSX1 U1_Q3_i_reg_19_ ( .D(n3928), .CK(clk), .SN(rst_n), .QN(Q7[19]) );
  DFFSX1 U1_Q3_i_reg_18_ ( .D(n3927), .CK(clk), .SN(rst_n), .QN(Q7[18]) );
  DFFSX1 U1_Q3_i_reg_17_ ( .D(n3926), .CK(clk), .SN(rst_n), .QN(Q7[17]) );
  DFFSX1 U1_Q3_i_reg_16_ ( .D(n3925), .CK(clk), .SN(rst_n), .QN(Q7[16]) );
  DFFSX1 U1_Q3_i_reg_15_ ( .D(n3924), .CK(clk), .SN(rst_n), .QN(Q7[15]) );
  DFFSX1 U1_Q3_i_reg_14_ ( .D(n3923), .CK(clk), .SN(rst_n), .QN(Q7[14]) );
  DFFSX1 U1_Q3_i_reg_13_ ( .D(n3922), .CK(clk), .SN(rst_n), .QN(Q7[13]) );
  DFFSX1 U1_Q3_i_reg_12_ ( .D(n3921), .CK(clk), .SN(rst_n), .QN(Q7[12]) );
  DFFSX1 U1_Q3_i_reg_11_ ( .D(n3920), .CK(clk), .SN(rst_n), .QN(Q7[11]) );
  DFFSX1 U1_Q3_i_reg_10_ ( .D(n3919), .CK(clk), .SN(rst_n), .QN(Q7[10]) );
  DFFSX1 U1_Q3_i_reg_9_ ( .D(n3918), .CK(clk), .SN(rst_n), .QN(Q7[9]) );
  DFFSX1 U1_Q3_i_reg_8_ ( .D(n3917), .CK(clk), .SN(rst_n), .QN(Q7[8]) );
  DFFSX1 U1_Q3_i_reg_7_ ( .D(n3916), .CK(clk), .SN(rst_n), .QN(Q7[7]) );
  DFFSX1 U1_Q3_i_reg_6_ ( .D(n3915), .CK(clk), .SN(rst_n), .QN(Q7[6]) );
  DFFSX1 U1_Q3_i_reg_5_ ( .D(n3914), .CK(clk), .SN(rst_n), .QN(Q7[5]) );
  DFFSX1 U1_Q3_i_reg_4_ ( .D(n3913), .CK(clk), .SN(rst_n), .QN(Q7[4]) );
  DFFSX1 U1_Q3_i_reg_3_ ( .D(n3912), .CK(clk), .SN(rst_n), .QN(Q7[3]) );
  DFFSX1 U1_Q3_i_reg_2_ ( .D(n3911), .CK(clk), .SN(rst_n), .QN(Q7[2]) );
  DFFSX1 U1_Q3_i_reg_1_ ( .D(n3910), .CK(clk), .SN(rst_n), .QN(Q7[1]) );
  DFFSX1 U1_Q3_i_reg_0_ ( .D(n3909), .CK(clk), .SN(rst_n), .QN(Q7[0]) );
  DFFSX1 U1_Q3_r_reg_25_ ( .D(n3908), .CK(clk), .SN(rst_n), .QN(Q7[53]) );
  DFFSX1 U1_Q3_r_reg_24_ ( .D(n3907), .CK(clk), .SN(rst_n), .QN(Q7[52]) );
  DFFSX1 U1_Q3_r_reg_23_ ( .D(n3906), .CK(clk), .SN(rst_n), .QN(Q7[51]) );
  DFFSX1 U1_Q3_r_reg_22_ ( .D(n3905), .CK(clk), .SN(rst_n), .QN(Q7[50]) );
  DFFSX1 U1_Q3_r_reg_21_ ( .D(n3904), .CK(clk), .SN(rst_n), .QN(Q7[49]) );
  DFFSX1 U1_Q3_r_reg_20_ ( .D(n3903), .CK(clk), .SN(rst_n), .QN(Q7[48]) );
  DFFSX1 U1_Q3_r_reg_19_ ( .D(n3902), .CK(clk), .SN(rst_n), .QN(Q7[47]) );
  DFFSX1 U1_Q3_r_reg_18_ ( .D(n3901), .CK(clk), .SN(rst_n), .QN(Q7[46]) );
  DFFSX1 U1_Q3_r_reg_17_ ( .D(n3900), .CK(clk), .SN(rst_n), .QN(Q7[45]) );
  DFFSX1 U1_Q3_r_reg_16_ ( .D(n3899), .CK(clk), .SN(rst_n), .QN(Q7[44]) );
  DFFSX1 U1_Q3_r_reg_15_ ( .D(n3898), .CK(clk), .SN(rst_n), .QN(Q7[43]) );
  DFFSX1 U1_Q3_r_reg_14_ ( .D(n3897), .CK(clk), .SN(rst_n), .QN(Q7[42]) );
  DFFSX1 U1_Q3_r_reg_13_ ( .D(n3896), .CK(clk), .SN(rst_n), .QN(Q7[41]) );
  DFFSX1 U1_Q3_r_reg_12_ ( .D(n3895), .CK(clk), .SN(rst_n), .QN(Q7[40]) );
  DFFSX1 U1_Q3_r_reg_11_ ( .D(n3894), .CK(clk), .SN(rst_n), .QN(Q7[39]) );
  DFFSX1 U1_Q3_r_reg_10_ ( .D(n3893), .CK(clk), .SN(rst_n), .QN(Q7[38]) );
  DFFSX1 U1_Q3_r_reg_9_ ( .D(n3892), .CK(clk), .SN(rst_n), .QN(Q7[37]) );
  DFFSX1 U1_Q3_r_reg_8_ ( .D(n3891), .CK(clk), .SN(rst_n), .QN(Q7[36]) );
  DFFSX1 U1_Q3_r_reg_7_ ( .D(n3890), .CK(clk), .SN(rst_n), .QN(Q7[35]) );
  DFFSX1 U1_Q3_r_reg_6_ ( .D(n3889), .CK(clk), .SN(rst_n), .QN(Q7[34]) );
  DFFSX1 U1_Q3_r_reg_5_ ( .D(n3888), .CK(clk), .SN(rst_n), .QN(Q7[33]) );
  DFFSX1 U1_Q3_r_reg_4_ ( .D(n3887), .CK(clk), .SN(rst_n), .QN(Q7[32]) );
  DFFSX1 U1_Q3_r_reg_3_ ( .D(n3886), .CK(clk), .SN(rst_n), .QN(Q7[31]) );
  DFFSX1 U1_Q3_r_reg_2_ ( .D(n3885), .CK(clk), .SN(rst_n), .QN(Q7[30]) );
  DFFSX1 U1_Q3_r_reg_1_ ( .D(n3884), .CK(clk), .SN(rst_n), .QN(Q7[29]) );
  DFFSX1 U1_Q3_r_reg_0_ ( .D(n3883), .CK(clk), .SN(rst_n), .QN(Q7[28]) );
  DFFSX1 U1_Q2_i_reg_25_ ( .D(n3882), .CK(clk), .SN(rst_n), .QN(Q6[25]) );
  DFFSX1 U1_Q2_i_reg_24_ ( .D(n3881), .CK(clk), .SN(rst_n), .QN(Q6[24]) );
  DFFSX1 U1_Q2_i_reg_23_ ( .D(n3880), .CK(clk), .SN(rst_n), .QN(Q6[23]) );
  DFFSX1 U1_Q2_i_reg_22_ ( .D(n3879), .CK(clk), .SN(rst_n), .QN(Q6[22]) );
  DFFSX1 U1_Q2_i_reg_21_ ( .D(n3878), .CK(clk), .SN(rst_n), .QN(Q6[21]) );
  DFFSX1 U1_Q2_i_reg_20_ ( .D(n3877), .CK(clk), .SN(rst_n), .QN(Q6[20]) );
  DFFSX1 U1_Q2_i_reg_19_ ( .D(n3876), .CK(clk), .SN(rst_n), .QN(Q6[19]) );
  DFFSX1 U1_Q2_i_reg_18_ ( .D(n3875), .CK(clk), .SN(rst_n), .QN(Q6[18]) );
  DFFSX1 U1_Q2_i_reg_17_ ( .D(n3874), .CK(clk), .SN(rst_n), .QN(Q6[17]) );
  DFFSX1 U1_Q2_i_reg_16_ ( .D(n3873), .CK(clk), .SN(rst_n), .QN(Q6[16]) );
  DFFSX1 U1_Q2_i_reg_15_ ( .D(n3872), .CK(clk), .SN(rst_n), .QN(Q6[15]) );
  DFFSX1 U1_Q2_i_reg_14_ ( .D(n3871), .CK(clk), .SN(rst_n), .QN(Q6[14]) );
  DFFSX1 U1_Q2_i_reg_13_ ( .D(n3870), .CK(clk), .SN(rst_n), .QN(Q6[13]) );
  DFFSX1 U1_Q2_i_reg_12_ ( .D(n3869), .CK(clk), .SN(rst_n), .QN(Q6[12]) );
  DFFSX1 U1_Q2_i_reg_11_ ( .D(n3868), .CK(clk), .SN(rst_n), .QN(Q6[11]) );
  DFFSX1 U1_Q2_i_reg_10_ ( .D(n3867), .CK(clk), .SN(rst_n), .QN(Q6[10]) );
  DFFSX1 U1_Q2_i_reg_9_ ( .D(n3866), .CK(clk), .SN(rst_n), .QN(Q6[9]) );
  DFFSX1 U1_Q2_i_reg_8_ ( .D(n3865), .CK(clk), .SN(rst_n), .QN(Q6[8]) );
  DFFSX1 U1_Q2_i_reg_7_ ( .D(n3864), .CK(clk), .SN(rst_n), .QN(Q6[7]) );
  DFFSX1 U1_Q2_i_reg_6_ ( .D(n3863), .CK(clk), .SN(rst_n), .QN(Q6[6]) );
  DFFSX1 U1_Q2_i_reg_5_ ( .D(n3862), .CK(clk), .SN(rst_n), .QN(Q6[5]) );
  DFFSX1 U1_Q2_i_reg_4_ ( .D(n3861), .CK(clk), .SN(rst_n), .QN(Q6[4]) );
  DFFSX1 U1_Q2_i_reg_3_ ( .D(n3860), .CK(clk), .SN(rst_n), .QN(Q6[3]) );
  DFFSX1 U1_Q2_i_reg_2_ ( .D(n3859), .CK(clk), .SN(rst_n), .QN(Q6[2]) );
  DFFSX1 U1_Q2_i_reg_1_ ( .D(n3858), .CK(clk), .SN(rst_n), .QN(Q6[1]) );
  DFFSX1 U1_Q2_i_reg_0_ ( .D(n3857), .CK(clk), .SN(rst_n), .QN(Q6[0]) );
  DFFSX1 U1_Q2_r_reg_25_ ( .D(n3856), .CK(clk), .SN(rst_n), .QN(Q6[53]) );
  DFFSX1 U1_Q2_r_reg_24_ ( .D(n3855), .CK(clk), .SN(rst_n), .QN(Q6[52]) );
  DFFSX1 U1_Q2_r_reg_23_ ( .D(n3854), .CK(clk), .SN(rst_n), .QN(Q6[51]) );
  DFFSX1 U1_Q2_r_reg_22_ ( .D(n3853), .CK(clk), .SN(rst_n), .QN(Q6[50]) );
  DFFSX1 U1_Q2_r_reg_21_ ( .D(n3852), .CK(clk), .SN(rst_n), .QN(Q6[49]) );
  DFFSX1 U1_Q2_r_reg_20_ ( .D(n3851), .CK(clk), .SN(rst_n), .QN(Q6[48]) );
  DFFSX1 U1_Q2_r_reg_19_ ( .D(n3850), .CK(clk), .SN(rst_n), .QN(Q6[47]) );
  DFFSX1 U1_Q2_r_reg_18_ ( .D(n3849), .CK(clk), .SN(rst_n), .QN(Q6[46]) );
  DFFSX1 U1_Q2_r_reg_17_ ( .D(n3848), .CK(clk), .SN(rst_n), .QN(Q6[45]) );
  DFFSX1 U1_Q2_r_reg_16_ ( .D(n3847), .CK(clk), .SN(rst_n), .QN(Q6[44]) );
  DFFSX1 U1_Q2_r_reg_15_ ( .D(n3846), .CK(clk), .SN(rst_n), .QN(Q6[43]) );
  DFFSX1 U1_Q2_r_reg_14_ ( .D(n3845), .CK(clk), .SN(rst_n), .QN(Q6[42]) );
  DFFSX1 U1_Q2_r_reg_13_ ( .D(n3844), .CK(clk), .SN(rst_n), .QN(Q6[41]) );
  DFFSX1 R9_A_reg_9_ ( .D(n3843), .CK(clk), .SN(rst_n), .Q(n29036), .QN(
        BOPA[9]) );
  DFFSX2 R9_C_reg_9_ ( .D(n3841), .CK(clk), .SN(rst_n), .Q(n8117), .QN(BOPC[9]) );
  DFFSX1 R9_A_reg_8_ ( .D(n3839), .CK(clk), .SN(rst_n), .Q(n29035), .QN(
        BOPA[8]) );
  DFFSX2 R9_C_reg_7_ ( .D(n3833), .CK(clk), .SN(rst_n), .QN(BOPC[7]) );
  DFFSX2 R9_B_reg_7_ ( .D(n3832), .CK(clk), .SN(rst_n), .QN(BOPB[7]) );
  DFFSX2 R9_C_reg_6_ ( .D(n3829), .CK(clk), .SN(rst_n), .Q(n8124), .QN(BOPC[6]) );
  DFFSX2 R9_B_reg_6_ ( .D(n3828), .CK(clk), .SN(rst_n), .Q(n8123), .QN(BOPB[6]) );
  DFFSX1 R9_A_reg_51_ ( .D(n3823), .CK(clk), .SN(rst_n), .Q(n28749), .QN(
        BOPA[51]) );
  DFFSX1 R9_D_reg_51_ ( .D(n3822), .CK(clk), .SN(rst_n), .Q(n8131), .QN(
        BOPD[51]) );
  DFFSX1 R9_C_reg_51_ ( .D(n3821), .CK(clk), .SN(rst_n), .Q(n8130), .QN(
        BOPC[51]) );
  DFFSX1 R9_B_reg_51_ ( .D(n3820), .CK(clk), .SN(rst_n), .Q(n8129), .QN(
        BOPB[51]) );
  DFFSX1 R9_A_reg_50_ ( .D(n3819), .CK(clk), .SN(rst_n), .Q(n28687), .QN(
        BOPA[50]) );
  DFFSX1 R9_D_reg_50_ ( .D(n3818), .CK(clk), .SN(rst_n), .QN(BOPD[50]) );
  DFFSX1 R9_C_reg_50_ ( .D(n3817), .CK(clk), .SN(rst_n), .QN(BOPC[50]) );
  DFFSX1 R9_B_reg_50_ ( .D(n3816), .CK(clk), .SN(rst_n), .QN(BOPB[50]) );
  DFFSX2 R9_D_reg_4_ ( .D(n3814), .CK(clk), .SN(rst_n), .Q(n8134), .QN(BOPD[4]) );
  DFFSX1 R9_A_reg_49_ ( .D(n3811), .CK(clk), .SN(rst_n), .Q(n28684), .QN(
        BOPA[49]) );
  DFFSX1 R9_D_reg_49_ ( .D(n3810), .CK(clk), .SN(rst_n), .QN(BOPD[49]) );
  DFFSX1 R9_C_reg_49_ ( .D(n3809), .CK(clk), .SN(rst_n), .QN(BOPC[49]) );
  DFFSX1 R9_B_reg_49_ ( .D(n3808), .CK(clk), .SN(rst_n), .QN(BOPB[49]) );
  DFFSX1 R9_A_reg_48_ ( .D(n3807), .CK(clk), .SN(rst_n), .Q(n28710), .QN(
        BOPA[48]) );
  DFFSX1 R9_D_reg_48_ ( .D(n3806), .CK(clk), .SN(rst_n), .QN(BOPD[48]) );
  DFFSX1 R9_C_reg_48_ ( .D(n3805), .CK(clk), .SN(rst_n), .QN(BOPC[48]) );
  DFFSX1 R9_B_reg_48_ ( .D(n3804), .CK(clk), .SN(rst_n), .QN(BOPB[48]) );
  DFFSX1 R9_D_reg_47_ ( .D(n3802), .CK(clk), .SN(rst_n), .QN(BOPD[47]) );
  DFFSX1 R9_C_reg_47_ ( .D(n3801), .CK(clk), .SN(rst_n), .QN(BOPC[47]) );
  DFFSX1 R9_B_reg_47_ ( .D(n3800), .CK(clk), .SN(rst_n), .QN(BOPB[47]) );
  DFFSX1 R9_D_reg_46_ ( .D(n3798), .CK(clk), .SN(rst_n), .QN(BOPD[46]) );
  DFFSX1 R9_C_reg_46_ ( .D(n3797), .CK(clk), .SN(rst_n), .QN(BOPC[46]) );
  DFFSX1 R9_B_reg_46_ ( .D(n3796), .CK(clk), .SN(rst_n), .QN(BOPB[46]) );
  DFFSX1 R9_D_reg_44_ ( .D(n3790), .CK(clk), .SN(rst_n), .QN(BOPD[44]) );
  DFFSX1 R9_B_reg_44_ ( .D(n3788), .CK(clk), .SN(rst_n), .QN(BOPB[44]) );
  DFFSX2 R9_B_reg_43_ ( .D(n3784), .CK(clk), .SN(rst_n), .QN(BOPB[43]) );
  DFFSX2 R9_C_reg_42_ ( .D(n3781), .CK(clk), .SN(rst_n), .QN(BOPC[42]) );
  DFFSX1 R9_B_reg_41_ ( .D(n3776), .CK(clk), .SN(rst_n), .QN(BOPB[41]) );
  DFFSX4 R9_D_reg_3_ ( .D(n3770), .CK(clk), .SN(rst_n), .Q(n8137), .QN(BOPD[3]) );
  DFFSX4 R9_B_reg_3_ ( .D(n3768), .CK(clk), .SN(rst_n), .Q(n8135), .QN(BOPB[3]) );
  DFFSX2 R9_D_reg_39_ ( .D(n3766), .CK(clk), .SN(rst_n), .QN(BOPD[39]) );
  DFFSX2 R9_B_reg_39_ ( .D(n3764), .CK(clk), .SN(rst_n), .QN(BOPB[39]) );
  DFFSX4 R9_A_reg_38_ ( .D(n3763), .CK(clk), .SN(rst_n), .Q(n28713), .QN(
        BOPA[38]) );
  DFFSX2 R9_B_reg_38_ ( .D(n3760), .CK(clk), .SN(rst_n), .QN(BOPB[38]) );
  DFFSX2 R9_B_reg_37_ ( .D(n3756), .CK(clk), .SN(rst_n), .QN(BOPB[37]) );
  DFFSX2 R9_B_reg_35_ ( .D(n3748), .CK(clk), .SN(rst_n), .QN(BOPB[35]) );
  DFFSX4 R9_A_reg_34_ ( .D(n3747), .CK(clk), .SN(rst_n), .Q(n6910), .QN(
        BOPA[34]) );
  DFFSX2 R9_D_reg_34_ ( .D(n3746), .CK(clk), .SN(rst_n), .QN(BOPD[34]) );
  DFFSX2 R9_B_reg_34_ ( .D(n3744), .CK(clk), .SN(rst_n), .QN(BOPB[34]) );
  DFFSX4 R9_A_reg_33_ ( .D(n3743), .CK(clk), .SN(rst_n), .Q(n29100), .QN(
        BOPA[33]) );
  DFFSX1 R9_D_reg_33_ ( .D(n3742), .CK(clk), .SN(rst_n), .QN(BOPD[33]) );
  DFFSX4 R9_A_reg_32_ ( .D(n3739), .CK(clk), .SN(rst_n), .Q(n28750), .QN(
        BOPA[32]) );
  DFFSX4 R9_A_reg_31_ ( .D(n3735), .CK(clk), .SN(rst_n), .Q(n29105), .QN(
        BOPA[31]) );
  DFFSX4 R9_D_reg_2_ ( .D(n3726), .CK(clk), .SN(rst_n), .Q(n8139), .QN(BOPD[2]) );
  DFFSX4 R9_C_reg_2_ ( .D(n3725), .CK(clk), .SN(rst_n), .Q(n8138), .QN(BOPC[2]) );
  DFFSX4 R9_B_reg_2_ ( .D(n3724), .CK(clk), .SN(rst_n), .Q(n7051), .QN(BOPB[2]) );
  DFFSX4 R9_A_reg_29_ ( .D(n3723), .CK(clk), .SN(rst_n), .Q(n29103), .QN(
        BOPA[29]) );
  DFFSX4 R9_A_reg_28_ ( .D(n3719), .CK(clk), .SN(rst_n), .Q(n29102), .QN(
        BOPA[28]) );
  DFFSX2 R9_D_reg_28_ ( .D(n3718), .CK(clk), .SN(rst_n), .QN(BOPD[28]) );
  DFFSX2 R9_B_reg_28_ ( .D(n3716), .CK(clk), .SN(rst_n), .QN(BOPB[28]) );
  DFFSX4 R9_A_reg_27_ ( .D(n3715), .CK(clk), .SN(rst_n), .Q(n28682), .QN(
        BOPA[27]) );
  DFFSX2 R9_D_reg_27_ ( .D(n3714), .CK(clk), .SN(rst_n), .QN(BOPD[27]) );
  DFFSX4 R9_A_reg_26_ ( .D(n3711), .CK(clk), .SN(rst_n), .Q(n28751), .QN(
        BOPA[26]) );
  DFFSX2 R9_D_reg_26_ ( .D(n3710), .CK(clk), .SN(rst_n), .QN(BOPD[26]) );
  DFFSX2 R9_C_reg_26_ ( .D(n3709), .CK(clk), .SN(rst_n), .QN(BOPC[26]) );
  DFFSX2 R9_B_reg_26_ ( .D(n3708), .CK(clk), .SN(rst_n), .QN(BOPB[26]) );
  DFFSX1 R9_A_reg_25_ ( .D(n3707), .CK(clk), .SN(rst_n), .Q(n29031), .QN(
        BOPA[25]) );
  DFFSX1 R9_D_reg_25_ ( .D(n3706), .CK(clk), .SN(rst_n), .QN(BOPD[25]) );
  DFFSX1 R9_C_reg_25_ ( .D(n3705), .CK(clk), .SN(rst_n), .QN(BOPC[25]) );
  DFFSX1 R9_B_reg_25_ ( .D(n3704), .CK(clk), .SN(rst_n), .QN(BOPB[25]) );
  DFFSX1 R9_A_reg_24_ ( .D(n3703), .CK(clk), .SN(rst_n), .Q(n29030), .QN(
        BOPA[24]) );
  DFFSX1 R9_D_reg_24_ ( .D(n3702), .CK(clk), .SN(rst_n), .Q(n8152), .QN(
        BOPD[24]) );
  DFFSX1 R9_C_reg_24_ ( .D(n3701), .CK(clk), .SN(rst_n), .Q(n8151), .QN(
        BOPC[24]) );
  DFFSX1 R9_B_reg_24_ ( .D(n3700), .CK(clk), .SN(rst_n), .Q(n8150), .QN(
        BOPB[24]) );
  DFFSX1 R9_A_reg_23_ ( .D(n3699), .CK(clk), .SN(rst_n), .Q(n29029), .QN(
        BOPA[23]) );
  DFFSX1 R9_D_reg_23_ ( .D(n3698), .CK(clk), .SN(rst_n), .Q(n8155), .QN(
        BOPD[23]) );
  DFFSX1 R9_C_reg_23_ ( .D(n3697), .CK(clk), .SN(rst_n), .Q(n8154), .QN(
        BOPC[23]) );
  DFFSX1 R9_B_reg_23_ ( .D(n3696), .CK(clk), .SN(rst_n), .Q(n8153), .QN(
        BOPB[23]) );
  DFFSX1 R9_A_reg_22_ ( .D(n3695), .CK(clk), .SN(rst_n), .Q(n29028), .QN(
        BOPA[22]) );
  DFFSX1 R9_D_reg_22_ ( .D(n3694), .CK(clk), .SN(rst_n), .Q(n8159), .QN(
        BOPD[22]) );
  DFFSX1 R9_C_reg_22_ ( .D(n3693), .CK(clk), .SN(rst_n), .Q(n8158), .QN(
        BOPC[22]) );
  DFFSX1 R9_B_reg_22_ ( .D(n3692), .CK(clk), .SN(rst_n), .Q(n8157), .QN(
        BOPB[22]) );
  DFFSX1 R9_A_reg_21_ ( .D(n3691), .CK(clk), .SN(rst_n), .Q(n29027), .QN(
        BOPA[21]) );
  DFFSX1 R9_A_reg_20_ ( .D(n3687), .CK(clk), .SN(rst_n), .Q(n29026), .QN(
        BOPA[20]) );
  DFFSX1 R9_D_reg_20_ ( .D(n3686), .CK(clk), .SN(rst_n), .Q(n8165), .QN(
        BOPD[20]) );
  DFFSX1 R9_C_reg_20_ ( .D(n3685), .CK(clk), .SN(rst_n), .Q(n8164), .QN(
        BOPC[20]) );
  DFFSX1 R9_B_reg_20_ ( .D(n3684), .CK(clk), .SN(rst_n), .Q(n8163), .QN(
        BOPB[20]) );
  DFFSX4 R9_D_reg_1_ ( .D(n3682), .CK(clk), .SN(rst_n), .Q(n8168), .QN(BOPD[1]) );
  DFFSX2 R9_C_reg_1_ ( .D(n3681), .CK(clk), .SN(rst_n), .Q(n8167), .QN(BOPC[1]) );
  DFFSX1 R9_A_reg_19_ ( .D(n3679), .CK(clk), .SN(rst_n), .Q(n29025), .QN(
        BOPA[19]) );
  DFFSX1 R9_A_reg_18_ ( .D(n3675), .CK(clk), .SN(rst_n), .Q(n29024), .QN(
        BOPA[18]) );
  DFFSX1 R9_A_reg_17_ ( .D(n3671), .CK(clk), .SN(rst_n), .Q(n29023), .QN(
        BOPA[17]) );
  DFFSX1 R9_A_reg_16_ ( .D(n3667), .CK(clk), .SN(rst_n), .Q(n29022), .QN(
        BOPA[16]) );
  DFFSX1 R9_A_reg_15_ ( .D(n3663), .CK(clk), .SN(rst_n), .Q(n29015), .QN(
        BOPA[15]) );
  DFFSX2 R9_B_reg_15_ ( .D(n3660), .CK(clk), .SN(rst_n), .Q(n8179), .QN(
        BOPB[15]) );
  DFFSX1 R9_A_reg_14_ ( .D(n3659), .CK(clk), .SN(rst_n), .Q(n29021), .QN(
        BOPA[14]) );
  DFFSX2 R9_B_reg_14_ ( .D(n3656), .CK(clk), .SN(rst_n), .Q(n6944), .QN(
        BOPB[14]) );
  DFFSX1 R9_A_reg_13_ ( .D(n3655), .CK(clk), .SN(rst_n), .Q(n29014), .QN(
        BOPA[13]) );
  DFFSX1 R9_A_reg_12_ ( .D(n3651), .CK(clk), .SN(rst_n), .Q(n29020), .QN(
        BOPA[12]) );
  DFFSX2 R9_C_reg_12_ ( .D(n3649), .CK(clk), .SN(rst_n), .Q(n8185), .QN(
        BOPC[12]) );
  DFFSX1 R9_A_reg_11_ ( .D(n3647), .CK(clk), .SN(rst_n), .Q(n29019), .QN(
        BOPA[11]) );
  DFFSX1 R9_A_reg_10_ ( .D(n3643), .CK(clk), .SN(rst_n), .Q(n29018), .QN(
        BOPA[10]) );
  DFFSX4 R9_D_reg_0_ ( .D(n3638), .CK(clk), .SN(rst_n), .Q(n7991), .QN(BOPD[0]) );
  DFFSX1 U0_Q2_r_reg_13_ ( .D(n3635), .CK(clk), .SN(rst_n), .QN(Q2[41]) );
  DFFSX1 U0_Q2_r_reg_14_ ( .D(n3634), .CK(clk), .SN(rst_n), .QN(Q2[42]) );
  DFFSX1 U0_Q2_r_reg_15_ ( .D(n3633), .CK(clk), .SN(rst_n), .QN(Q2[43]) );
  DFFSX1 U0_Q2_r_reg_16_ ( .D(n3632), .CK(clk), .SN(rst_n), .QN(Q2[44]) );
  DFFSX1 U0_Q2_r_reg_17_ ( .D(n3631), .CK(clk), .SN(rst_n), .QN(Q2[45]) );
  DFFSX1 U0_Q2_r_reg_18_ ( .D(n3630), .CK(clk), .SN(rst_n), .QN(Q2[46]) );
  DFFSX1 U0_Q2_r_reg_19_ ( .D(n3629), .CK(clk), .SN(rst_n), .QN(Q2[47]) );
  DFFSX1 U0_Q2_r_reg_20_ ( .D(n3628), .CK(clk), .SN(rst_n), .QN(Q2[48]) );
  DFFSX1 U0_Q2_r_reg_21_ ( .D(n3627), .CK(clk), .SN(rst_n), .QN(Q2[49]) );
  DFFSX1 U0_Q2_r_reg_22_ ( .D(n3626), .CK(clk), .SN(rst_n), .QN(Q2[50]) );
  DFFSX1 U0_Q2_r_reg_23_ ( .D(n3625), .CK(clk), .SN(rst_n), .QN(Q2[51]) );
  DFFSX1 U0_Q2_r_reg_24_ ( .D(n3624), .CK(clk), .SN(rst_n), .QN(Q2[52]) );
  DFFSX1 U0_Q2_r_reg_25_ ( .D(n3623), .CK(clk), .SN(rst_n), .QN(Q2[53]) );
  DFFSX1 U0_Q2_i_reg_0_ ( .D(n3622), .CK(clk), .SN(rst_n), .QN(Q2[0]) );
  DFFSX1 U0_Q2_i_reg_1_ ( .D(n3621), .CK(clk), .SN(rst_n), .QN(Q2[1]) );
  DFFSX1 U0_Q2_i_reg_2_ ( .D(n3620), .CK(clk), .SN(rst_n), .QN(Q2[2]) );
  DFFSX1 U0_Q2_i_reg_3_ ( .D(n3619), .CK(clk), .SN(rst_n), .QN(Q2[3]) );
  DFFSX1 U0_Q2_i_reg_4_ ( .D(n3618), .CK(clk), .SN(rst_n), .QN(Q2[4]) );
  DFFSX1 U0_Q2_i_reg_5_ ( .D(n3617), .CK(clk), .SN(rst_n), .QN(Q2[5]) );
  DFFSX1 U0_Q2_i_reg_6_ ( .D(n3616), .CK(clk), .SN(rst_n), .QN(Q2[6]) );
  DFFSX1 U0_Q2_i_reg_7_ ( .D(n3615), .CK(clk), .SN(rst_n), .QN(Q2[7]) );
  DFFSX1 U0_Q2_i_reg_8_ ( .D(n3614), .CK(clk), .SN(rst_n), .QN(Q2[8]) );
  DFFSX1 U0_Q2_i_reg_9_ ( .D(n3613), .CK(clk), .SN(rst_n), .QN(Q2[9]) );
  DFFSX1 U0_Q2_i_reg_10_ ( .D(n3612), .CK(clk), .SN(rst_n), .QN(Q2[10]) );
  DFFSX1 U0_Q2_i_reg_11_ ( .D(n3611), .CK(clk), .SN(rst_n), .QN(Q2[11]) );
  DFFSX1 U0_Q2_i_reg_12_ ( .D(n3610), .CK(clk), .SN(rst_n), .QN(Q2[12]) );
  DFFSX1 U0_Q2_i_reg_13_ ( .D(n3609), .CK(clk), .SN(rst_n), .QN(Q2[13]) );
  DFFSX1 U0_Q2_i_reg_14_ ( .D(n3608), .CK(clk), .SN(rst_n), .QN(Q2[14]) );
  DFFSX1 U0_Q2_i_reg_15_ ( .D(n3607), .CK(clk), .SN(rst_n), .QN(Q2[15]) );
  DFFSX1 U0_Q2_i_reg_16_ ( .D(n3606), .CK(clk), .SN(rst_n), .QN(Q2[16]) );
  DFFSX1 U0_Q2_i_reg_17_ ( .D(n3605), .CK(clk), .SN(rst_n), .QN(Q2[17]) );
  DFFSX1 U0_Q2_i_reg_18_ ( .D(n3604), .CK(clk), .SN(rst_n), .QN(Q2[18]) );
  DFFSX1 U0_Q2_i_reg_19_ ( .D(n3603), .CK(clk), .SN(rst_n), .QN(Q2[19]) );
  DFFSX1 U0_Q2_i_reg_20_ ( .D(n3602), .CK(clk), .SN(rst_n), .QN(Q2[20]) );
  DFFSX1 U0_Q2_i_reg_21_ ( .D(n3601), .CK(clk), .SN(rst_n), .QN(Q2[21]) );
  DFFSX1 U0_Q2_i_reg_22_ ( .D(n3600), .CK(clk), .SN(rst_n), .QN(Q2[22]) );
  DFFSX1 U0_Q2_i_reg_23_ ( .D(n3599), .CK(clk), .SN(rst_n), .QN(Q2[23]) );
  DFFSX1 U0_Q2_i_reg_24_ ( .D(n3598), .CK(clk), .SN(rst_n), .QN(Q2[24]) );
  DFFSX1 U0_Q2_i_reg_25_ ( .D(n3597), .CK(clk), .SN(rst_n), .QN(Q2[25]) );
  DFFSX1 U0_Q3_r_reg_0_ ( .D(n3596), .CK(clk), .SN(rst_n), .QN(Q3[28]) );
  DFFSX1 U0_Q3_r_reg_1_ ( .D(n3595), .CK(clk), .SN(rst_n), .QN(Q3[29]) );
  DFFSX1 U0_Q3_r_reg_2_ ( .D(n3594), .CK(clk), .SN(rst_n), .QN(Q3[30]) );
  DFFSX1 U0_Q3_r_reg_3_ ( .D(n3593), .CK(clk), .SN(rst_n), .QN(Q3[31]) );
  DFFSX1 U0_Q3_r_reg_4_ ( .D(n3592), .CK(clk), .SN(rst_n), .QN(Q3[32]) );
  DFFSX1 U0_Q3_r_reg_5_ ( .D(n3591), .CK(clk), .SN(rst_n), .QN(Q3[33]) );
  DFFSX1 U0_Q3_r_reg_6_ ( .D(n3590), .CK(clk), .SN(rst_n), .QN(Q3[34]) );
  DFFSX1 U0_Q3_r_reg_7_ ( .D(n3589), .CK(clk), .SN(rst_n), .QN(Q3[35]) );
  DFFSX1 U0_Q3_r_reg_8_ ( .D(n3588), .CK(clk), .SN(rst_n), .QN(Q3[36]) );
  DFFSX1 U0_Q3_r_reg_9_ ( .D(n3587), .CK(clk), .SN(rst_n), .QN(Q3[37]) );
  DFFSX1 U0_Q3_r_reg_10_ ( .D(n3586), .CK(clk), .SN(rst_n), .QN(Q3[38]) );
  DFFSX1 U0_Q3_r_reg_11_ ( .D(n3585), .CK(clk), .SN(rst_n), .QN(Q3[39]) );
  DFFSX1 U0_Q3_r_reg_12_ ( .D(n3584), .CK(clk), .SN(rst_n), .QN(Q3[40]) );
  DFFSX1 U0_Q3_r_reg_13_ ( .D(n3583), .CK(clk), .SN(rst_n), .QN(Q3[41]) );
  DFFSX1 U0_Q3_r_reg_14_ ( .D(n3582), .CK(clk), .SN(rst_n), .QN(Q3[42]) );
  DFFSX1 U0_Q3_r_reg_15_ ( .D(n3581), .CK(clk), .SN(rst_n), .QN(Q3[43]) );
  DFFSX1 U0_Q3_r_reg_16_ ( .D(n3580), .CK(clk), .SN(rst_n), .QN(Q3[44]) );
  DFFSX1 U0_Q3_r_reg_17_ ( .D(n3579), .CK(clk), .SN(rst_n), .QN(Q3[45]) );
  DFFSX1 U0_Q3_r_reg_18_ ( .D(n3578), .CK(clk), .SN(rst_n), .QN(Q3[46]) );
  DFFSX1 U0_Q3_r_reg_19_ ( .D(n3577), .CK(clk), .SN(rst_n), .QN(Q3[47]) );
  DFFSX1 U0_Q3_r_reg_20_ ( .D(n3576), .CK(clk), .SN(rst_n), .QN(Q3[48]) );
  DFFSX1 U0_Q3_r_reg_21_ ( .D(n3575), .CK(clk), .SN(rst_n), .QN(Q3[49]) );
  DFFSX1 U0_Q3_r_reg_22_ ( .D(n3574), .CK(clk), .SN(rst_n), .QN(Q3[50]) );
  DFFSX1 U0_Q3_r_reg_23_ ( .D(n3573), .CK(clk), .SN(rst_n), .QN(Q3[51]) );
  DFFSX1 U0_Q3_r_reg_24_ ( .D(n3572), .CK(clk), .SN(rst_n), .QN(Q3[52]) );
  DFFSX1 U0_Q3_r_reg_25_ ( .D(n3571), .CK(clk), .SN(rst_n), .QN(Q3[53]) );
  DFFSX1 U0_Q3_i_reg_0_ ( .D(n3570), .CK(clk), .SN(rst_n), .QN(Q3[0]) );
  DFFSX1 U0_Q3_i_reg_1_ ( .D(n3569), .CK(clk), .SN(rst_n), .QN(Q3[1]) );
  DFFSX1 U0_Q3_i_reg_2_ ( .D(n3568), .CK(clk), .SN(rst_n), .QN(Q3[2]) );
  DFFSX1 U0_Q3_i_reg_3_ ( .D(n3567), .CK(clk), .SN(rst_n), .QN(Q3[3]) );
  DFFSX1 U0_Q3_i_reg_4_ ( .D(n3566), .CK(clk), .SN(rst_n), .QN(Q3[4]) );
  DFFSX1 U0_Q3_i_reg_5_ ( .D(n3565), .CK(clk), .SN(rst_n), .QN(Q3[5]) );
  DFFSX1 U0_Q3_i_reg_6_ ( .D(n3564), .CK(clk), .SN(rst_n), .QN(Q3[6]) );
  DFFSX1 U0_Q3_i_reg_7_ ( .D(n3563), .CK(clk), .SN(rst_n), .QN(Q3[7]) );
  DFFSX1 U0_Q3_i_reg_8_ ( .D(n3562), .CK(clk), .SN(rst_n), .QN(Q3[8]) );
  DFFSX1 U0_Q3_i_reg_9_ ( .D(n3561), .CK(clk), .SN(rst_n), .QN(Q3[9]) );
  DFFSX1 U0_Q3_i_reg_10_ ( .D(n3560), .CK(clk), .SN(rst_n), .QN(Q3[10]) );
  DFFSX1 U0_Q3_i_reg_11_ ( .D(n3559), .CK(clk), .SN(rst_n), .QN(Q3[11]) );
  DFFSX1 U0_Q3_i_reg_12_ ( .D(n3558), .CK(clk), .SN(rst_n), .QN(Q3[12]) );
  DFFSX1 U0_Q3_i_reg_13_ ( .D(n3557), .CK(clk), .SN(rst_n), .QN(Q3[13]) );
  DFFSX1 U0_Q3_i_reg_14_ ( .D(n3556), .CK(clk), .SN(rst_n), .QN(Q3[14]) );
  DFFSX1 U0_Q3_i_reg_15_ ( .D(n3555), .CK(clk), .SN(rst_n), .QN(Q3[15]) );
  DFFSX1 U0_Q3_i_reg_16_ ( .D(n3554), .CK(clk), .SN(rst_n), .QN(Q3[16]) );
  DFFSX1 U0_Q3_i_reg_17_ ( .D(n3553), .CK(clk), .SN(rst_n), .QN(Q3[17]) );
  DFFSX1 U0_Q3_i_reg_18_ ( .D(n3552), .CK(clk), .SN(rst_n), .QN(Q3[18]) );
  DFFSX1 U0_Q3_i_reg_19_ ( .D(n3551), .CK(clk), .SN(rst_n), .QN(Q3[19]) );
  DFFSX1 U0_Q3_i_reg_20_ ( .D(n3550), .CK(clk), .SN(rst_n), .QN(Q3[20]) );
  DFFSX1 U0_Q3_i_reg_21_ ( .D(n3549), .CK(clk), .SN(rst_n), .QN(Q3[21]) );
  DFFSX1 U0_Q3_i_reg_22_ ( .D(n3548), .CK(clk), .SN(rst_n), .QN(Q3[22]) );
  DFFSX1 U0_Q3_i_reg_23_ ( .D(n3547), .CK(clk), .SN(rst_n), .QN(Q3[23]) );
  DFFSX1 U0_Q3_i_reg_24_ ( .D(n3546), .CK(clk), .SN(rst_n), .QN(Q3[24]) );
  DFFSX1 U0_Q3_i_reg_25_ ( .D(n3545), .CK(clk), .SN(rst_n), .QN(Q3[25]) );
  DFFSX1 U0_Q0_r_reg_0_ ( .D(n3544), .CK(clk), .SN(rst_n), .QN(Q0[28]) );
  DFFSX1 U0_Q0_i_reg_0_ ( .D(n3543), .CK(clk), .SN(rst_n), .QN(Q0[0]) );
  DFFSX1 U0_Q0_i_reg_1_ ( .D(n3542), .CK(clk), .SN(rst_n), .QN(Q0[1]) );
  DFFSX1 U0_Q0_i_reg_2_ ( .D(n3541), .CK(clk), .SN(rst_n), .QN(Q0[2]) );
  DFFSX1 U0_Q0_i_reg_3_ ( .D(n3540), .CK(clk), .SN(rst_n), .QN(Q0[3]) );
  DFFSX1 U0_Q0_i_reg_4_ ( .D(n3539), .CK(clk), .SN(rst_n), .QN(Q0[4]) );
  DFFSX1 U0_Q0_i_reg_5_ ( .D(n3538), .CK(clk), .SN(rst_n), .QN(Q0[5]) );
  DFFSX1 U0_Q0_i_reg_6_ ( .D(n3537), .CK(clk), .SN(rst_n), .QN(Q0[6]) );
  DFFSX1 U0_Q0_i_reg_7_ ( .D(n3536), .CK(clk), .SN(rst_n), .QN(Q0[7]) );
  DFFSX1 U0_Q0_i_reg_8_ ( .D(n3535), .CK(clk), .SN(rst_n), .QN(Q0[8]) );
  DFFSX1 U0_Q0_i_reg_9_ ( .D(n3534), .CK(clk), .SN(rst_n), .QN(Q0[9]) );
  DFFSX1 U0_Q0_i_reg_10_ ( .D(n3533), .CK(clk), .SN(rst_n), .QN(Q0[10]) );
  DFFSX1 U0_Q0_i_reg_11_ ( .D(n3532), .CK(clk), .SN(rst_n), .QN(Q0[11]) );
  DFFSX1 U0_Q0_i_reg_12_ ( .D(n3531), .CK(clk), .SN(rst_n), .QN(Q0[12]) );
  DFFSX1 U0_Q0_i_reg_13_ ( .D(n3530), .CK(clk), .SN(rst_n), .QN(Q0[13]) );
  DFFSX1 U0_Q0_i_reg_14_ ( .D(n3529), .CK(clk), .SN(rst_n), .QN(Q0[14]) );
  DFFSX1 U0_Q0_i_reg_15_ ( .D(n3528), .CK(clk), .SN(rst_n), .QN(Q0[15]) );
  DFFSX1 U0_Q0_i_reg_16_ ( .D(n3527), .CK(clk), .SN(rst_n), .QN(Q0[16]) );
  DFFSX1 U0_Q0_i_reg_17_ ( .D(n3526), .CK(clk), .SN(rst_n), .QN(Q0[17]) );
  DFFSX1 U0_Q0_i_reg_18_ ( .D(n3525), .CK(clk), .SN(rst_n), .QN(Q0[18]) );
  DFFSX1 U0_Q0_i_reg_19_ ( .D(n3524), .CK(clk), .SN(rst_n), .QN(Q0[19]) );
  DFFSX1 U0_Q0_i_reg_20_ ( .D(n3523), .CK(clk), .SN(rst_n), .QN(Q0[20]) );
  DFFSX1 U0_Q0_i_reg_21_ ( .D(n3522), .CK(clk), .SN(rst_n), .QN(Q0[21]) );
  DFFSX1 U0_Q0_i_reg_22_ ( .D(n3521), .CK(clk), .SN(rst_n), .QN(Q0[22]) );
  DFFSX1 U0_Q0_i_reg_23_ ( .D(n3520), .CK(clk), .SN(rst_n), .QN(Q0[23]) );
  DFFSX1 U0_Q0_i_reg_24_ ( .D(n3519), .CK(clk), .SN(rst_n), .QN(Q0[24]) );
  DFFSX1 U0_Q0_i_reg_25_ ( .D(n3518), .CK(clk), .SN(rst_n), .QN(Q0[25]) );
  DFFSX1 U0_Q1_r_reg_0_ ( .D(n3517), .CK(clk), .SN(rst_n), .QN(Q1[28]) );
  DFFSX1 U0_Q1_r_reg_1_ ( .D(n3516), .CK(clk), .SN(rst_n), .QN(Q1[29]) );
  DFFSX1 U0_Q1_r_reg_2_ ( .D(n3515), .CK(clk), .SN(rst_n), .QN(Q1[30]) );
  DFFSX1 U0_Q1_r_reg_3_ ( .D(n3514), .CK(clk), .SN(rst_n), .QN(Q1[31]) );
  DFFSX1 U0_Q1_r_reg_4_ ( .D(n3513), .CK(clk), .SN(rst_n), .QN(Q1[32]) );
  DFFSX1 U0_Q1_r_reg_5_ ( .D(n3512), .CK(clk), .SN(rst_n), .QN(Q1[33]) );
  DFFSX1 U0_Q1_r_reg_6_ ( .D(n3511), .CK(clk), .SN(rst_n), .QN(Q1[34]) );
  DFFSX1 U0_Q1_r_reg_7_ ( .D(n3510), .CK(clk), .SN(rst_n), .QN(Q1[35]) );
  DFFSX1 U0_Q1_r_reg_8_ ( .D(n3509), .CK(clk), .SN(rst_n), .QN(Q1[36]) );
  DFFSX1 U0_Q1_r_reg_9_ ( .D(n3508), .CK(clk), .SN(rst_n), .QN(Q1[37]) );
  DFFSX1 U0_Q1_r_reg_10_ ( .D(n3507), .CK(clk), .SN(rst_n), .QN(Q1[38]) );
  DFFSX1 U0_Q1_r_reg_11_ ( .D(n3506), .CK(clk), .SN(rst_n), .QN(Q1[39]) );
  DFFSX1 U0_Q1_r_reg_12_ ( .D(n3505), .CK(clk), .SN(rst_n), .QN(Q1[40]) );
  DFFSX1 U0_Q1_r_reg_13_ ( .D(n3504), .CK(clk), .SN(rst_n), .QN(Q1[41]) );
  DFFSX1 U0_Q1_r_reg_14_ ( .D(n3503), .CK(clk), .SN(rst_n), .QN(Q1[42]) );
  DFFSX1 U0_Q1_r_reg_15_ ( .D(n3502), .CK(clk), .SN(rst_n), .QN(Q1[43]) );
  DFFSX1 U0_Q1_r_reg_16_ ( .D(n3501), .CK(clk), .SN(rst_n), .QN(Q1[44]) );
  DFFSX1 U0_Q1_r_reg_17_ ( .D(n3500), .CK(clk), .SN(rst_n), .QN(Q1[45]) );
  DFFSX1 U0_Q1_r_reg_18_ ( .D(n3499), .CK(clk), .SN(rst_n), .QN(Q1[46]) );
  DFFSX1 U0_Q1_r_reg_19_ ( .D(n3498), .CK(clk), .SN(rst_n), .QN(Q1[47]) );
  DFFSX1 U0_Q1_r_reg_20_ ( .D(n3497), .CK(clk), .SN(rst_n), .QN(Q1[48]) );
  DFFSX1 U0_Q1_r_reg_21_ ( .D(n3496), .CK(clk), .SN(rst_n), .QN(Q1[49]) );
  DFFSX1 U0_Q1_r_reg_22_ ( .D(n3495), .CK(clk), .SN(rst_n), .QN(Q1[50]) );
  DFFSX1 U0_Q1_r_reg_23_ ( .D(n3494), .CK(clk), .SN(rst_n), .QN(Q1[51]) );
  DFFSX1 U0_Q1_r_reg_24_ ( .D(n3493), .CK(clk), .SN(rst_n), .QN(Q1[52]) );
  DFFSX1 U0_Q1_r_reg_25_ ( .D(n3492), .CK(clk), .SN(rst_n), .QN(Q1[53]) );
  DFFSX1 U0_Q1_i_reg_0_ ( .D(n3491), .CK(clk), .SN(rst_n), .QN(Q1[0]) );
  DFFSX1 U0_Q1_i_reg_1_ ( .D(n3490), .CK(clk), .SN(rst_n), .QN(Q1[1]) );
  DFFSX1 U0_Q1_i_reg_2_ ( .D(n3489), .CK(clk), .SN(rst_n), .QN(Q1[2]) );
  DFFSX1 U0_Q1_i_reg_3_ ( .D(n3488), .CK(clk), .SN(rst_n), .QN(Q1[3]) );
  DFFSX1 U0_Q1_i_reg_4_ ( .D(n3487), .CK(clk), .SN(rst_n), .QN(Q1[4]) );
  DFFSX1 U0_Q1_i_reg_5_ ( .D(n3486), .CK(clk), .SN(rst_n), .QN(Q1[5]) );
  DFFSX1 U0_Q1_i_reg_6_ ( .D(n3485), .CK(clk), .SN(rst_n), .QN(Q1[6]) );
  DFFSX1 U0_Q1_i_reg_7_ ( .D(n3484), .CK(clk), .SN(rst_n), .QN(Q1[7]) );
  DFFSX1 U0_Q1_i_reg_8_ ( .D(n3483), .CK(clk), .SN(rst_n), .QN(Q1[8]) );
  DFFSX1 U0_Q1_i_reg_9_ ( .D(n3482), .CK(clk), .SN(rst_n), .QN(Q1[9]) );
  DFFSX1 U0_Q1_i_reg_10_ ( .D(n3481), .CK(clk), .SN(rst_n), .QN(Q1[10]) );
  DFFSX1 U0_Q1_i_reg_11_ ( .D(n3480), .CK(clk), .SN(rst_n), .QN(Q1[11]) );
  DFFSX1 U0_Q1_i_reg_12_ ( .D(n3479), .CK(clk), .SN(rst_n), .QN(Q1[12]) );
  DFFSX1 U0_Q1_i_reg_13_ ( .D(n3478), .CK(clk), .SN(rst_n), .QN(Q1[13]) );
  DFFSX1 U0_Q1_i_reg_14_ ( .D(n3477), .CK(clk), .SN(rst_n), .QN(Q1[14]) );
  DFFSX1 U0_Q1_i_reg_15_ ( .D(n3476), .CK(clk), .SN(rst_n), .QN(Q1[15]) );
  DFFSX1 U0_Q1_i_reg_16_ ( .D(n3475), .CK(clk), .SN(rst_n), .QN(Q1[16]) );
  DFFSX1 U0_Q1_i_reg_17_ ( .D(n3474), .CK(clk), .SN(rst_n), .QN(Q1[17]) );
  DFFSX1 U0_Q1_i_reg_18_ ( .D(n3473), .CK(clk), .SN(rst_n), .QN(Q1[18]) );
  DFFSX1 U0_Q1_i_reg_19_ ( .D(n3472), .CK(clk), .SN(rst_n), .QN(Q1[19]) );
  DFFSX1 U0_Q1_i_reg_20_ ( .D(n3471), .CK(clk), .SN(rst_n), .QN(Q1[20]) );
  DFFSX1 U0_Q1_i_reg_21_ ( .D(n3470), .CK(clk), .SN(rst_n), .QN(Q1[21]) );
  DFFSX1 U0_Q1_i_reg_22_ ( .D(n3469), .CK(clk), .SN(rst_n), .QN(Q1[22]) );
  DFFSX1 U0_Q1_i_reg_23_ ( .D(n3468), .CK(clk), .SN(rst_n), .QN(Q1[23]) );
  DFFSX1 U0_Q1_i_reg_24_ ( .D(n3467), .CK(clk), .SN(rst_n), .QN(Q1[24]) );
  DFFSX1 U0_Q1_i_reg_25_ ( .D(n3466), .CK(clk), .SN(rst_n), .QN(Q1[25]) );
  DFFSX1 U0_Q2_r_reg_0_ ( .D(n3465), .CK(clk), .SN(rst_n), .QN(Q2[28]) );
  DFFSX1 U0_Q2_r_reg_1_ ( .D(n3464), .CK(clk), .SN(rst_n), .QN(Q2[29]) );
  DFFSX1 U0_Q2_r_reg_2_ ( .D(n3463), .CK(clk), .SN(rst_n), .QN(Q2[30]) );
  DFFSX1 U0_Q2_r_reg_3_ ( .D(n3462), .CK(clk), .SN(rst_n), .QN(Q2[31]) );
  DFFSX1 U0_Q2_r_reg_4_ ( .D(n3461), .CK(clk), .SN(rst_n), .QN(Q2[32]) );
  DFFSX1 U0_Q2_r_reg_5_ ( .D(n3460), .CK(clk), .SN(rst_n), .QN(Q2[33]) );
  DFFSX1 U0_Q2_r_reg_6_ ( .D(n3459), .CK(clk), .SN(rst_n), .QN(Q2[34]) );
  DFFSX1 U0_Q2_r_reg_7_ ( .D(n3458), .CK(clk), .SN(rst_n), .QN(Q2[35]) );
  DFFSX1 U0_Q2_r_reg_8_ ( .D(n3457), .CK(clk), .SN(rst_n), .QN(Q2[36]) );
  DFFSX1 U0_Q2_r_reg_9_ ( .D(n3456), .CK(clk), .SN(rst_n), .QN(Q2[37]) );
  DFFSX1 U0_Q2_r_reg_10_ ( .D(n3455), .CK(clk), .SN(rst_n), .QN(Q2[38]) );
  DFFSX1 U0_Q2_r_reg_11_ ( .D(n3454), .CK(clk), .SN(rst_n), .QN(Q2[39]) );
  DFFSX1 U0_Q2_r_reg_12_ ( .D(n3453), .CK(clk), .SN(rst_n), .QN(Q2[40]) );
  DFFSX1 U0_Q0_r_reg_1_ ( .D(n3452), .CK(clk), .SN(rst_n), .QN(Q0[29]) );
  DFFSX1 U0_Q0_r_reg_3_ ( .D(n3451), .CK(clk), .SN(rst_n), .QN(Q0[31]) );
  DFFSX1 U0_Q0_r_reg_4_ ( .D(n3450), .CK(clk), .SN(rst_n), .QN(Q0[32]) );
  DFFSX1 U0_Q0_r_reg_5_ ( .D(n3449), .CK(clk), .SN(rst_n), .QN(Q0[33]) );
  DFFSX1 U0_Q0_r_reg_6_ ( .D(n3448), .CK(clk), .SN(rst_n), .QN(Q0[34]) );
  DFFSX1 U0_Q0_r_reg_7_ ( .D(n3447), .CK(clk), .SN(rst_n), .QN(Q0[35]) );
  DFFSX1 U0_Q0_r_reg_8_ ( .D(n3446), .CK(clk), .SN(rst_n), .QN(Q0[36]) );
  DFFSX1 U0_Q0_r_reg_9_ ( .D(n3445), .CK(clk), .SN(rst_n), .QN(Q0[37]) );
  DFFSX1 U0_Q0_r_reg_10_ ( .D(n3444), .CK(clk), .SN(rst_n), .QN(Q0[38]) );
  DFFSX1 U0_Q0_r_reg_11_ ( .D(n3443), .CK(clk), .SN(rst_n), .QN(Q0[39]) );
  DFFSX1 U0_Q0_r_reg_12_ ( .D(n3442), .CK(clk), .SN(rst_n), .QN(Q0[40]) );
  DFFSX1 U0_Q0_r_reg_13_ ( .D(n3441), .CK(clk), .SN(rst_n), .QN(Q0[41]) );
  DFFSX1 U0_Q0_r_reg_14_ ( .D(n3440), .CK(clk), .SN(rst_n), .QN(Q0[42]) );
  DFFSX1 U0_Q0_r_reg_15_ ( .D(n3439), .CK(clk), .SN(rst_n), .QN(Q0[43]) );
  DFFSX1 U0_Q0_r_reg_16_ ( .D(n3438), .CK(clk), .SN(rst_n), .QN(Q0[44]) );
  DFFSX1 U0_Q0_r_reg_17_ ( .D(n3437), .CK(clk), .SN(rst_n), .QN(Q0[45]) );
  DFFSX1 U0_Q0_r_reg_18_ ( .D(n3436), .CK(clk), .SN(rst_n), .QN(Q0[46]) );
  DFFSX1 U0_Q0_r_reg_19_ ( .D(n3435), .CK(clk), .SN(rst_n), .QN(Q0[47]) );
  DFFSX1 U0_Q0_r_reg_20_ ( .D(n3434), .CK(clk), .SN(rst_n), .QN(Q0[48]) );
  DFFSX1 U0_Q0_r_reg_21_ ( .D(n3433), .CK(clk), .SN(rst_n), .QN(Q0[49]) );
  DFFSX1 U0_Q0_r_reg_22_ ( .D(n3432), .CK(clk), .SN(rst_n), .QN(Q0[50]) );
  DFFSX1 U0_Q0_r_reg_23_ ( .D(n3431), .CK(clk), .SN(rst_n), .QN(Q0[51]) );
  DFFSX1 U0_Q0_r_reg_24_ ( .D(n3430), .CK(clk), .SN(rst_n), .QN(Q0[52]) );
  DFFSX1 U0_Q0_r_reg_25_ ( .D(n3429), .CK(clk), .SN(rst_n), .QN(Q0[53]) );
  DFFSX1 U0_Q0_r_reg_2_ ( .D(n3428), .CK(clk), .SN(rst_n), .QN(Q0[30]) );
  DFFSX1 R7_A_reg_9_ ( .D(n3427), .CK(clk), .SN(rst_n), .Q(n29088), .QN(
        AOPA[9]) );
  DFFSX1 R7_A_reg_8_ ( .D(n3423), .CK(clk), .SN(rst_n), .Q(n29087), .QN(
        AOPA[8]) );
  DFFSX4 R7_C_reg_8_ ( .D(n3421), .CK(clk), .SN(rst_n), .Q(n8062), .QN(AOPC[8]) );
  DFFSX4 R7_B_reg_8_ ( .D(n3420), .CK(clk), .SN(rst_n), .Q(n8064), .QN(AOPB[8]) );
  DFFSX1 R7_A_reg_7_ ( .D(n3419), .CK(clk), .SN(rst_n), .Q(n29086), .QN(
        AOPA[7]) );
  DFFSX2 R7_C_reg_7_ ( .D(n3417), .CK(clk), .SN(rst_n), .Q(n7056), .QN(AOPC[7]) );
  DFFSX1 R7_A_reg_6_ ( .D(n3415), .CK(clk), .SN(rst_n), .Q(n29085), .QN(
        AOPA[6]) );
  DFFSX2 R7_B_reg_6_ ( .D(n3412), .CK(clk), .SN(rst_n), .Q(n8069), .QN(AOPB[6]) );
  DFFSX1 R7_A_reg_5_ ( .D(n3411), .CK(clk), .SN(rst_n), .Q(n29084), .QN(
        AOPA[5]) );
  DFFSX2 R7_C_reg_5_ ( .D(n3409), .CK(clk), .SN(rst_n), .Q(n8070), .QN(AOPC[5]) );
  DFFSX1 R7_A_reg_51_ ( .D(n3407), .CK(clk), .SN(rst_n), .Q(n29083), .QN(
        AOPA[51]) );
  DFFSX1 R7_D_reg_51_ ( .D(n3406), .CK(clk), .SN(rst_n), .Q(n8056), .QN(
        AOPD[51]) );
  DFFSX1 R7_C_reg_51_ ( .D(n3405), .CK(clk), .SN(rst_n), .Q(n8055), .QN(
        AOPC[51]) );
  DFFSX1 R7_B_reg_51_ ( .D(n3404), .CK(clk), .SN(rst_n), .Q(n8073), .QN(
        AOPB[51]) );
  DFFSX1 R7_A_reg_50_ ( .D(n3403), .CK(clk), .SN(rst_n), .Q(n29082), .QN(
        AOPA[50]) );
  DFFSX1 R7_D_reg_50_ ( .D(n3402), .CK(clk), .SN(rst_n), .QN(AOPD[50]) );
  DFFSX1 R7_C_reg_50_ ( .D(n3401), .CK(clk), .SN(rst_n), .QN(AOPC[50]) );
  DFFSX1 R7_B_reg_50_ ( .D(n3400), .CK(clk), .SN(rst_n), .QN(AOPB[50]) );
  DFFSX1 R7_A_reg_4_ ( .D(n3399), .CK(clk), .SN(rst_n), .Q(n29081), .QN(
        AOPA[4]) );
  DFFSX2 R7_C_reg_4_ ( .D(n3397), .CK(clk), .SN(rst_n), .Q(n8074), .QN(AOPC[4]) );
  DFFSX2 R7_B_reg_4_ ( .D(n3396), .CK(clk), .SN(rst_n), .Q(n8076), .QN(AOPB[4]) );
  DFFSX1 R7_A_reg_49_ ( .D(n3395), .CK(clk), .SN(rst_n), .Q(n29080), .QN(
        AOPA[49]) );
  DFFSX1 R7_D_reg_49_ ( .D(n3394), .CK(clk), .SN(rst_n), .QN(AOPD[49]) );
  DFFSX1 R7_C_reg_49_ ( .D(n3393), .CK(clk), .SN(rst_n), .QN(AOPC[49]) );
  DFFSX1 R7_B_reg_49_ ( .D(n3392), .CK(clk), .SN(rst_n), .QN(AOPB[49]) );
  DFFSX1 R7_A_reg_48_ ( .D(n3391), .CK(clk), .SN(rst_n), .Q(n29079), .QN(
        AOPA[48]) );
  DFFSX1 R7_D_reg_48_ ( .D(n3390), .CK(clk), .SN(rst_n), .QN(AOPD[48]) );
  DFFSX1 R7_C_reg_48_ ( .D(n3389), .CK(clk), .SN(rst_n), .QN(AOPC[48]) );
  DFFSX1 R7_B_reg_48_ ( .D(n3388), .CK(clk), .SN(rst_n), .QN(AOPB[48]) );
  DFFSX1 R7_A_reg_47_ ( .D(n3387), .CK(clk), .SN(rst_n), .Q(n29078), .QN(
        AOPA[47]) );
  DFFSX1 R7_D_reg_47_ ( .D(n3386), .CK(clk), .SN(rst_n), .QN(AOPD[47]) );
  DFFSX1 R7_C_reg_47_ ( .D(n3385), .CK(clk), .SN(rst_n), .QN(AOPC[47]) );
  DFFSX1 R7_B_reg_47_ ( .D(n3384), .CK(clk), .SN(rst_n), .QN(AOPB[47]) );
  DFFSX1 R7_A_reg_46_ ( .D(n3383), .CK(clk), .SN(rst_n), .Q(n29077), .QN(
        AOPA[46]) );
  DFFSX1 R7_D_reg_46_ ( .D(n3382), .CK(clk), .SN(rst_n), .QN(AOPD[46]) );
  DFFSX1 R7_C_reg_46_ ( .D(n3381), .CK(clk), .SN(rst_n), .QN(AOPC[46]) );
  DFFSX1 R7_B_reg_46_ ( .D(n3380), .CK(clk), .SN(rst_n), .QN(AOPB[46]) );
  DFFSX1 R7_A_reg_45_ ( .D(n3379), .CK(clk), .SN(rst_n), .Q(n29076), .QN(
        AOPA[45]) );
  DFFSX1 R7_C_reg_45_ ( .D(n3377), .CK(clk), .SN(rst_n), .QN(AOPC[45]) );
  DFFSX1 R7_B_reg_45_ ( .D(n3376), .CK(clk), .SN(rst_n), .QN(AOPB[45]) );
  DFFSX1 R7_A_reg_44_ ( .D(n3375), .CK(clk), .SN(rst_n), .Q(n29075), .QN(
        AOPA[44]) );
  DFFSX1 R7_C_reg_44_ ( .D(n3373), .CK(clk), .SN(rst_n), .QN(AOPC[44]) );
  DFFSX1 R7_B_reg_44_ ( .D(n3372), .CK(clk), .SN(rst_n), .QN(AOPB[44]) );
  DFFSX1 R7_A_reg_43_ ( .D(n3371), .CK(clk), .SN(rst_n), .Q(n29074), .QN(
        AOPA[43]) );
  DFFSX1 R7_A_reg_42_ ( .D(n3367), .CK(clk), .SN(rst_n), .Q(n29073), .QN(
        AOPA[42]) );
  DFFSX1 R7_A_reg_41_ ( .D(n3363), .CK(clk), .SN(rst_n), .Q(n29072), .QN(
        AOPA[41]) );
  DFFSX1 R7_D_reg_41_ ( .D(n3362), .CK(clk), .SN(rst_n), .QN(AOPD[41]) );
  DFFSX1 R7_A_reg_40_ ( .D(n3359), .CK(clk), .SN(rst_n), .Q(n29071), .QN(
        AOPA[40]) );
  DFFSX1 R7_B_reg_40_ ( .D(n3356), .CK(clk), .SN(rst_n), .QN(AOPB[40]) );
  DFFSX1 R7_A_reg_3_ ( .D(n3355), .CK(clk), .SN(rst_n), .Q(n29070), .QN(
        AOPA[3]) );
  DFFSX4 R7_D_reg_3_ ( .D(n3354), .CK(clk), .SN(rst_n), .Q(n8080), .QN(AOPD[3]) );
  DFFSX1 R7_A_reg_39_ ( .D(n3351), .CK(clk), .SN(rst_n), .Q(n29069), .QN(
        AOPA[39]) );
  DFFSX2 R7_D_reg_39_ ( .D(n3350), .CK(clk), .SN(rst_n), .QN(AOPD[39]) );
  DFFSX2 R7_B_reg_39_ ( .D(n3348), .CK(clk), .SN(rst_n), .QN(AOPB[39]) );
  DFFSX1 R7_A_reg_38_ ( .D(n3347), .CK(clk), .SN(rst_n), .Q(n29068), .QN(
        AOPA[38]) );
  DFFSX2 R7_D_reg_38_ ( .D(n3346), .CK(clk), .SN(rst_n), .QN(AOPD[38]) );
  DFFSX2 R7_B_reg_38_ ( .D(n3344), .CK(clk), .SN(rst_n), .QN(AOPB[38]) );
  DFFSX1 R7_A_reg_37_ ( .D(n3343), .CK(clk), .SN(rst_n), .Q(n29067), .QN(
        AOPA[37]) );
  DFFSX2 R7_C_reg_37_ ( .D(n3341), .CK(clk), .SN(rst_n), .QN(AOPC[37]) );
  DFFSX2 R7_B_reg_37_ ( .D(n3340), .CK(clk), .SN(rst_n), .QN(AOPB[37]) );
  DFFSX1 R7_A_reg_36_ ( .D(n3339), .CK(clk), .SN(rst_n), .Q(n29066), .QN(
        AOPA[36]) );
  DFFSX1 R7_D_reg_36_ ( .D(n3338), .CK(clk), .SN(rst_n), .QN(AOPD[36]) );
  DFFSX2 R7_C_reg_36_ ( .D(n3337), .CK(clk), .SN(rst_n), .QN(AOPC[36]) );
  DFFSX1 R7_A_reg_35_ ( .D(n3335), .CK(clk), .SN(rst_n), .Q(n29065), .QN(
        AOPA[35]) );
  DFFSX2 R7_D_reg_35_ ( .D(n3334), .CK(clk), .SN(rst_n), .QN(AOPD[35]) );
  DFFSX1 R7_A_reg_34_ ( .D(n3331), .CK(clk), .SN(rst_n), .Q(n29064), .QN(
        AOPA[34]) );
  DFFSX2 R7_B_reg_34_ ( .D(n3328), .CK(clk), .SN(rst_n), .QN(AOPB[34]) );
  DFFSX1 R7_A_reg_33_ ( .D(n3327), .CK(clk), .SN(rst_n), .Q(n29063), .QN(
        AOPA[33]) );
  DFFSX1 R7_A_reg_32_ ( .D(n3323), .CK(clk), .SN(rst_n), .Q(n29062), .QN(
        AOPA[32]) );
  DFFSX1 R7_A_reg_31_ ( .D(n3319), .CK(clk), .SN(rst_n), .Q(n29061), .QN(
        AOPA[31]) );
  DFFSX1 R7_A_reg_30_ ( .D(n3315), .CK(clk), .SN(rst_n), .Q(n29060), .QN(
        AOPA[30]) );
  DFFSX1 R7_A_reg_2_ ( .D(n3311), .CK(clk), .SN(rst_n), .Q(n29059), .QN(
        AOPA[2]) );
  DFFSX4 R7_D_reg_2_ ( .D(n3310), .CK(clk), .SN(rst_n), .Q(n5777), .QN(AOPD[2]) );
  DFFSX4 R7_C_reg_2_ ( .D(n3309), .CK(clk), .SN(rst_n), .Q(n8084), .QN(AOPC[2]) );
  DFFSX1 R7_A_reg_29_ ( .D(n3307), .CK(clk), .SN(rst_n), .Q(n29058), .QN(
        AOPA[29]) );
  DFFSX2 R7_D_reg_29_ ( .D(n3306), .CK(clk), .SN(rst_n), .QN(AOPD[29]) );
  DFFSX2 R7_C_reg_29_ ( .D(n3305), .CK(clk), .SN(rst_n), .QN(AOPC[29]) );
  DFFSX2 R7_B_reg_29_ ( .D(n3304), .CK(clk), .SN(rst_n), .QN(AOPB[29]) );
  DFFSX1 R7_A_reg_28_ ( .D(n3303), .CK(clk), .SN(rst_n), .Q(n29057), .QN(
        AOPA[28]) );
  DFFSX2 R7_D_reg_28_ ( .D(n3302), .CK(clk), .SN(rst_n), .QN(AOPD[28]) );
  DFFSX2 R7_C_reg_28_ ( .D(n3301), .CK(clk), .SN(rst_n), .QN(AOPC[28]) );
  DFFSX2 R7_B_reg_28_ ( .D(n3300), .CK(clk), .SN(rst_n), .QN(AOPB[28]) );
  DFFSX1 R7_A_reg_27_ ( .D(n3299), .CK(clk), .SN(rst_n), .Q(n29056), .QN(
        AOPA[27]) );
  DFFSX2 R7_D_reg_27_ ( .D(n3298), .CK(clk), .SN(rst_n), .QN(AOPD[27]) );
  DFFSX2 R7_C_reg_27_ ( .D(n3297), .CK(clk), .SN(rst_n), .QN(AOPC[27]) );
  DFFSX1 R7_A_reg_26_ ( .D(n3295), .CK(clk), .SN(rst_n), .Q(n29055), .QN(
        AOPA[26]) );
  DFFSX2 R7_D_reg_26_ ( .D(n3294), .CK(clk), .SN(rst_n), .QN(AOPD[26]) );
  DFFSX2 R7_C_reg_26_ ( .D(n3293), .CK(clk), .SN(rst_n), .QN(AOPC[26]) );
  DFFSX1 R7_A_reg_25_ ( .D(n3291), .CK(clk), .SN(rst_n), .Q(n29054), .QN(
        AOPA[25]) );
  DFFSX1 R7_D_reg_25_ ( .D(n3290), .CK(clk), .SN(rst_n), .QN(AOPD[25]) );
  DFFSX1 R7_C_reg_25_ ( .D(n3289), .CK(clk), .SN(rst_n), .QN(AOPC[25]) );
  DFFSX1 R7_B_reg_25_ ( .D(n3288), .CK(clk), .SN(rst_n), .QN(AOPB[25]) );
  DFFSX1 R7_A_reg_24_ ( .D(n3287), .CK(clk), .SN(rst_n), .Q(n29053), .QN(
        AOPA[24]) );
  DFFSX1 R7_D_reg_24_ ( .D(n3286), .CK(clk), .SN(rst_n), .Q(n8088), .QN(
        AOPD[24]) );
  DFFSX1 R7_C_reg_24_ ( .D(n3285), .CK(clk), .SN(rst_n), .Q(n8087), .QN(
        AOPC[24]) );
  DFFSX1 R7_B_reg_24_ ( .D(n3284), .CK(clk), .SN(rst_n), .Q(n8089), .QN(
        AOPB[24]) );
  DFFSX1 R7_A_reg_23_ ( .D(n3283), .CK(clk), .SN(rst_n), .Q(n29052), .QN(
        AOPA[23]) );
  DFFSX1 R7_D_reg_23_ ( .D(n3282), .CK(clk), .SN(rst_n), .Q(n8091), .QN(
        AOPD[23]) );
  DFFSX1 R7_C_reg_23_ ( .D(n3281), .CK(clk), .SN(rst_n), .Q(n8090), .QN(
        AOPC[23]) );
  DFFSX1 R7_B_reg_23_ ( .D(n3280), .CK(clk), .SN(rst_n), .Q(n8092), .QN(
        AOPB[23]) );
  DFFSX1 R7_A_reg_22_ ( .D(n3279), .CK(clk), .SN(rst_n), .Q(n29051), .QN(
        AOPA[22]) );
  DFFSX1 R7_D_reg_22_ ( .D(n3278), .CK(clk), .SN(rst_n), .Q(n8094), .QN(
        AOPD[22]) );
  DFFSX1 R7_C_reg_22_ ( .D(n3277), .CK(clk), .SN(rst_n), .Q(n8093), .QN(
        AOPC[22]) );
  DFFSX1 R7_B_reg_22_ ( .D(n3276), .CK(clk), .SN(rst_n), .Q(n8095), .QN(
        AOPB[22]) );
  DFFSX1 R7_A_reg_21_ ( .D(n3275), .CK(clk), .SN(rst_n), .Q(n29050), .QN(
        AOPA[21]) );
  DFFSX1 R7_A_reg_20_ ( .D(n3271), .CK(clk), .SN(rst_n), .Q(n29049), .QN(
        AOPA[20]) );
  DFFSX1 R7_D_reg_20_ ( .D(n3270), .CK(clk), .SN(rst_n), .Q(n8100), .QN(
        AOPD[20]) );
  DFFSX1 R7_C_reg_20_ ( .D(n3269), .CK(clk), .SN(rst_n), .Q(n8099), .QN(
        AOPC[20]) );
  DFFSX1 R7_B_reg_20_ ( .D(n3268), .CK(clk), .SN(rst_n), .Q(n8101), .QN(
        AOPB[20]) );
  DFFSX1 R7_A_reg_1_ ( .D(n3267), .CK(clk), .SN(rst_n), .Q(n29048), .QN(
        AOPA[1]) );
  DFFSX4 R7_B_reg_1_ ( .D(n3264), .CK(clk), .SN(rst_n), .Q(n8104), .QN(AOPB[1]) );
  DFFSX1 R7_A_reg_19_ ( .D(n3263), .CK(clk), .SN(rst_n), .Q(n29047), .QN(
        AOPA[19]) );
  DFFSX1 R7_A_reg_18_ ( .D(n3259), .CK(clk), .SN(rst_n), .Q(n29046), .QN(
        AOPA[18]) );
  DFFSX1 R7_A_reg_17_ ( .D(n3255), .CK(clk), .SN(rst_n), .Q(n29045), .QN(
        AOPA[17]) );
  DFFSX1 R7_A_reg_16_ ( .D(n3251), .CK(clk), .SN(rst_n), .Q(n29044), .QN(
        AOPA[16]) );
  DFFSX1 R7_A_reg_15_ ( .D(n3247), .CK(clk), .SN(rst_n), .Q(n29043), .QN(
        AOPA[15]) );
  DFFSX1 R7_A_reg_14_ ( .D(n3243), .CK(clk), .SN(rst_n), .Q(n29042), .QN(
        AOPA[14]) );
  DFFSX2 R7_B_reg_14_ ( .D(n3240), .CK(clk), .SN(rst_n), .Q(n7990), .QN(
        AOPB[14]) );
  DFFSX1 R7_A_reg_13_ ( .D(n3239), .CK(clk), .SN(rst_n), .Q(n29041), .QN(
        AOPA[13]) );
  DFFSX1 R7_A_reg_12_ ( .D(n3235), .CK(clk), .SN(rst_n), .Q(n29040), .QN(
        AOPA[12]) );
  DFFSX2 R7_C_reg_12_ ( .D(n3233), .CK(clk), .SN(rst_n), .Q(n7062), .QN(
        AOPC[12]) );
  DFFSX1 R7_A_reg_11_ ( .D(n3231), .CK(clk), .SN(rst_n), .Q(n29039), .QN(
        AOPA[11]) );
  DFFSX1 R7_A_reg_10_ ( .D(n3227), .CK(clk), .SN(rst_n), .Q(n29038), .QN(
        AOPA[10]) );
  DFFSX2 R7_D_reg_10_ ( .D(n3226), .CK(clk), .SN(rst_n), .Q(n8204), .QN(
        AOPD[10]) );
  DFFSX1 R7_A_reg_0_ ( .D(n3223), .CK(clk), .SN(rst_n), .Q(n29037), .QN(
        AOPA[0]) );
  DFFSX4 R7_D_reg_0_ ( .D(n3222), .CK(clk), .SN(rst_n), .Q(n8207), .QN(AOPD[0]) );
  DFFSX4 R7_B_reg_0_ ( .D(n3220), .CK(clk), .SN(rst_n), .Q(n8208), .QN(AOPB[0]) );
  FFT2048_DW02_mult_2_stage_J1_0 U0_U0_A2_U0 ( .A(AOPB[25:0]), .B({U0_U0_z2, 
        n12003, U0_U0_z1[0]}), .TC(1'b1), .CLK(clk), .PRODUCT({
        SYNOPSYS_UNCONNECTED_417, SYNOPSYS_UNCONNECTED_418, U0_U0_y2}) );
  FFT2048_DW02_mult_2_stage_J1_1 U0_U1_A1_U0 ( .A(AOPC[51:26]), .B({
        U1_U1_z1[16:6], n5766, U1_U1_z1[4:2], n29097, U1_U1_z1[0]}), .TC(1'b1), 
        .CLK(clk), .PRODUCT({SYNOPSYS_UNCONNECTED_419, 
        SYNOPSYS_UNCONNECTED_420, U0_U1_y1}) );
  FFT2048_DW02_mult_2_stage_J1_2 U0_U1_A2_U0 ( .A(AOPC[25:0]), .B({
        U1_U1_z2[16], n6902, U1_U1_z2[14:11], n6909, U1_U1_z2[9:4], n6877, 
        U1_U1_z2[2:1], U1_U1_z1[0]}), .TC(1'b1), .CLK(clk), .PRODUCT({
        SYNOPSYS_UNCONNECTED_421, SYNOPSYS_UNCONNECTED_422, U0_U1_y2}) );
  FFT2048_DW02_mult_2_stage_J1_3 U0_U2_A1_U0 ( .A(AOPD[51:26]), .B({
        U1_U2_z1[16:2], n29098, U1_U2_z1[0]}), .TC(1'b1), .CLK(clk), .PRODUCT(
        {SYNOPSYS_UNCONNECTED_423, SYNOPSYS_UNCONNECTED_424, U0_U2_y1}) );
  FFT2048_DW02_mult_2_stage_J1_4 U0_U2_A2_U0 ( .A(AOPD[25:0]), .B({
        U1_U2_z2[16:10], n5771, U1_U2_z2[8:1], U1_U2_z1[0]}), .TC(1'b1), .CLK(
        clk), .PRODUCT({SYNOPSYS_UNCONNECTED_425, SYNOPSYS_UNCONNECTED_426, 
        U0_U2_y2}) );
  FFT2048_DW02_mult_2_stage_J1_5 U1_U0_A1_U0 ( .A(BOPB[51:26]), .B({
        U0_U0_z1[16], n6945, U0_U0_z1[14:2], n6879, U0_U0_z1[0]}), .TC(1'b1), 
        .CLK(clk), .PRODUCT({SYNOPSYS_UNCONNECTED_427, 
        SYNOPSYS_UNCONNECTED_428, U1_U0_y1}) );
  FFT2048_DW02_mult_2_stage_J1_6 U1_U0_A2_U0 ( .A(BOPB[25:0]), .B({U0_U0_z2, 
        n12003, U0_U0_z1[0]}), .TC(1'b1), .CLK(clk), .PRODUCT({
        SYNOPSYS_UNCONNECTED_429, SYNOPSYS_UNCONNECTED_430, U1_U0_y2}) );
  FFT2048_DW02_mult_2_stage_J1_7 U1_U1_A1_U0 ( .A(BOPC[51:26]), .B({
        U1_U1_z1[16:6], n5766, U1_U1_z1[4:2], n29097, U1_U1_z1[0]}), .TC(1'b1), 
        .CLK(clk), .PRODUCT({SYNOPSYS_UNCONNECTED_431, 
        SYNOPSYS_UNCONNECTED_432, U1_U1_y1}) );
  FFT2048_DW02_mult_2_stage_J1_8 U1_U1_A2_U0 ( .A(BOPC[25:0]), .B({
        U1_U1_z2[16], n6902, U1_U1_z2[14:11], n6909, U1_U1_z2[9:4], n6877, 
        U1_U1_z2[2:1], U1_U1_z1[0]}), .TC(1'b1), .CLK(clk), .PRODUCT({
        SYNOPSYS_UNCONNECTED_433, SYNOPSYS_UNCONNECTED_434, U1_U1_y2}) );
  FFT2048_DW02_mult_2_stage_J1_9 U1_U2_A1_U0 ( .A(BOPD[51:26]), .B({
        U1_U2_z1[16:2], n29098, U1_U2_z1[0]}), .TC(1'b1), .CLK(clk), .PRODUCT(
        {SYNOPSYS_UNCONNECTED_435, SYNOPSYS_UNCONNECTED_436, U1_U2_y1}) );
  FFT2048_DW02_mult_2_stage_J1_10 U1_U2_A2_U0 ( .A(BOPD[25:0]), .B({
        U1_U2_z2[16:10], n5771, U1_U2_z2[8:1], U1_U2_z1[0]}), .TC(1'b1), .CLK(
        clk), .PRODUCT({SYNOPSYS_UNCONNECTED_437, SYNOPSYS_UNCONNECTED_438, 
        U1_U2_y2}) );
  FFT2048_DW02_mult_2_stage_J1_11 U2_U0_A1_U0 ( .A({U2_B_r[25:23], n7118, 
        U2_B_r[21:9], n7130, U2_B_r[7:6], n7088, U2_B_r[4:0]}), .B(U2_U0_z1), 
        .TC(1'b1), .CLK(clk), .PRODUCT({SYNOPSYS_UNCONNECTED_439, 
        SYNOPSYS_UNCONNECTED_440, SYNOPSYS_UNCONNECTED_441, U2_U0_y1}) );
  FFT2048_DW02_mult_2_stage_J1_12 U2_U0_A2_U0 ( .A({U2_B_i[25:4], n29101, 
        U2_B_i[2:0]}), .B({U2_U0_z2, U2_U0_z1[0]}), .TC(1'b1), .CLK(clk), 
        .PRODUCT({SYNOPSYS_UNCONNECTED_442, SYNOPSYS_UNCONNECTED_443, 
        SYNOPSYS_UNCONNECTED_444, U2_U0_y2}) );
  FFT2048_DW02_mult_2_stage_J1_13 U0_U1_A0_U0 ( .A(W1[15:0]), .B(U0_U1_z0), 
        .TC(1'b1), .CLK(clk), .PRODUCT({SYNOPSYS_UNCONNECTED_445, 
        SYNOPSYS_UNCONNECTED_446, U0_U1_y0}) );
  FFT2048_DW02_mult_2_stage_J1_14 U0_U2_A0_U0 ( .A(W2[15:0]), .B(U0_U2_z0), 
        .TC(1'b1), .CLK(clk), .PRODUCT({SYNOPSYS_UNCONNECTED_447, 
        SYNOPSYS_UNCONNECTED_448, U0_U2_y0}) );
  FFT2048_DW02_mult_2_stage_J1_15 U1_U0_A0_U0 ( .A({n6897, W0[14:3], n6876, 
        W0[1:0]}), .B(U1_U0_z0), .TC(1'b1), .CLK(clk), .PRODUCT({
        SYNOPSYS_UNCONNECTED_449, SYNOPSYS_UNCONNECTED_450, U1_U0_y0}) );
  FFT2048_DW02_mult_2_stage_J1_16 U1_U1_A0_U0 ( .A({W1[15:4], n7143, W1[2:0]}), 
        .B(U1_U1_z0), .TC(1'b1), .CLK(clk), .PRODUCT({SYNOPSYS_UNCONNECTED_451, 
        SYNOPSYS_UNCONNECTED_452, U1_U1_y0}) );
  FFT2048_DW02_mult_2_stage_J1_17 U1_U2_A0_U0 ( .A(W2[15:0]), .B(U1_U2_z0), 
        .TC(1'b1), .CLK(clk), .PRODUCT({SYNOPSYS_UNCONNECTED_453, 
        SYNOPSYS_UNCONNECTED_454, U1_U2_y0}) );
  FFT2048_DW02_mult_2_stage_J1_18 U2_U0_A0_U0 ( .A(W3[15:0]), .B({
        U2_U0_z0[26:17], n6889, U2_U0_z0[15:8], n6890, U2_U0_z0[6:0]}), .TC(
        1'b1), .CLK(clk), .PRODUCT({SYNOPSYS_UNCONNECTED_455, 
        SYNOPSYS_UNCONNECTED_456, SYNOPSYS_UNCONNECTED_457, U2_U0_y0}) );
  FFT2048_DW02_mult_2_stage_J1_19 U0_U0_A1_U0 ( .A(AOPB[51:26]), .B({
        U0_U0_z1[16], n6945, U0_U0_z1[14:2], n6879, U0_U0_z1[0]}), .TC(1'b1), 
        .CLK(clk), .PRODUCT({SYNOPSYS_UNCONNECTED_458, 
        SYNOPSYS_UNCONNECTED_459, U0_U0_y1}) );
  FFT2048_DW02_mult_2_stage_J1_20 U0_U0_A0_U0 ( .A({n6897, W0[14:3], n6876, 
        W0[1:0]}), .B(U0_U0_z0), .TC(1'b1), .CLK(clk), .PRODUCT({
        SYNOPSYS_UNCONNECTED_460, SYNOPSYS_UNCONNECTED_461, U0_U0_y0}) );
  DFFSX1 U1_A_r_d0_reg_1_ ( .D(n28682), .CK(clk), .SN(rst_n), .QN(U1_A_r_d0[1]) );
  DFFSX2 T1_W2_reg_15_ ( .D(n29170), .CK(clk), .SN(rst_n), .Q(n8001), .QN(
        W2[15]) );
  DFFSX4 T1_W3_reg_7_ ( .D(n29115), .CK(clk), .SN(rst_n), .Q(n8015), .QN(W3[7]) );
  DFFSX4 R9_A_reg_36_ ( .D(n3755), .CK(clk), .SN(rst_n), .Q(n28748), .QN(
        BOPA[36]) );
  DFFSX4 R9_A_reg_41_ ( .D(n3779), .CK(clk), .SN(rst_n), .Q(n28746), .QN(
        BOPA[41]) );
  DFFSX4 T1_W3_reg_11_ ( .D(n29142), .CK(clk), .SN(rst_n), .Q(n8018), .QN(
        W3[11]) );
  DFFSX4 R9_A_reg_30_ ( .D(n3731), .CK(clk), .SN(rst_n), .Q(n29104), .QN(
        BOPA[30]) );
  DFFSX1 C_sel_reg_reg_0__0_ ( .D(n5412), .CK(clk), .SN(rst_n), .Q(n28707), 
        .QN(C_sel_reg[0]) );
  DFFSX4 R9_A_reg_40_ ( .D(n3775), .CK(clk), .SN(rst_n), .Q(n28683), .QN(
        BOPA[40]) );
  DFFSX1 cnt_reg_3_ ( .D(n5676), .CK(clk), .SN(rst_n), .Q(n28679), .QN(cnt[3])
         );
  DFFSX1 cnt_reg_5_ ( .D(n5674), .CK(clk), .SN(rst_n), .Q(n28673), .QN(cnt[5])
         );
  DFFSX1 U1_pipe2_reg_26_ ( .D(n5038), .CK(clk), .SN(rst_n), .QN(U1_pipe2[26])
         );
  DFFSX1 U1_pipe0_reg_26_ ( .D(n5129), .CK(clk), .SN(rst_n), .QN(U1_pipe0[26])
         );
  DFFSX1 U1_pipe14_reg_26_ ( .D(n4777), .CK(clk), .SN(rst_n), .QN(
        U1_pipe14[26]) );
  DFFSX1 U1_pipe4_reg_26_ ( .D(n5094), .CK(clk), .SN(rst_n), .QN(U1_pipe4[26])
         );
  DFFSX1 U1_pipe10_reg_26_ ( .D(n4864), .CK(clk), .SN(rst_n), .QN(
        U1_pipe10[26]) );
  DFFSX1 U1_pipe2_reg_24_ ( .D(n5036), .CK(clk), .SN(rst_n), .QN(U1_pipe2[24])
         );
  DFFSX1 U1_pipe10_reg_25_ ( .D(n4863), .CK(clk), .SN(rst_n), .QN(
        U1_pipe10[25]) );
  DFFSX1 U1_pipe10_reg_24_ ( .D(n4862), .CK(clk), .SN(rst_n), .QN(
        U1_pipe10[24]) );
  DFFSX1 U1_pipe2_reg_25_ ( .D(n5037), .CK(clk), .SN(rst_n), .QN(U1_pipe2[25])
         );
  DFFSX1 U1_pipe2_reg_23_ ( .D(n5035), .CK(clk), .SN(rst_n), .QN(U1_pipe2[23])
         );
  DFFSX1 U1_pipe2_reg_22_ ( .D(n5034), .CK(clk), .SN(rst_n), .QN(U1_pipe2[22])
         );
  DFFSX1 U1_pipe14_reg_25_ ( .D(n4776), .CK(clk), .SN(rst_n), .QN(
        U1_pipe14[25]) );
  DFFSX1 U1_pipe14_reg_23_ ( .D(n4774), .CK(clk), .SN(rst_n), .QN(
        U1_pipe14[23]) );
  DFFSX1 U1_pipe14_reg_22_ ( .D(n4773), .CK(clk), .SN(rst_n), .QN(
        U1_pipe14[22]) );
  DFFSX1 U1_pipe10_reg_23_ ( .D(n4861), .CK(clk), .SN(rst_n), .QN(
        U1_pipe10[23]) );
  DFFSX1 U1_pipe10_reg_22_ ( .D(n4860), .CK(clk), .SN(rst_n), .QN(
        U1_pipe10[22]) );
  DFFSX1 U1_pipe10_reg_21_ ( .D(n4859), .CK(clk), .SN(rst_n), .QN(
        U1_pipe10[21]) );
  DFFSX1 out_valid_reg ( .D(n28700), .CK(clk), .SN(rst_n), .QN(out_valid) );
  DFFSX1 O_im_reg_9_ ( .D(n5739), .CK(clk), .SN(rst_n), .QN(O_im[9]) );
  DFFSX1 O_im_reg_8_ ( .D(n5740), .CK(clk), .SN(rst_n), .QN(O_im[8]) );
  DFFSX1 O_im_reg_7_ ( .D(n5741), .CK(clk), .SN(rst_n), .QN(O_im[7]) );
  DFFSX1 O_im_reg_6_ ( .D(n5742), .CK(clk), .SN(rst_n), .QN(O_im[6]) );
  DFFSX1 O_im_reg_5_ ( .D(n5743), .CK(clk), .SN(rst_n), .QN(O_im[5]) );
  DFFSX1 O_re_reg_25_ ( .D(n5697), .CK(clk), .SN(rst_n), .QN(O_re[25]) );
  DFFSX1 O_re_reg_24_ ( .D(n5698), .CK(clk), .SN(rst_n), .QN(O_re[24]) );
  DFFSX1 O_im_reg_4_ ( .D(n5744), .CK(clk), .SN(rst_n), .QN(O_im[4]) );
  DFFSX1 O_re_reg_23_ ( .D(n5699), .CK(clk), .SN(rst_n), .QN(O_re[23]) );
  DFFSX1 O_re_reg_22_ ( .D(n5700), .CK(clk), .SN(rst_n), .QN(O_re[22]) );
  DFFSX1 O_re_reg_21_ ( .D(n5701), .CK(clk), .SN(rst_n), .QN(O_re[21]) );
  DFFSX1 O_re_reg_20_ ( .D(n5702), .CK(clk), .SN(rst_n), .QN(O_re[20]) );
  DFFSX1 O_re_reg_19_ ( .D(n5703), .CK(clk), .SN(rst_n), .QN(O_re[19]) );
  DFFSX1 O_re_reg_18_ ( .D(n5704), .CK(clk), .SN(rst_n), .QN(O_re[18]) );
  DFFSX1 O_re_reg_17_ ( .D(n5705), .CK(clk), .SN(rst_n), .QN(O_re[17]) );
  DFFSX1 O_re_reg_16_ ( .D(n5706), .CK(clk), .SN(rst_n), .QN(O_re[16]) );
  DFFSX1 O_re_reg_15_ ( .D(n5707), .CK(clk), .SN(rst_n), .QN(O_re[15]) );
  DFFSX1 O_re_reg_14_ ( .D(n5708), .CK(clk), .SN(rst_n), .QN(O_re[14]) );
  DFFSX1 O_im_reg_3_ ( .D(n5745), .CK(clk), .SN(rst_n), .QN(O_im[3]) );
  DFFSX1 O_re_reg_13_ ( .D(n5709), .CK(clk), .SN(rst_n), .QN(O_re[13]) );
  DFFSX1 O_re_reg_12_ ( .D(n5710), .CK(clk), .SN(rst_n), .QN(O_re[12]) );
  DFFSX1 O_re_reg_11_ ( .D(n5711), .CK(clk), .SN(rst_n), .QN(O_re[11]) );
  DFFSX1 O_re_reg_10_ ( .D(n5712), .CK(clk), .SN(rst_n), .QN(O_re[10]) );
  DFFSX1 O_re_reg_9_ ( .D(n5713), .CK(clk), .SN(rst_n), .QN(O_re[9]) );
  DFFSX1 O_re_reg_8_ ( .D(n5714), .CK(clk), .SN(rst_n), .QN(O_re[8]) );
  DFFSX1 O_re_reg_7_ ( .D(n5715), .CK(clk), .SN(rst_n), .QN(O_re[7]) );
  DFFSX1 O_re_reg_6_ ( .D(n5716), .CK(clk), .SN(rst_n), .QN(O_re[6]) );
  DFFSX1 O_re_reg_5_ ( .D(n5717), .CK(clk), .SN(rst_n), .QN(O_re[5]) );
  DFFSX1 O_re_reg_4_ ( .D(n5718), .CK(clk), .SN(rst_n), .QN(O_re[4]) );
  DFFSX1 O_im_reg_2_ ( .D(n5746), .CK(clk), .SN(rst_n), .QN(O_im[2]) );
  DFFSX1 O_re_reg_3_ ( .D(n5719), .CK(clk), .SN(rst_n), .QN(O_re[3]) );
  DFFSX1 O_re_reg_2_ ( .D(n5720), .CK(clk), .SN(rst_n), .QN(O_re[2]) );
  DFFSX1 O_re_reg_1_ ( .D(n5721), .CK(clk), .SN(rst_n), .QN(O_re[1]) );
  DFFSX1 O_re_reg_0_ ( .D(n5722), .CK(clk), .SN(rst_n), .QN(O_re[0]) );
  DFFSX1 O_im_reg_25_ ( .D(n5723), .CK(clk), .SN(rst_n), .QN(O_im[25]) );
  DFFSX1 O_im_reg_24_ ( .D(n5724), .CK(clk), .SN(rst_n), .QN(O_im[24]) );
  DFFSX1 O_im_reg_23_ ( .D(n5725), .CK(clk), .SN(rst_n), .QN(O_im[23]) );
  DFFSX1 O_im_reg_22_ ( .D(n5726), .CK(clk), .SN(rst_n), .QN(O_im[22]) );
  DFFSX1 O_im_reg_21_ ( .D(n5727), .CK(clk), .SN(rst_n), .QN(O_im[21]) );
  DFFSX1 O_im_reg_20_ ( .D(n5728), .CK(clk), .SN(rst_n), .QN(O_im[20]) );
  DFFSX1 O_im_reg_1_ ( .D(n5747), .CK(clk), .SN(rst_n), .QN(O_im[1]) );
  DFFSX1 O_im_reg_19_ ( .D(n5729), .CK(clk), .SN(rst_n), .QN(O_im[19]) );
  DFFSX1 O_im_reg_18_ ( .D(n5730), .CK(clk), .SN(rst_n), .QN(O_im[18]) );
  DFFSX1 O_im_reg_17_ ( .D(n5731), .CK(clk), .SN(rst_n), .QN(O_im[17]) );
  DFFSX1 O_im_reg_16_ ( .D(n5732), .CK(clk), .SN(rst_n), .QN(O_im[16]) );
  DFFSX1 O_im_reg_15_ ( .D(n5733), .CK(clk), .SN(rst_n), .QN(O_im[15]) );
  DFFSX1 O_im_reg_14_ ( .D(n5734), .CK(clk), .SN(rst_n), .QN(O_im[14]) );
  DFFSX1 O_im_reg_13_ ( .D(n5735), .CK(clk), .SN(rst_n), .QN(O_im[13]) );
  DFFSX1 O_im_reg_12_ ( .D(n5736), .CK(clk), .SN(rst_n), .QN(O_im[12]) );
  DFFSX1 O_im_reg_11_ ( .D(n5737), .CK(clk), .SN(rst_n), .QN(O_im[11]) );
  DFFSX1 O_im_reg_10_ ( .D(n5738), .CK(clk), .SN(rst_n), .QN(O_im[10]) );
  DFFSX1 O_im_reg_0_ ( .D(n5748), .CK(clk), .SN(rst_n), .QN(O_im[0]) );
  DFFSX1 R9_A_reg_3_ ( .D(n3771), .CK(clk), .SN(rst_n), .Q(n29032), .QN(
        BOPA[3]) );
  DFFSX1 R9_A_reg_2_ ( .D(n3727), .CK(clk), .SN(rst_n), .Q(n29016), .QN(
        BOPA[2]) );
  DFFSX1 R9_A_reg_1_ ( .D(n3683), .CK(clk), .SN(rst_n), .Q(n29013), .QN(
        BOPA[1]) );
  DFFSX1 R9_A_reg_7_ ( .D(n3835), .CK(clk), .SN(rst_n), .Q(n29034), .QN(
        BOPA[7]) );
  DFFSX1 R9_A_reg_6_ ( .D(n3831), .CK(clk), .SN(rst_n), .Q(n29033), .QN(
        BOPA[6]) );
  DFFSX1 R9_A_reg_5_ ( .D(n3827), .CK(clk), .SN(rst_n), .Q(n29017), .QN(
        BOPA[5]) );
  DFFSX1 R9_A_reg_4_ ( .D(n3815), .CK(clk), .SN(rst_n), .Q(n29011), .QN(
        BOPA[4]) );
  DFFSX4 R9_B_reg_40_ ( .D(n3772), .CK(clk), .SN(rst_n), .QN(BOPB[40]) );
  DFFSX4 R9_D_reg_36_ ( .D(n3754), .CK(clk), .SN(rst_n), .QN(BOPD[36]) );
  DFFSX4 T1_W0_reg_19_ ( .D(n29230), .CK(clk), .SN(rst_n), .QN(W0[19]) );
  DFFSX4 R7_C_reg_39_ ( .D(n3349), .CK(clk), .SN(rst_n), .QN(AOPC[39]) );
  DFFSX2 R7_B_reg_31_ ( .D(n3316), .CK(clk), .SN(rst_n), .QN(AOPB[31]) );
  DFFSX4 T1_W1_reg_18_ ( .D(n29199), .CK(clk), .SN(rst_n), .QN(W1[18]) );
  DFFSX2 R7_C_reg_31_ ( .D(n3317), .CK(clk), .SN(rst_n), .QN(AOPC[31]) );
  DFFSX4 R9_D_reg_41_ ( .D(n3778), .CK(clk), .SN(rst_n), .QN(BOPD[41]) );
  DFFSX2 R9_B_reg_30_ ( .D(n3728), .CK(clk), .SN(rst_n), .QN(BOPB[30]) );
  DFFSX4 T1_W1_reg_19_ ( .D(n29198), .CK(clk), .SN(rst_n), .Q(n7083), .QN(
        W1[19]) );
  DFFSX2 R9_C_reg_45_ ( .D(n3793), .CK(clk), .SN(rst_n), .QN(BOPC[45]) );
  DFFSX4 R9_B_reg_36_ ( .D(n3752), .CK(clk), .SN(rst_n), .QN(BOPB[36]) );
  DFFSX4 T1_W2_reg_26_ ( .D(n29158), .CK(clk), .SN(rst_n), .QN(W2[26]) );
  DFFSX2 R9_C_reg_36_ ( .D(n3753), .CK(clk), .SN(rst_n), .QN(BOPC[36]) );
  DFFSX2 R7_D_reg_30_ ( .D(n3314), .CK(clk), .SN(rst_n), .QN(AOPD[30]) );
  DFFSX2 R9_C_reg_35_ ( .D(n3749), .CK(clk), .SN(rst_n), .QN(BOPC[35]) );
  DFFSX2 R7_C_reg_30_ ( .D(n3313), .CK(clk), .SN(rst_n), .QN(AOPC[30]) );
  DFFSX2 out_start1_reg ( .D(n29091), .CK(clk), .SN(rst_n), .Q(n28700), .QN(
        n29112) );
  DFFSX4 U0_pipe13_reg_26_ ( .D(n4666), .CK(clk), .SN(rst_n), .Q(n29001), .QN(
        U0_pipe13[26]) );
  DFFSX4 U0_pipe10_reg_27_ ( .D(n4550), .CK(clk), .SN(rst_n), .Q(n28995), .QN(
        U0_pipe10[27]) );
  DFFSX4 U0_pipe3_reg_20_ ( .D(n4355), .CK(clk), .SN(rst_n), .Q(n28777), .QN(
        U0_pipe3[20]) );
  DFFSX4 U1_pipe8_reg_27_ ( .D(n4809), .CK(clk), .SN(rst_n), .Q(n28987), .QN(
        U1_pipe8[27]) );
  DFFSX4 U0_pipe7_reg_27_ ( .D(n4435), .CK(clk), .SN(rst_n), .Q(n28692), .QN(
        U0_pipe7[27]) );
  DFFSX4 U1_pipe15_reg_20_ ( .D(n4799), .CK(clk), .SN(rst_n), .Q(n28873), .QN(
        U1_pipe15[20]) );
  DFFSX4 U1_pipe1_reg_27_ ( .D(n5011), .CK(clk), .SN(rst_n), .Q(n28693), .QN(
        U1_pipe1[27]) );
  DFFSX4 U1_pipe15_reg_26_ ( .D(n4805), .CK(clk), .SN(rst_n), .Q(n29006), .QN(
        U1_pipe15[26]) );
  DFFSX4 U1_pipe9_reg_26_ ( .D(n4836), .CK(clk), .SN(rst_n), .Q(n29003), .QN(
        U1_pipe9[26]) );
  DFFSX4 U0_pipe12_reg_27_ ( .D(n4693), .CK(clk), .SN(rst_n), .Q(n28916), .QN(
        U0_pipe12[27]) );
  DFFSX4 U0_pipe9_reg_26_ ( .D(n4579), .CK(clk), .SN(rst_n), .Q(n28999), .QN(
        U0_pipe9[26]) );
  DFFSX4 U1_pipe13_reg_24_ ( .D(n4747), .CK(clk), .SN(rst_n), .Q(n28948), .QN(
        U1_pipe13[24]) );
  DFFSX4 U0_pipe15_reg_25_ ( .D(n4611), .CK(clk), .SN(rst_n), .Q(n28935), .QN(
        U0_pipe15[25]) );
  DFFSX4 U0_pipe2_reg_27_ ( .D(n4376), .CK(clk), .SN(rst_n), .Q(n28915), .QN(
        U0_pipe2[27]) );
  DFFSX4 U1_pipe13_reg_26_ ( .D(n4749), .CK(clk), .SN(rst_n), .Q(n29005), .QN(
        U1_pipe13[26]) );
  DFFSX4 U0_pipe15_reg_26_ ( .D(n4610), .CK(clk), .SN(rst_n), .Q(n29002), .QN(
        U0_pipe15[26]) );
  DFFSX4 U0_pipe14_reg_27_ ( .D(n4637), .CK(clk), .SN(rst_n), .Q(n28917), .QN(
        U0_pipe14[27]) );
  DFFSX4 U0_pipe11_reg_27_ ( .D(n4522), .CK(clk), .SN(rst_n), .Q(n28691), .QN(
        U0_pipe11[27]) );
  DFFSX4 U1_pipe4_reg_27_ ( .D(n5095), .CK(clk), .SN(rst_n), .Q(n28990), .QN(
        U1_pipe4[27]) );
  DFFSX1 R9_A_reg_0_ ( .D(n3639), .CK(clk), .SN(rst_n), .Q(n28676), .QN(
        BOPA[0]) );
  DFFSX1 T1_W3_reg_8_ ( .D(n29114), .CK(clk), .SN(rst_n), .Q(n8023), .QN(W3[8]) );
  DFFSX4 R9_D_reg_32_ ( .D(n3738), .CK(clk), .SN(rst_n), .QN(BOPD[32]) );
  DFFSX4 R9_B_reg_31_ ( .D(n3732), .CK(clk), .SN(rst_n), .QN(BOPB[31]) );
  DFFSX4 R7_B_reg_33_ ( .D(n3324), .CK(clk), .SN(rst_n), .QN(AOPB[33]) );
  DFFSX4 R7_D_reg_32_ ( .D(n3322), .CK(clk), .SN(rst_n), .QN(AOPD[32]) );
  DFFSX4 R7_B_reg_32_ ( .D(n3320), .CK(clk), .SN(rst_n), .QN(AOPB[32]) );
  DFFSX4 R9_B_reg_27_ ( .D(n3712), .CK(clk), .SN(rst_n), .QN(BOPB[27]) );
  DFFSX4 R9_C_reg_28_ ( .D(n3717), .CK(clk), .SN(rst_n), .QN(BOPC[28]) );
  DFFSX4 R9_C_reg_30_ ( .D(n3729), .CK(clk), .SN(rst_n), .QN(BOPC[30]) );
  DFFSX4 T1_W1_reg_23_ ( .D(n29193), .CK(clk), .SN(rst_n), .QN(W1[23]) );
  DFFSX4 R9_C_reg_29_ ( .D(n3721), .CK(clk), .SN(rst_n), .QN(BOPC[29]) );
  DFFSX4 R7_D_reg_37_ ( .D(n3342), .CK(clk), .SN(rst_n), .QN(AOPD[37]) );
  DFFSX4 T1_W2_reg_23_ ( .D(n29161), .CK(clk), .SN(rst_n), .QN(W2[23]) );
  DFFSX4 T1_W0_reg_23_ ( .D(n29225), .CK(clk), .SN(rst_n), .QN(W0[23]) );
  DFFSX4 R7_B_reg_7_ ( .D(n3416), .CK(clk), .SN(rst_n), .Q(n8066), .QN(AOPB[7]) );
  DFFSX4 T1_W0_reg_25_ ( .D(n29223), .CK(clk), .SN(rst_n), .QN(W0[25]) );
  DFFSX4 R7_B_reg_35_ ( .D(n3332), .CK(clk), .SN(rst_n), .QN(AOPB[35]) );
  DFFSX4 T1_W1_reg_25_ ( .D(n29191), .CK(clk), .SN(rst_n), .QN(W1[25]) );
  DFFSX4 R9_C_reg_5_ ( .D(n3825), .CK(clk), .SN(rst_n), .Q(n8127), .QN(BOPC[5]) );
  DFFSX4 R9_B_reg_29_ ( .D(n3720), .CK(clk), .SN(rst_n), .QN(BOPB[29]) );
  DFFSX4 R9_C_reg_13_ ( .D(n3653), .CK(clk), .SN(rst_n), .Q(n7060), .QN(
        BOPC[13]) );
  DFFSX2 T1_W1_reg_27_ ( .D(n29189), .CK(clk), .SN(rst_n), .QN(W1[27]) );
  DFFSX2 U2_out_valid_reg ( .D(n28697), .CK(clk), .SN(rst_n), .Q(n28922), .QN(
        OP_done1) );
  DFFSX2 U2_valid_reg_1_ ( .D(n28998), .CK(clk), .SN(rst_n), .Q(n28697), .QN(
        U2_valid_1_) );
  DFFSX2 cnt_reg_6_ ( .D(n5673), .CK(clk), .SN(rst_n), .Q(n28704), .QN(cnt[6])
         );
  DFFSX2 R7_valid_reg ( .D(n29242), .CK(clk), .SN(rst_n), .Q(n28985), .QN(
        R7_valid) );
  DFFSX2 R9_C_reg_0_ ( .D(n3637), .CK(clk), .SN(rst_n), .Q(n8194), .QN(BOPC[0]) );
  DFFSX1 R9_D_reg_11_ ( .D(n3646), .CK(clk), .SN(rst_n), .Q(n8189), .QN(
        BOPD[11]) );
  DFFSX4 T1_W1_reg_9_ ( .D(n29177), .CK(clk), .SN(rst_n), .Q(n8050), .QN(W1[9]) );
  DFFSX2 U1_done_reg ( .D(n28997), .CK(clk), .SN(rst_n), .Q(n28921), .QN(
        OP2_done0) );
  DFFSX2 U1_valid_reg_1_ ( .D(n8053), .CK(clk), .SN(rst_n), .Q(n28997), .QN(
        U1_valid[1]) );
  DFFSX2 T1_W3_reg_15_ ( .D(n29138), .CK(clk), .SN(rst_n), .Q(n8000), .QN(
        W3[15]) );
  DFFSX2 cnt_reg_7_ ( .D(n5672), .CK(clk), .SN(rst_n), .Q(n28703), .QN(cnt[7])
         );
  DFFSX2 cnt_reg_0_ ( .D(n5679), .CK(clk), .SN(rst_n), .Q(n28709), .QN(cnt[0])
         );
  DFFSX1 R9_C_reg_19_ ( .D(n3677), .CK(clk), .SN(rst_n), .Q(n7061), .QN(
        BOPC[19]) );
  DFFSX1 R9_C_reg_18_ ( .D(n3673), .CK(clk), .SN(rst_n), .Q(n7059), .QN(
        BOPC[18]) );
  DFFSX1 R9_D_reg_15_ ( .D(n3662), .CK(clk), .SN(rst_n), .Q(n7058), .QN(
        BOPD[15]) );
  DFFSX1 R9_C_reg_16_ ( .D(n3665), .CK(clk), .SN(rst_n), .Q(n7052), .QN(
        BOPC[16]) );
  DFFSX2 R9_B_reg_33_ ( .D(n3740), .CK(clk), .SN(rst_n), .Q(n7045), .QN(
        BOPB[33]) );
  DFFSX2 R9_A_reg_37_ ( .D(n3759), .CK(clk), .SN(rst_n), .Q(n28747), .QN(
        BOPA[37]) );
  DFFSX1 R7_D_reg_18_ ( .D(n3258), .CK(clk), .SN(rst_n), .Q(n6950), .QN(
        AOPD[18]) );
  DFFSX1 R7_B_reg_19_ ( .D(n3260), .CK(clk), .SN(rst_n), .Q(n8108), .QN(
        AOPB[19]) );
  DFFSX1 cs_reg_1_ ( .D(n5683), .CK(clk), .SN(rst_n), .Q(n29111), .QN(cs[1])
         );
  DFFSX1 cs_reg_0_ ( .D(n5681), .CK(clk), .SN(rst_n), .Q(n29110), .QN(cs[0])
         );
  DFFSX2 T1_W3_reg_2_ ( .D(n29122), .CK(clk), .SN(rst_n), .Q(n8036), .QN(W3[2]) );
  DFFSX2 T1_W3_reg_19_ ( .D(n29134), .CK(clk), .SN(rst_n), .QN(W3[19]) );
  DFFSX1 T1_W1_reg_14_ ( .D(n29203), .CK(clk), .SN(rst_n), .Q(n8004), .QN(
        W1[14]) );
  DFFSX1 T1_W2_reg_14_ ( .D(n29171), .CK(clk), .SN(rst_n), .Q(n8012), .QN(
        W2[14]) );
  DFFSX2 T1_W2_reg_12_ ( .D(n29173), .CK(clk), .SN(rst_n), .Q(n7988), .QN(
        W2[12]) );
  DFFSX2 T1_W2_reg_11_ ( .D(n29174), .CK(clk), .SN(rst_n), .Q(n7997), .QN(
        W2[11]) );
  DFFSX2 R9_D_reg_9_ ( .D(n3842), .CK(clk), .SN(rst_n), .Q(n8118), .QN(BOPD[9]) );
  DFFSX2 R9_B_reg_9_ ( .D(n3840), .CK(clk), .SN(rst_n), .Q(n8116), .QN(BOPB[9]) );
  DFFSX2 R9_D_reg_8_ ( .D(n3838), .CK(clk), .SN(rst_n), .Q(n8121), .QN(BOPD[8]) );
  DFFSX2 R9_B_reg_8_ ( .D(n3836), .CK(clk), .SN(rst_n), .Q(n8119), .QN(BOPB[8]) );
  DFFSX2 R9_A_reg_44_ ( .D(n3791), .CK(clk), .SN(rst_n), .Q(n28711), .QN(
        BOPA[44]) );
  DFFSX1 R9_D_reg_43_ ( .D(n3786), .CK(clk), .SN(rst_n), .QN(BOPD[43]) );
  DFFSX1 R9_D_reg_42_ ( .D(n3782), .CK(clk), .SN(rst_n), .QN(BOPD[42]) );
  DFFSX1 R9_C_reg_34_ ( .D(n3745), .CK(clk), .SN(rst_n), .QN(BOPC[34]) );
  DFFSX1 R9_D_reg_21_ ( .D(n3690), .CK(clk), .SN(rst_n), .Q(n8162), .QN(
        BOPD[21]) );
  DFFSX1 R9_C_reg_21_ ( .D(n3689), .CK(clk), .SN(rst_n), .Q(n8161), .QN(
        BOPC[21]) );
  DFFSX1 R9_D_reg_19_ ( .D(n3678), .CK(clk), .SN(rst_n), .Q(n8170), .QN(
        BOPD[19]) );
  DFFSX1 R9_D_reg_18_ ( .D(n3674), .CK(clk), .SN(rst_n), .Q(n8172), .QN(
        BOPD[18]) );
  DFFSX1 R9_C_reg_17_ ( .D(n3669), .CK(clk), .SN(rst_n), .Q(n8176), .QN(
        BOPC[17]) );
  DFFSX1 R9_D_reg_14_ ( .D(n3658), .CK(clk), .SN(rst_n), .QN(BOPD[14]) );
  DFFSX2 R9_B_reg_12_ ( .D(n3648), .CK(clk), .SN(rst_n), .Q(n8184), .QN(
        BOPB[12]) );
  DFFSX2 R9_B_reg_11_ ( .D(n3644), .CK(clk), .SN(rst_n), .Q(n8187), .QN(
        BOPB[11]) );
  DFFSX2 R9_B_reg_10_ ( .D(n3640), .CK(clk), .SN(rst_n), .Q(n8190), .QN(
        BOPB[10]) );
  DFFSX2 R7_D_reg_9_ ( .D(n3426), .CK(clk), .SN(rst_n), .Q(n8060), .QN(AOPD[9]) );
  DFFSX2 R7_D_reg_8_ ( .D(n3422), .CK(clk), .SN(rst_n), .Q(n8063), .QN(AOPD[8]) );
  DFFSX2 R7_B_reg_5_ ( .D(n3408), .CK(clk), .SN(rst_n), .Q(n8072), .QN(AOPB[5]) );
  DFFSX1 R7_D_reg_4_ ( .D(n3398), .CK(clk), .SN(rst_n), .Q(n8075), .QN(AOPD[4]) );
  DFFSX1 R7_C_reg_43_ ( .D(n3369), .CK(clk), .SN(rst_n), .QN(AOPC[43]) );
  DFFSX1 R7_B_reg_43_ ( .D(n3368), .CK(clk), .SN(rst_n), .QN(AOPB[43]) );
  DFFSX1 R7_C_reg_42_ ( .D(n3365), .CK(clk), .SN(rst_n), .QN(AOPC[42]) );
  DFFSX1 R7_C_reg_41_ ( .D(n3361), .CK(clk), .SN(rst_n), .QN(AOPC[41]) );
  DFFSX1 R7_C_reg_40_ ( .D(n3357), .CK(clk), .SN(rst_n), .QN(AOPC[40]) );
  DFFSX2 R7_C_reg_3_ ( .D(n3353), .CK(clk), .SN(rst_n), .Q(n8079), .QN(AOPC[3]) );
  DFFSX2 R7_B_reg_3_ ( .D(n3352), .CK(clk), .SN(rst_n), .Q(n8081), .QN(AOPB[3]) );
  DFFSX1 R7_B_reg_36_ ( .D(n3336), .CK(clk), .SN(rst_n), .QN(AOPB[36]) );
  DFFSX1 R7_D_reg_21_ ( .D(n3274), .CK(clk), .SN(rst_n), .Q(n8097), .QN(
        AOPD[21]) );
  DFFSX1 R7_C_reg_21_ ( .D(n3273), .CK(clk), .SN(rst_n), .Q(n8096), .QN(
        AOPC[21]) );
  DFFSX1 R7_B_reg_21_ ( .D(n3272), .CK(clk), .SN(rst_n), .Q(n8098), .QN(
        AOPB[21]) );
  DFFSX1 R7_C_reg_19_ ( .D(n3261), .CK(clk), .SN(rst_n), .Q(n8106), .QN(
        AOPC[19]) );
  DFFSX1 R7_C_reg_18_ ( .D(n3257), .CK(clk), .SN(rst_n), .Q(n8109), .QN(
        AOPC[18]) );
  DFFSX1 R7_B_reg_18_ ( .D(n3256), .CK(clk), .SN(rst_n), .Q(n8110), .QN(
        AOPB[18]) );
  DFFSX1 R7_C_reg_17_ ( .D(n3253), .CK(clk), .SN(rst_n), .Q(n8111), .QN(
        AOPC[17]) );
  DFFSX1 R7_C_reg_16_ ( .D(n3249), .CK(clk), .SN(rst_n), .Q(n8114), .QN(
        AOPC[16]) );
  DFFSX1 R7_D_reg_15_ ( .D(n3246), .CK(clk), .SN(rst_n), .Q(n8196), .QN(
        AOPD[15]) );
  DFFSX1 R7_C_reg_15_ ( .D(n3245), .CK(clk), .SN(rst_n), .Q(n8195), .QN(
        AOPC[15]) );
  DFFSX1 R7_C_reg_14_ ( .D(n3241), .CK(clk), .SN(rst_n), .Q(n7992), .QN(
        AOPC[14]) );
  DFFSX2 R7_D_reg_13_ ( .D(n3238), .CK(clk), .SN(rst_n), .Q(n7989), .QN(
        AOPD[13]) );
  DFFSX2 R7_C_reg_13_ ( .D(n3237), .CK(clk), .SN(rst_n), .Q(n7954), .QN(
        AOPC[13]) );
  DFFSX2 R7_B_reg_13_ ( .D(n3236), .CK(clk), .SN(rst_n), .Q(n8198), .QN(
        AOPB[13]) );
  DFFSX1 R7_D_reg_12_ ( .D(n3234), .CK(clk), .SN(rst_n), .Q(n8199), .QN(
        AOPD[12]) );
  DFFSX2 R7_B_reg_12_ ( .D(n3232), .CK(clk), .SN(rst_n), .Q(n7955), .QN(
        AOPB[12]) );
  DFFSX2 R7_D_reg_11_ ( .D(n3230), .CK(clk), .SN(rst_n), .Q(n8201), .QN(
        AOPD[11]) );
  DFFSX2 R7_C_reg_11_ ( .D(n3229), .CK(clk), .SN(rst_n), .Q(n8200), .QN(
        AOPC[11]) );
  DFFSX2 R7_B_reg_11_ ( .D(n3228), .CK(clk), .SN(rst_n), .Q(n8202), .QN(
        AOPB[11]) );
  DFFSX2 R7_C_reg_10_ ( .D(n3225), .CK(clk), .SN(rst_n), .Q(n8203), .QN(
        AOPC[10]) );
  DFFSX2 R7_B_reg_10_ ( .D(n3224), .CK(clk), .SN(rst_n), .Q(n8205), .QN(
        AOPB[10]) );
  DFFSX2 R7_C_reg_0_ ( .D(n3221), .CK(clk), .SN(rst_n), .Q(n8206), .QN(AOPC[0]) );
  DFFSX1 R9_A_reg_46_ ( .D(n3799), .CK(clk), .SN(rst_n), .Q(n28708), .QN(
        BOPA[46]) );
  DFFSX1 R9_A_reg_45_ ( .D(n3795), .CK(clk), .SN(rst_n), .Q(n28686), .QN(
        BOPA[45]) );
  DFFSX1 R9_A_reg_47_ ( .D(n3803), .CK(clk), .SN(rst_n), .Q(n28685), .QN(
        BOPA[47]) );
  DFFSX1 cs_reg_2_ ( .D(n5682), .CK(clk), .SN(rst_n), .Q(n28912), .QN(cs[2])
         );
  DFFSX2 R7_C_reg_38_ ( .D(n3345), .CK(clk), .SN(rst_n), .QN(AOPC[38]) );
  DFFSX2 T1_W2_reg_27_ ( .D(n29157), .CK(clk), .SN(rst_n), .QN(W2[27]) );
  DFFSX2 R9_C_reg_38_ ( .D(n3761), .CK(clk), .SN(rst_n), .QN(BOPC[38]) );
  DFFSX1 cnt_reg_8_ ( .D(n5671), .CK(clk), .SN(rst_n), .Q(n28706), .QN(cnt[8])
         );
  DFFSX2 R9_C_reg_33_ ( .D(n3741), .CK(clk), .SN(rst_n), .QN(BOPC[33]) );
  DFFSX1 U1_pipe4_reg_23_ ( .D(n5091), .CK(clk), .SN(rst_n), .QN(U1_pipe4[23])
         );
  DFFSX1 U1_pipe6_reg_22_ ( .D(n4947), .CK(clk), .SN(rst_n), .QN(U1_pipe6[22])
         );
  DFFSX1 U1_pipe3_reg_17_ ( .D(n5057), .CK(clk), .SN(rst_n), .Q(n28844), .QN(
        U1_pipe3[17]) );
  DFFSX1 U1_pipe3_reg_19_ ( .D(n5059), .CK(clk), .SN(rst_n), .Q(n28842), .QN(
        U1_pipe3[19]) );
  DFFSX1 U0_pipe3_reg_17_ ( .D(n4358), .CK(clk), .SN(rst_n), .Q(n28780), .QN(
        U0_pipe3[17]) );
  DFFSX1 U1_pipe3_reg_16_ ( .D(n5056), .CK(clk), .SN(rst_n), .Q(n28845), .QN(
        U1_pipe3[16]) );
  DFFSX1 U0_pipe15_reg_22_ ( .D(n4614), .CK(clk), .SN(rst_n), .Q(n28938), .QN(
        U0_pipe15[22]) );
  DFFSX1 U1_pipe2_reg_27_ ( .D(n5039), .CK(clk), .SN(rst_n), .Q(n28913), .QN(
        U1_pipe2[27]) );
  DFFSX1 U0_pipe3_reg_24_ ( .D(n4351), .CK(clk), .SN(rst_n), .Q(n28928), .QN(
        U0_pipe3[24]) );
  DFFSX1 U0_pipe15_reg_23_ ( .D(n4613), .CK(clk), .SN(rst_n), .Q(n28937), .QN(
        U0_pipe15[23]) );
  DFFSX1 U0_pipe3_reg_18_ ( .D(n4357), .CK(clk), .SN(rst_n), .Q(n28779), .QN(
        U0_pipe3[18]) );
  DFFSX1 U0_pipe3_reg_23_ ( .D(n4352), .CK(clk), .SN(rst_n), .Q(n28929), .QN(
        U0_pipe3[23]) );
  DFFSX1 U1_pipe3_reg_18_ ( .D(n5058), .CK(clk), .SN(rst_n), .Q(n28843), .QN(
        U1_pipe3[18]) );
  DFFSX1 U1_pipe9_reg_20_ ( .D(n4830), .CK(clk), .SN(rst_n), .Q(n28825), .QN(
        U1_pipe9[20]) );
  DFFSX1 U0_pipe3_reg_22_ ( .D(n4353), .CK(clk), .SN(rst_n), .Q(n28930), .QN(
        U0_pipe3[22]) );
  DFFSX1 U0_pipe13_reg_22_ ( .D(n4670), .CK(clk), .SN(rst_n), .Q(n28934), .QN(
        U0_pipe13[22]) );
  DFFSX1 U0_pipe13_reg_23_ ( .D(n4669), .CK(clk), .SN(rst_n), .Q(n28933), .QN(
        U0_pipe13[23]) );
  DFFSX1 U0_pipe13_reg_24_ ( .D(n4668), .CK(clk), .SN(rst_n), .Q(n28932), .QN(
        U0_pipe13[24]) );
  DFFSX1 U1_pipe6_reg_27_ ( .D(n4952), .CK(clk), .SN(rst_n), .Q(n28992), .QN(
        U1_pipe6[27]) );
  DFFSX1 U1_pipe3_reg_20_ ( .D(n5060), .CK(clk), .SN(rst_n), .Q(n28841), .QN(
        U1_pipe3[20]) );
  DFFSX1 U0_pipe5_reg_27_ ( .D(n4491), .CK(clk), .SN(rst_n), .Q(n28690), .QN(
        U0_pipe5[27]) );
  DFFSX1 U1_pipe12_reg_27_ ( .D(n4722), .CK(clk), .SN(rst_n), .Q(n28918), .QN(
        U1_pipe12[27]) );
  DFFSX1 U0_pipe0_reg_27_ ( .D(n4285), .CK(clk), .SN(rst_n), .Q(n28993), .QN(
        U0_pipe0[27]) );
  DFFSX1 U1_pipe0_reg_27_ ( .D(n5130), .CK(clk), .SN(rst_n), .Q(n28989), .QN(
        U1_pipe0[27]) );
  DFFSX2 R7_B_reg_30_ ( .D(n3312), .CK(clk), .SN(rst_n), .QN(AOPB[30]) );
  DFFSX2 R7_B_reg_27_ ( .D(n3296), .CK(clk), .SN(rst_n), .QN(AOPB[27]) );
  DFFSX2 R9_C_reg_31_ ( .D(n3733), .CK(clk), .SN(rst_n), .QN(BOPC[31]) );
  DFFSX2 R9_C_reg_43_ ( .D(n3785), .CK(clk), .SN(rst_n), .QN(BOPC[43]) );
  DFFSX2 R9_B_reg_4_ ( .D(n3812), .CK(clk), .SN(rst_n), .Q(n8132), .QN(BOPB[4]) );
  DFFSHQX4 T1_W0_reg_2_ ( .D(n29218), .CK(clk), .SN(rst_n), .Q(n6875) );
  DFFSX2 T1_W3_reg_23_ ( .D(n29129), .CK(clk), .SN(rst_n), .QN(W3[23]) );
  DFFSX4 T1_W1_reg_11_ ( .D(n29206), .CK(clk), .SN(rst_n), .Q(n8024), .QN(
        W1[11]) );
  DFFSX4 R7_C_reg_34_ ( .D(n3329), .CK(clk), .SN(rst_n), .QN(AOPC[34]) );
  DFFSX4 R9_D_reg_29_ ( .D(n3722), .CK(clk), .SN(rst_n), .QN(BOPD[29]) );
  DFFSX2 R9_C_reg_41_ ( .D(n3777), .CK(clk), .SN(rst_n), .QN(BOPC[41]) );
  DFFSX1 R7_D_reg_5_ ( .D(n3410), .CK(clk), .SN(rst_n), .Q(n8071), .QN(AOPD[5]) );
  DFFSX2 T1_W3_reg_0_ ( .D(n29144), .CK(clk), .SN(rst_n), .Q(n8019), .QN(W3[0]) );
  DFFSX2 R9_B_reg_5_ ( .D(n3824), .CK(clk), .SN(rst_n), .Q(n8126), .QN(BOPB[5]) );
  DFFSX2 R9_C_reg_4_ ( .D(n3813), .CK(clk), .SN(rst_n), .Q(n8133), .QN(BOPC[4]) );
  DFFSX1 R9_D_reg_38_ ( .D(n3762), .CK(clk), .SN(rst_n), .QN(BOPD[38]) );
  DFFSX1 R9_B_reg_21_ ( .D(n3688), .CK(clk), .SN(rst_n), .Q(n8160), .QN(
        BOPB[21]) );
  DFFSX2 R9_B_reg_0_ ( .D(n3636), .CK(clk), .SN(rst_n), .Q(n8193), .QN(BOPB[0]) );
  DFFSX2 R7_B_reg_9_ ( .D(n3424), .CK(clk), .SN(rst_n), .Q(n8061), .QN(AOPB[9]) );
  DFFSX1 R7_D_reg_45_ ( .D(n3378), .CK(clk), .SN(rst_n), .QN(AOPD[45]) );
  DFFSX1 R7_C_reg_32_ ( .D(n3321), .CK(clk), .SN(rst_n), .QN(AOPC[32]) );
  DFFSX2 R9_D_reg_45_ ( .D(n3794), .CK(clk), .SN(rst_n), .QN(BOPD[45]) );
  DFFSX1 U1_pipe7_reg_27_ ( .D(n4980), .CK(clk), .SN(rst_n), .Q(n28696), .QN(
        U1_pipe7[27]) );
  DFFSX2 R9_B_reg_32_ ( .D(n3736), .CK(clk), .SN(rst_n), .QN(BOPB[32]) );
  DFFSX1 cnt_reg_4_ ( .D(n5675), .CK(clk), .SN(rst_n), .Q(n28680), .QN(cnt[4])
         );
  DFFSX1 R9_D_reg_40_ ( .D(n3774), .CK(clk), .SN(rst_n), .Q(n7053), .QN(
        BOPD[40]) );
  DFFSX1 R9_D_reg_16_ ( .D(n3666), .CK(clk), .SN(rst_n), .Q(n8178), .QN(
        BOPD[16]) );
  DFFSX1 R7_B_reg_17_ ( .D(n3252), .CK(clk), .SN(rst_n), .Q(n8113), .QN(
        AOPB[17]) );
  DFFSX1 T1_W3_reg_25_ ( .D(n29127), .CK(clk), .SN(rst_n), .QN(W3[25]) );
  DFFSX2 R9_A_reg_35_ ( .D(n3751), .CK(clk), .SN(rst_n), .Q(n6932), .QN(
        BOPA[35]) );
  DFFSX2 T1_W1_reg_24_ ( .D(n29192), .CK(clk), .SN(rst_n), .QN(W1[24]) );
  DFFSX2 R9_A_reg_39_ ( .D(n3767), .CK(clk), .SN(rst_n), .Q(n28681), .QN(
        BOPA[39]) );
  DFFSX2 R9_C_reg_27_ ( .D(n3713), .CK(clk), .SN(rst_n), .QN(BOPC[27]) );
  DFFSX2 R9_C_reg_3_ ( .D(n3769), .CK(clk), .SN(rst_n), .Q(n8136), .QN(BOPC[3]) );
  DFFSX1 R9_A_reg_43_ ( .D(n3787), .CK(clk), .SN(rst_n), .Q(n28688), .QN(
        BOPA[43]) );
  DFFSX1 R9_A_reg_42_ ( .D(n3783), .CK(clk), .SN(rst_n), .Q(n28712), .QN(
        BOPA[42]) );
  DFFSX2 R9_C_reg_44_ ( .D(n3789), .CK(clk), .SN(rst_n), .QN(BOPC[44]) );
  DFFSX2 R7_D_reg_1_ ( .D(n3266), .CK(clk), .SN(rst_n), .Q(n8103), .QN(AOPD[1]) );
  DFFSX2 R9_B_reg_1_ ( .D(n3680), .CK(clk), .SN(rst_n), .Q(n8166), .QN(BOPB[1]) );
  DFFSX1 R7_D_reg_34_ ( .D(n3330), .CK(clk), .SN(rst_n), .QN(AOPD[34]) );
  DFFSX2 R9_C_reg_10_ ( .D(n3641), .CK(clk), .SN(rst_n), .Q(n8191), .QN(
        BOPC[10]) );
  DFFSX2 R9_C_reg_39_ ( .D(n3765), .CK(clk), .SN(rst_n), .QN(BOPC[39]) );
  DFFSX2 R9_C_reg_11_ ( .D(n3645), .CK(clk), .SN(rst_n), .Q(n8188), .QN(
        BOPC[11]) );
  DFFSX2 R9_B_reg_13_ ( .D(n3652), .CK(clk), .SN(rst_n), .Q(n8183), .QN(
        BOPB[13]) );
  DFFSX2 R9_C_reg_37_ ( .D(n3757), .CK(clk), .SN(rst_n), .QN(BOPC[37]) );
  DFFSX2 R7_C_reg_1_ ( .D(n3265), .CK(clk), .SN(rst_n), .Q(n8102), .QN(AOPC[1]) );
  DFFSX2 T1_W3_reg_17_ ( .D(n29136), .CK(clk), .SN(rst_n), .QN(W3[17]) );
  DFFSX2 T1_W1_reg_10_ ( .D(n29207), .CK(clk), .SN(rst_n), .Q(n7952), .QN(
        W1[10]) );
  DFFSX1 R9_D_reg_31_ ( .D(n3734), .CK(clk), .SN(rst_n), .QN(BOPD[31]) );
  DFFSX1 R9_D_reg_30_ ( .D(n3730), .CK(clk), .SN(rst_n), .QN(BOPD[30]) );
  DFFSX1 R9_D_reg_6_ ( .D(n3830), .CK(clk), .SN(rst_n), .Q(n8125), .QN(BOPD[6]) );
  DFFSX1 R9_D_reg_5_ ( .D(n3826), .CK(clk), .SN(rst_n), .Q(n8128), .QN(BOPD[5]) );
  DFFSX1 R9_D_reg_17_ ( .D(n3670), .CK(clk), .SN(rst_n), .Q(n8177), .QN(
        BOPD[17]) );
  DFFSX1 R9_C_reg_15_ ( .D(n3661), .CK(clk), .SN(rst_n), .Q(n8180), .QN(
        BOPC[15]) );
  DFFSX1 R9_C_reg_32_ ( .D(n3737), .CK(clk), .SN(rst_n), .QN(BOPC[32]) );
  DFFSX1 R7_B_reg_42_ ( .D(n3364), .CK(clk), .SN(rst_n), .QN(AOPB[42]) );
  DFFSX1 R9_C_reg_8_ ( .D(n3837), .CK(clk), .SN(rst_n), .Q(n8120), .QN(BOPC[8]) );
  DFFSX1 R9_C_reg_40_ ( .D(n3773), .CK(clk), .SN(rst_n), .QN(BOPC[40]) );
  DFFSX1 R7_B_reg_16_ ( .D(n3248), .CK(clk), .SN(rst_n), .Q(n7057), .QN(
        AOPB[16]) );
  DFFSX1 R9_D_reg_7_ ( .D(n3834), .CK(clk), .SN(rst_n), .Q(n8122), .QN(BOPD[7]) );
  DFFSX1 R9_C_reg_14_ ( .D(n3657), .CK(clk), .SN(rst_n), .Q(n8181), .QN(
        BOPC[14]) );
  DFFSX1 T1_W0_reg_14_ ( .D(n29235), .CK(clk), .SN(rst_n), .Q(n7975), .QN(
        W0[14]) );
  DFFSX1 R7_D_reg_7_ ( .D(n3418), .CK(clk), .SN(rst_n), .Q(n8065), .QN(AOPD[7]) );
  DFFSX2 R7_B_reg_26_ ( .D(n3292), .CK(clk), .SN(rst_n), .QN(AOPB[26]) );
  DFFSX2 R7_B_reg_2_ ( .D(n3308), .CK(clk), .SN(rst_n), .Q(n8085), .QN(AOPB[2]) );
  DFFSX2 R7_C_reg_6_ ( .D(n3413), .CK(clk), .SN(rst_n), .Q(n8067), .QN(AOPC[6]) );
  DFFSX2 R7_D_reg_33_ ( .D(n3326), .CK(clk), .SN(rst_n), .QN(AOPD[33]) );
  DFFSX2 T1_W1_reg_12_ ( .D(n29205), .CK(clk), .SN(rst_n), .Q(n7972), .QN(
        W1[12]) );
  DFFSX1 R7_D_reg_31_ ( .D(n3318), .CK(clk), .SN(rst_n), .QN(AOPD[31]) );
  DFFSX1 R7_D_reg_40_ ( .D(n3358), .CK(clk), .SN(rst_n), .QN(AOPD[40]) );
  DFFSX1 R7_D_reg_14_ ( .D(n3242), .CK(clk), .SN(rst_n), .Q(n7054), .QN(
        AOPD[14]) );
  DFFSX1 R7_C_reg_33_ ( .D(n3325), .CK(clk), .SN(rst_n), .QN(AOPC[33]) );
  DFFSX1 R7_D_reg_6_ ( .D(n3414), .CK(clk), .SN(rst_n), .Q(n8068), .QN(AOPD[6]) );
  DFFSX1 R7_D_reg_16_ ( .D(n3250), .CK(clk), .SN(rst_n), .Q(n8115), .QN(
        AOPD[16]) );
  DFFSX2 R9_D_reg_13_ ( .D(n3654), .CK(clk), .SN(rst_n), .Q(n8182), .QN(
        BOPD[13]) );
  DFFSX2 R7_D_reg_44_ ( .D(n3374), .CK(clk), .SN(rst_n), .QN(AOPD[44]) );
  DFFSX1 R7_D_reg_42_ ( .D(n3366), .CK(clk), .SN(rst_n), .QN(AOPD[42]) );
  DFFSX1 R7_B_reg_41_ ( .D(n3360), .CK(clk), .SN(rst_n), .QN(AOPB[41]) );
  DFFSX1 R7_D_reg_19_ ( .D(n3262), .CK(clk), .SN(rst_n), .Q(n8107), .QN(
        AOPD[19]) );
  DFFSX1 R9_D_reg_12_ ( .D(n3650), .CK(clk), .SN(rst_n), .Q(n8186), .QN(
        BOPD[12]) );
  DFFSX1 R9_D_reg_10_ ( .D(n3642), .CK(clk), .SN(rst_n), .Q(n8192), .QN(
        BOPD[10]) );
  DFFSX1 R7_B_reg_15_ ( .D(n3244), .CK(clk), .SN(rst_n), .Q(n8197), .QN(
        AOPB[15]) );
  DFFSX1 R9_D_reg_37_ ( .D(n3758), .CK(clk), .SN(rst_n), .QN(BOPD[37]) );
  DFFSX1 R9_D_reg_35_ ( .D(n3750), .CK(clk), .SN(rst_n), .QN(BOPD[35]) );
  DFFSX1 R7_D_reg_43_ ( .D(n3370), .CK(clk), .SN(rst_n), .QN(AOPD[43]) );
  DFFSX1 R7_D_reg_17_ ( .D(n3254), .CK(clk), .SN(rst_n), .Q(n8112), .QN(
        AOPD[17]) );
  DFFSX1 R9_B_reg_19_ ( .D(n3676), .CK(clk), .SN(rst_n), .Q(n8169), .QN(
        BOPB[19]) );
  DFFSX2 R9_B_reg_17_ ( .D(n3668), .CK(clk), .SN(rst_n), .Q(n8175), .QN(
        BOPB[17]) );
  DFFSX2 R9_B_reg_45_ ( .D(n3792), .CK(clk), .SN(rst_n), .QN(BOPB[45]) );
  DFFSX2 R7_C_reg_35_ ( .D(n3333), .CK(clk), .SN(rst_n), .QN(AOPC[35]) );
  DFFSX2 R7_C_reg_9_ ( .D(n3425), .CK(clk), .SN(rst_n), .Q(n8059), .QN(AOPC[9]) );
  DFFSX1 R9_B_reg_42_ ( .D(n3780), .CK(clk), .SN(rst_n), .QN(BOPB[42]) );
  DFFSX1 R9_B_reg_16_ ( .D(n3664), .CK(clk), .SN(rst_n), .Q(n7055), .QN(
        BOPB[16]) );
  DFFSX1 R9_B_reg_18_ ( .D(n3672), .CK(clk), .SN(rst_n), .Q(n8171), .QN(
        BOPB[18]) );
  DFFSX1 T1_W3_reg_13_ ( .D(n29140), .CK(clk), .SN(rst_n), .Q(n8016), .QN(
        W3[13]) );
  DFFSX1 U0_pipe3_reg_16_ ( .D(n4359), .CK(clk), .SN(rst_n), .Q(n28781), .QN(
        U0_pipe3[16]) );
  DFFSX1 U0_pipe13_reg_18_ ( .D(n4674), .CK(clk), .SN(rst_n), .Q(n28795), .QN(
        U0_pipe13[18]) );
  DFFSX1 U0_pipe15_reg_20_ ( .D(n4616), .CK(clk), .SN(rst_n), .Q(n28809), .QN(
        U0_pipe15[20]) );
  DFFSX1 U0_pipe13_reg_20_ ( .D(n4672), .CK(clk), .SN(rst_n), .Q(n28793), .QN(
        U0_pipe13[20]) );
  DFFSX1 U1_pipe13_reg_22_ ( .D(n4745), .CK(clk), .SN(rst_n), .Q(n28950), .QN(
        U1_pipe13[22]) );
  DFFSX1 U1_pipe3_reg_22_ ( .D(n5062), .CK(clk), .SN(rst_n), .Q(n28946), .QN(
        U1_pipe3[22]) );
  DFFSX1 U1_pipe13_reg_23_ ( .D(n4746), .CK(clk), .SN(rst_n), .Q(n28949), .QN(
        U1_pipe13[23]) );
  DFFSX1 U1_pipe3_reg_23_ ( .D(n5063), .CK(clk), .SN(rst_n), .Q(n28945), .QN(
        U1_pipe3[23]) );
  DFFSX1 U1_pipe3_reg_24_ ( .D(n5064), .CK(clk), .SN(rst_n), .Q(n28944), .QN(
        U1_pipe3[24]) );
  DFFSX1 U1_pipe9_reg_25_ ( .D(n4835), .CK(clk), .SN(rst_n), .Q(n28939), .QN(
        U1_pipe9[25]) );
  DFFSX1 U0_pipe3_reg_25_ ( .D(n4350), .CK(clk), .SN(rst_n), .Q(n28927), .QN(
        U0_pipe3[25]) );
  DFFSX1 U1_pipe15_reg_25_ ( .D(n4804), .CK(clk), .SN(rst_n), .Q(n28951), .QN(
        U1_pipe15[25]) );
  DFFSX1 U1_pipe0_reg_25_ ( .D(n5128), .CK(clk), .SN(rst_n), .QN(U1_pipe0[25])
         );
  DFFSX1 U1_pipe3_reg_26_ ( .D(n5066), .CK(clk), .SN(rst_n), .Q(n29004), .QN(
        U1_pipe3[26]) );
  DFFSX1 U0_pipe1_reg_27_ ( .D(n4404), .CK(clk), .SN(rst_n), .Q(n28689), .QN(
        U0_pipe1[27]) );
  DFFSX1 U1_pipe14_reg_27_ ( .D(n4778), .CK(clk), .SN(rst_n), .Q(n28988), .QN(
        U1_pipe14[27]) );
  DFFSX1 U0_pipe8_reg_27_ ( .D(n4606), .CK(clk), .SN(rst_n), .Q(n28914), .QN(
        U0_pipe8[27]) );
  DFFSX1 U1_pipe10_reg_27_ ( .D(n4865), .CK(clk), .SN(rst_n), .Q(n28991), .QN(
        U1_pipe10[27]) );
  DFFSX1 U0_pipe4_reg_27_ ( .D(n4320), .CK(clk), .SN(rst_n), .Q(n28994), .QN(
        U0_pipe4[27]) );
  DFFSX2 U2_valid_reg_0_ ( .D(n28702), .CK(clk), .SN(rst_n), .Q(n28998), .QN(
        n8054) );
  OAI21XL U6295 ( .A0(n21811), .A1(n6728), .B0(n6727), .Y(n4464) );
  BUFX4 U6296 ( .A(n25330), .Y(n6887) );
  XOR2X1 U6297 ( .A(n22461), .B(n7555), .Y(n22462) );
  XOR2X1 U6298 ( .A(n7446), .B(n19574), .Y(n7268) );
  XOR2X1 U6299 ( .A(n12339), .B(n7715), .Y(n9606) );
  XOR2X2 U6300 ( .A(n6805), .B(n7731), .Y(n21947) );
  AOI211XL U6301 ( .A0(n28252), .A1(n27659), .B0(n28459), .C0(n27444), .Y(
        n27445) );
  AOI211XL U6302 ( .A0(n28252), .A1(n27513), .B0(n28299), .C0(n27395), .Y(
        n27396) );
  AOI211XL U6303 ( .A0(n28252), .A1(n27525), .B0(n28313), .C0(n27399), .Y(
        n27400) );
  AOI211XL U6304 ( .A0(n28252), .A1(n27580), .B0(n28378), .C0(n27417), .Y(
        n27418) );
  AOI211XL U6305 ( .A0(n28252), .A1(n27696), .B0(n28501), .C0(n27456), .Y(
        n27457) );
  AOI211XL U6306 ( .A0(n28252), .A1(n27714), .B0(n28522), .C0(n27462), .Y(
        n27463) );
  AOI211XL U6307 ( .A0(n28252), .A1(n27507), .B0(n28291), .C0(n27393), .Y(
        n27394) );
  AOI211XL U6308 ( .A0(n28252), .A1(n27531), .B0(n28320), .C0(n27401), .Y(
        n27402) );
  AOI211XL U6309 ( .A0(n28252), .A1(n27574), .B0(n28371), .C0(n27415), .Y(
        n27416) );
  AOI211XL U6310 ( .A0(n28252), .A1(n27586), .B0(n28385), .C0(n27419), .Y(
        n27420) );
  AOI211XL U6311 ( .A0(n28252), .A1(n27665), .B0(n28466), .C0(n27446), .Y(
        n27447) );
  AOI211XL U6312 ( .A0(n28252), .A1(n27702), .B0(n28508), .C0(n27458), .Y(
        n27459) );
  AOI211XL U6313 ( .A0(n28322), .A1(n28321), .B0(n28320), .C0(n28319), .Y(
        n28323) );
  AOI211XL U6314 ( .A0(n5826), .A1(n28379), .B0(n28378), .C0(n27872), .Y(
        n27873) );
  AOI211XL U6315 ( .A0(n5826), .A1(n27696), .B0(n28501), .C0(n27202), .Y(
        n27203) );
  AOI211XL U6316 ( .A0(n5826), .A1(n27531), .B0(n28320), .C0(n27104), .Y(
        n27105) );
  AOI211XL U6317 ( .A0(n5826), .A1(n28460), .B0(n28459), .C0(n27936), .Y(
        n27937) );
  AOI211XL U6318 ( .A0(n5826), .A1(n27659), .B0(n28459), .C0(n27184), .Y(
        n27185) );
  AOI211XL U6319 ( .A0(n5826), .A1(n27525), .B0(n28313), .C0(n27101), .Y(
        n27102) );
  XOR2X2 U6320 ( .A(n6122), .B(n7902), .Y(n6121) );
  AOI211XL U6321 ( .A0(n27162), .A1(n27513), .B0(n28299), .C0(n27095), .Y(
        n27096) );
  AOI211XL U6322 ( .A0(n27162), .A1(n27580), .B0(n28378), .C0(n27132), .Y(
        n27133) );
  AOI211XL U6323 ( .A0(n27162), .A1(n27714), .B0(n28522), .C0(n27214), .Y(
        n27215) );
  AOI211XL U6324 ( .A0(n27162), .A1(n27507), .B0(n28291), .C0(n27092), .Y(
        n27093) );
  AOI211XL U6325 ( .A0(n27162), .A1(n28386), .B0(n28385), .C0(n27877), .Y(
        n27878) );
  AOI211XL U6326 ( .A0(n27162), .A1(n28467), .B0(n28466), .C0(n27940), .Y(
        n27941) );
  AOI211XL U6327 ( .A0(n27162), .A1(n27665), .B0(n28466), .C0(n27187), .Y(
        n27188) );
  AOI211XL U6328 ( .A0(n27162), .A1(n27793), .B0(n28625), .C0(n27267), .Y(
        n27268) );
  AOI211XL U6329 ( .A0(n27162), .A1(n28292), .B0(n28291), .C0(n27821), .Y(
        n27822) );
  AOI211XL U6330 ( .A0(n27162), .A1(n28372), .B0(n28371), .C0(n27867), .Y(
        n27868) );
  AOI211XL U6331 ( .A0(n27162), .A1(n27574), .B0(n28371), .C0(n27128), .Y(
        n27129) );
  AOI211XL U6332 ( .A0(n27162), .A1(n27586), .B0(n28385), .C0(n27136), .Y(
        n27137) );
  AOI211XL U6333 ( .A0(n27162), .A1(n27702), .B0(n28508), .C0(n27206), .Y(
        n27207) );
  AOI211XL U6334 ( .A0(n27631), .A1(n27659), .B0(n28459), .C0(n27658), .Y(
        n27660) );
  AOI211XL U6335 ( .A0(n27631), .A1(n28300), .B0(n28299), .C0(n28298), .Y(
        n28301) );
  AOI211XL U6336 ( .A0(n27631), .A1(n28314), .B0(n28313), .C0(n28312), .Y(
        n28315) );
  AOI211XL U6337 ( .A0(n27631), .A1(n28502), .B0(n28501), .C0(n28500), .Y(
        n28503) );
  AOI211XL U6338 ( .A0(n27631), .A1(n28523), .B0(n28522), .C0(n28521), .Y(
        n28524) );
  AOI211XL U6339 ( .A0(n27631), .A1(n27531), .B0(n28320), .C0(n27530), .Y(
        n27532) );
  AOI211XL U6340 ( .A0(n27631), .A1(n27586), .B0(n28385), .C0(n27585), .Y(
        n27587) );
  AOI211XL U6341 ( .A0(n27631), .A1(n27702), .B0(n28508), .C0(n27701), .Y(
        n27703) );
  AOI211XL U6342 ( .A0(n27631), .A1(n28509), .B0(n28508), .C0(n28507), .Y(
        n28510) );
  AOI211XL U6343 ( .A0(n27631), .A1(n27525), .B0(n28313), .C0(n27524), .Y(
        n27526) );
  AOI211XL U6344 ( .A0(n27631), .A1(n27580), .B0(n28378), .C0(n27579), .Y(
        n27581) );
  AOI211XL U6345 ( .A0(n27631), .A1(n27714), .B0(n28522), .C0(n27713), .Y(
        n27715) );
  AOI211XL U6346 ( .A0(n27631), .A1(n27665), .B0(n28466), .C0(n27664), .Y(
        n27666) );
  AOI211XL U6347 ( .A0(n27631), .A1(n27793), .B0(n28625), .C0(n27792), .Y(
        n27794) );
  AOI211XL U6348 ( .A0(n5921), .A1(n27586), .B0(n28385), .C0(n27311), .Y(
        n27312) );
  AOI211XL U6349 ( .A0(n5921), .A1(n27580), .B0(n28378), .C0(n27309), .Y(
        n27310) );
  AOI211XL U6350 ( .A0(n5921), .A1(n27574), .B0(n28371), .C0(n27307), .Y(
        n27308) );
  AOI211XL U6351 ( .A0(n5827), .A1(n27513), .B0(n28299), .C0(n27512), .Y(
        n27514) );
  AOI211XL U6352 ( .A0(n5798), .A1(n27507), .B0(n28291), .C0(n27506), .Y(
        n27508) );
  AOI211XL U6353 ( .A0(n5798), .A1(n27574), .B0(n28371), .C0(n27573), .Y(
        n27575) );
  AOI211XL U6354 ( .A0(n28143), .A1(n27659), .B0(n28459), .C0(n27335), .Y(
        n27336) );
  AOI211XL U6355 ( .A0(n28143), .A1(n27513), .B0(n28299), .C0(n27286), .Y(
        n27287) );
  AOI211XL U6356 ( .A0(n28143), .A1(n27525), .B0(n28313), .C0(n27290), .Y(
        n27291) );
  AOI211XL U6357 ( .A0(n28143), .A1(n27696), .B0(n28501), .C0(n27347), .Y(
        n27348) );
  AOI211XL U6358 ( .A0(n28143), .A1(n27714), .B0(n28522), .C0(n27353), .Y(
        n27354) );
  AOI211XL U6359 ( .A0(n28143), .A1(n27507), .B0(n28291), .C0(n27284), .Y(
        n27285) );
  AOI211XL U6360 ( .A0(n28143), .A1(n27531), .B0(n28320), .C0(n27292), .Y(
        n27293) );
  AOI211XL U6361 ( .A0(n28143), .A1(n27665), .B0(n28466), .C0(n27337), .Y(
        n27338) );
  AOI211XL U6362 ( .A0(n28143), .A1(n27702), .B0(n28508), .C0(n27349), .Y(
        n27350) );
  OAI21XL U6363 ( .A0(n20350), .A1(n20345), .B0(n20344), .Y(n20347) );
  OAI21XL U6364 ( .A0(n17072), .A1(n14011), .B0(n16818), .Y(n14013) );
  OAI21XL U6365 ( .A0(n17196), .A1(n17182), .B0(n17181), .Y(n17186) );
  OAI21XL U6366 ( .A0(n18649), .A1(n18700), .B0(n18703), .Y(n6269) );
  OAI21XL U6367 ( .A0(n17196), .A1(n17189), .B0(n17194), .Y(n17192) );
  OAI21XL U6368 ( .A0(n25016), .A1(n25011), .B0(n6343), .Y(n6365) );
  OAI21XL U6369 ( .A0(n20353), .A1(n20065), .B0(n20311), .Y(n14891) );
  OAI21XL U6370 ( .A0(n17476), .A1(n17470), .B0(n17469), .Y(n17473) );
  OAI2BB1XL U6371 ( .A0N(n7729), .A1N(n21946), .B0(n7730), .Y(n14582) );
  AOI2BB1XL U6372 ( .A0N(n17632), .A1N(n7215), .B0(n17633), .Y(n17636) );
  OAI21X2 U6373 ( .A0(n6237), .A1(n24371), .B0(n24370), .Y(n6338) );
  NAND3X1 U6374 ( .A(n7857), .B(n7856), .C(n14864), .Y(n6122) );
  OAI32X4 U6375 ( .A0(n7305), .A1(C_sel_reg[8]), .A2(n28672), .B0(n14998), 
        .B1(n11633), .Y(n16570) );
  BUFX3 U6376 ( .A(n5933), .Y(n15557) );
  INVX4 U6377 ( .A(n5813), .Y(n16344) );
  OAI21XL U6378 ( .A0(Q7[11]), .A1(n5927), .B0(n27123), .Y(n27566) );
  OAI21XL U6379 ( .A0(Q7[13]), .A1(n5927), .B0(n27131), .Y(n27578) );
  OAI21XL U6380 ( .A0(Q7[22]), .A1(n5927), .B0(n27168), .Y(n27633) );
  OAI21XL U6381 ( .A0(Q7[24]), .A1(n5927), .B0(n27176), .Y(n27645) );
  OAI21XL U6382 ( .A0(Q7[25]), .A1(n5927), .B0(n27180), .Y(n27651) );
  OAI21XL U6383 ( .A0(Q7[12]), .A1(n5927), .B0(n27127), .Y(n27572) );
  OAI21XL U6384 ( .A0(Q7[16]), .A1(n5840), .B0(n27143), .Y(n27596) );
  OAI21XL U6385 ( .A0(Q7[21]), .A1(n5927), .B0(n27164), .Y(n27626) );
  OAI21XL U6386 ( .A0(Q7[39]), .A1(n5927), .B0(n27220), .Y(n27724) );
  OAI21XL U6387 ( .A0(Q7[40]), .A1(n5927), .B0(n27224), .Y(n27730) );
  OAI21XL U6388 ( .A0(Q7[41]), .A1(n5840), .B0(n27228), .Y(n27736) );
  OAI21XL U6389 ( .A0(Q7[42]), .A1(n5927), .B0(n27232), .Y(n27742) );
  OAI21XL U6390 ( .A0(Q7[49]), .A1(n5927), .B0(n27261), .Y(n27785) );
  OAI21XL U6391 ( .A0(Q7[14]), .A1(n5840), .B0(n27135), .Y(n27584) );
  OAI21XL U6392 ( .A0(Q7[15]), .A1(n5840), .B0(n27139), .Y(n27590) );
  OAI21XL U6393 ( .A0(Q7[17]), .A1(n5840), .B0(n27147), .Y(n27602) );
  OAI21XL U6394 ( .A0(Q7[47]), .A1(n5840), .B0(n27253), .Y(n27773) );
  OAI21XL U6395 ( .A0(Q7[48]), .A1(n5840), .B0(n27257), .Y(n27779) );
  INVX1 U6396 ( .A(n19072), .Y(n19100) );
  OAI21XL U6397 ( .A0(n22773), .A1(n14131), .B0(n7296), .Y(n22771) );
  OAI21XL U6398 ( .A0(n17491), .A1(n17480), .B0(n17479), .Y(n17489) );
  OAI21XL U6399 ( .A0(n16823), .A1(n16811), .B0(n16810), .Y(n16821) );
  INVXL U6400 ( .A(n19392), .Y(n19404) );
  OAI21XL U6401 ( .A0(Q6[42]), .A1(n5840), .B0(n27232), .Y(n27741) );
  OAI21XL U6402 ( .A0(Q6[49]), .A1(n5927), .B0(n27261), .Y(n27789) );
  OAI2BB1X1 U6403 ( .A0N(n7291), .A1N(n7753), .B0(n6366), .Y(n25016) );
  AOI21X2 U6404 ( .A0(n19785), .A1(n6652), .B0(n6658), .Y(n19793) );
  NAND2X1 U6405 ( .A(n7377), .B(n7379), .Y(n6419) );
  OAI21X2 U6406 ( .A0(n22597), .A1(n6238), .B0(n6800), .Y(n6799) );
  NAND2XL U6407 ( .A(n7187), .B(n6949), .Y(n6128) );
  CLKINVX3 U6408 ( .A(n25123), .Y(n25528) );
  CLKINVX3 U6409 ( .A(n15027), .Y(n15025) );
  INVX1 U6410 ( .A(n16416), .Y(n7125) );
  CLKINVX3 U6411 ( .A(n27281), .Y(n28168) );
  OAI21XL U6412 ( .A0(n7167), .A1(n6519), .B0(n8687), .Y(n6602) );
  AND2X2 U6413 ( .A(n6949), .B(n7188), .Y(n6127) );
  INVX1 U6414 ( .A(n14974), .Y(n14897) );
  OAI21XL U6415 ( .A0(n25290), .A1(n12401), .B0(n12400), .Y(n12402) );
  NAND2X2 U6416 ( .A(n6777), .B(n24672), .Y(n24701) );
  CLKINVX3 U6417 ( .A(n27390), .Y(n27431) );
  NOR2X2 U6418 ( .A(n22301), .B(n6760), .Y(n6759) );
  OAI21X2 U6419 ( .A0(n25534), .A1(n25523), .B0(n25522), .Y(n25531) );
  OAI21X2 U6420 ( .A0(n6697), .A1(n22175), .B0(n22174), .Y(n22180) );
  OAI2BB1X1 U6421 ( .A0N(n20332), .A1N(n7896), .B0(n20331), .Y(n7491) );
  OAI21XL U6422 ( .A0(n19407), .A1(n7712), .B0(n7711), .Y(n19429) );
  INVX1 U6423 ( .A(n21946), .Y(n22972) );
  OAI21XL U6424 ( .A0(n17181), .A1(n17183), .B0(n17184), .Y(n9603) );
  INVX1 U6425 ( .A(n24414), .Y(n22456) );
  NAND2BX1 U6426 ( .AN(n12334), .B(n29008), .Y(n16629) );
  OAI21XL U6427 ( .A0(n17456), .A1(n9541), .B0(n9540), .Y(n7411) );
  OAI2BB1X1 U6428 ( .A0N(n8630), .A1N(n7537), .B0(n16636), .Y(n7536) );
  NAND2X1 U6429 ( .A(n9147), .B(n6276), .Y(n6277) );
  AOI2BB1X1 U6430 ( .A0N(n17063), .A1N(n13966), .B0(n13974), .Y(n17058) );
  AOI21X1 U6431 ( .A0(n22359), .A1(n22318), .B0(n22317), .Y(n22331) );
  OAI21X1 U6432 ( .A0(n14970), .A1(n16787), .B0(n14969), .Y(n6683) );
  OAI21XL U6433 ( .A0(n7478), .A1(n20327), .B0(n20326), .Y(n20328) );
  NOR2X1 U6434 ( .A(n5953), .B(n6874), .Y(n5952) );
  XOR2X1 U6435 ( .A(n6561), .B(n8461), .Y(n19790) );
  OR3XL U6436 ( .A(A_sel_reg[0]), .B(n27236), .C(C_sel_reg[1]), .Y(n14980) );
  OAI21XL U6437 ( .A0(n13457), .A1(n24478), .B0(n13456), .Y(n24450) );
  OAI21XL U6438 ( .A0(n6073), .A1(n17644), .B0(n6072), .Y(n14505) );
  XOR2X1 U6439 ( .A(n12361), .B(n12360), .Y(n25286) );
  OAI21XL U6440 ( .A0(n13462), .A1(n24452), .B0(n13461), .Y(n13463) );
  AND2X2 U6441 ( .A(n13561), .B(n7553), .Y(n6151) );
  OAI21XL U6442 ( .A0(n19073), .A1(n9719), .B0(n9718), .Y(n7677) );
  OAI21XL U6443 ( .A0(n14495), .A1(n14491), .B0(n14492), .Y(n7251) );
  OAI21XL U6444 ( .A0(n17627), .A1(n6038), .B0(n14501), .Y(n6037) );
  NOR2X1 U6445 ( .A(n5845), .B(n20041), .Y(n20327) );
  OAI21XL U6446 ( .A0(n14483), .A1(n25145), .B0(n7041), .Y(n6508) );
  NAND2BX1 U6447 ( .AN(n19749), .B(n6688), .Y(n19870) );
  NAND2XL U6448 ( .A(n6594), .B(n8673), .Y(n16655) );
  NAND2X1 U6449 ( .A(n6544), .B(n24435), .Y(n6229) );
  INVX1 U6450 ( .A(n17032), .Y(n7095) );
  OAI21X1 U6451 ( .A0(n19235), .A1(n7038), .B0(n14857), .Y(n7903) );
  AOI21X1 U6452 ( .A0(n14967), .A1(n16794), .B0(n6086), .Y(n16787) );
  OAI21XL U6453 ( .A0(n8639), .A1(n8635), .B0(n8636), .Y(n6561) );
  XNOR2X2 U6454 ( .A(n6804), .B(n13191), .Y(n21946) );
  OAI21XL U6455 ( .A0(n13524), .A1(n13999), .B0(n13523), .Y(n13525) );
  OAI21XL U6456 ( .A0(n14862), .A1(n14858), .B0(n14859), .Y(n7808) );
  OAI21XL U6457 ( .A0(n9509), .A1(n17503), .B0(n9508), .Y(n17477) );
  OAI21XL U6458 ( .A0(n9596), .A1(n13723), .B0(n9595), .Y(n9597) );
  OAI21XL U6459 ( .A0(n23932), .A1(n23931), .B0(n23930), .Y(n23933) );
  OAI21XL U6460 ( .A0(n17108), .A1(n13887), .B0(n13886), .Y(n13888) );
  OAI21XL U6461 ( .A0(n16799), .A1(n14965), .B0(n14964), .Y(n16794) );
  INVXL U6462 ( .A(n24692), .Y(n5846) );
  OAI21XL U6463 ( .A0(n9144), .A1(n25009), .B0(n9143), .Y(n9145) );
  OAI21XL U6464 ( .A0(n25208), .A1(n14390), .B0(n14389), .Y(n14391) );
  OAI21XL U6465 ( .A0(n13991), .A1(n13990), .B0(n13989), .Y(n5989) );
  XOR2X1 U6466 ( .A(n8639), .B(n8638), .Y(n12334) );
  NAND2BX1 U6467 ( .AN(n25703), .B(n25705), .Y(n12234) );
  XNOR2X2 U6468 ( .A(n11551), .B(n11550), .Y(U2_U0_z0[11]) );
  AOI21X1 U6469 ( .A0(n11506), .A1(n6178), .B0(n11505), .Y(n11511) );
  NOR2X1 U6470 ( .A(n7252), .B(n14269), .Y(n14495) );
  NOR2BX1 U6471 ( .AN(n25715), .B(n6476), .Y(n25700) );
  NOR2X1 U6472 ( .A(n9596), .B(n13722), .Y(n9598) );
  NOR2XL U6473 ( .A(n14138), .B(n14131), .Y(n14140) );
  AOI21X1 U6474 ( .A0(n7540), .A1(n26904), .B0(n26947), .Y(n7539) );
  NOR2X1 U6475 ( .A(n28707), .B(n27236), .Y(n11920) );
  AOI21X1 U6476 ( .A0(n24743), .A1(n24745), .B0(n6778), .Y(n24731) );
  OAI21XL U6477 ( .A0(n9546), .A1(n9542), .B0(n9543), .Y(n9349) );
  OAI21XL U6478 ( .A0(n19764), .A1(n19848), .B0(n6651), .Y(n19822) );
  OAI21XL U6479 ( .A0(n14872), .A1(n20419), .B0(n14871), .Y(n20388) );
  OAI21XL U6480 ( .A0(n22001), .A1(n14559), .B0(n14558), .Y(n21978) );
  OAI21XL U6481 ( .A0(n13518), .A1(n24900), .B0(n13517), .Y(n13996) );
  OAI21XL U6482 ( .A0(n9707), .A1(n19104), .B0(n9706), .Y(n9708) );
  OAI21XL U6483 ( .A0(n14046), .A1(n22501), .B0(n14045), .Y(n22442) );
  OAI21XL U6484 ( .A0(n22658), .A1(n12578), .B0(n12577), .Y(n12579) );
  NAND2BX1 U6485 ( .AN(n24662), .B(n22932), .Y(n23017) );
  OAI21XL U6486 ( .A0(n25508), .A1(n25554), .B0(n25507), .Y(n25509) );
  OAI21XL U6487 ( .A0(n19091), .A1(n9714), .B0(n9713), .Y(n19082) );
  XOR2X1 U6488 ( .A(n12280), .B(n12277), .Y(n14577) );
  CLKINVX4 U6489 ( .A(n27122), .Y(n27236) );
  XOR2X1 U6490 ( .A(n8634), .B(n6964), .Y(n12332) );
  NOR2X1 U6491 ( .A(n13524), .B(n13998), .Y(n13526) );
  AOI21X1 U6492 ( .A0(n13983), .A1(n13982), .B0(n13981), .Y(n13991) );
  AOI21X1 U6493 ( .A0(n24094), .A1(n6986), .B0(n24093), .Y(n24157) );
  AOI21X1 U6494 ( .A0(n8033), .A1(n9141), .B0(n8032), .Y(n25009) );
  AOI21X1 U6495 ( .A0(n6641), .A1(n6648), .B0(n6562), .Y(n8639) );
  XNOR2X2 U6496 ( .A(n9227), .B(n9218), .Y(n24677) );
  XOR2X2 U6497 ( .A(n13660), .B(n13650), .Y(n19233) );
  XNOR2X2 U6498 ( .A(n13485), .B(n13484), .Y(n22453) );
  XNOR2X1 U6499 ( .A(n6359), .B(n9230), .Y(n24692) );
  XOR2X2 U6500 ( .A(n13983), .B(n6720), .Y(n20032) );
  OAI21XL U6501 ( .A0(n11389), .A1(n11231), .B0(n11230), .Y(n11234) );
  CLKINVX3 U6502 ( .A(OP_done1), .Y(n27213) );
  OAI21XL U6503 ( .A0(n6878), .A1(n10705), .B0(n10704), .Y(n10708) );
  OAI21XL U6504 ( .A0(n9214), .A1(n9213), .B0(n9212), .Y(n9227) );
  NAND2BX2 U6505 ( .AN(n24662), .B(n24642), .Y(n24745) );
  INVXL U6506 ( .A(n25151), .Y(n21794) );
  OAI21XL U6507 ( .A0(n14477), .A1(n14473), .B0(n14474), .Y(n14481) );
  OAI21XL U6508 ( .A0(n22025), .A1(n14544), .B0(n14543), .Y(n14545) );
  OAI21XL U6509 ( .A0(n8929), .A1(n25072), .B0(n8928), .Y(n25048) );
  INVX1 U6510 ( .A(n20047), .Y(n5850) );
  OAI21XL U6511 ( .A0(n18704), .A1(n18703), .B0(n18702), .Y(n18705) );
  OAI21XL U6512 ( .A0(n12889), .A1(n17699), .B0(n12888), .Y(n17666) );
  XOR2X1 U6513 ( .A(n9161), .B(n9160), .Y(n24679) );
  OAI21XL U6514 ( .A0(n18594), .A1(n18593), .B0(n18592), .Y(n18706) );
  ADDFX2 U6515 ( .A(n18864), .B(n18863), .CI(U2_A_i_d[21]), .CO(n18866), .S(
        n18820) );
  NAND2BX1 U6516 ( .AN(n20007), .B(n5859), .Y(n7005) );
  XOR2X2 U6517 ( .A(n11287), .B(n6979), .Y(U0_U1_z0[17]) );
  XNOR2X2 U6518 ( .A(n11260), .B(n11259), .Y(U0_U1_z0[22]) );
  XNOR2X2 U6519 ( .A(n8264), .B(n8263), .Y(U1_U2_z0[21]) );
  OAI21X1 U6520 ( .A0(n24039), .A1(n24038), .B0(n24037), .Y(n24094) );
  NAND3BX1 U6521 ( .AN(n13513), .B(n24919), .C(n7326), .Y(n6553) );
  OAI2BB1X1 U6522 ( .A0N(W3[15]), .A1N(n7986), .B0(n6179), .Y(n10101) );
  XNOR2X1 U6523 ( .A(n9233), .B(n9224), .Y(n24687) );
  OAI21XL U6524 ( .A0(n6878), .A1(n8261), .B0(n8260), .Y(n8264) );
  INVX2 U6525 ( .A(n14948), .Y(n5817) );
  OAI21XL U6526 ( .A0(n6878), .A1(n10725), .B0(n10724), .Y(n10730) );
  INVX1 U6527 ( .A(n25174), .Y(n21781) );
  INVXL U6528 ( .A(n20002), .Y(n14946) );
  INVX1 U6529 ( .A(n14953), .Y(n5862) );
  INVXL U6530 ( .A(n14086), .Y(n13452) );
  INVX1 U6531 ( .A(n19993), .Y(n5859) );
  INVX1 U6532 ( .A(n24664), .Y(n5819) );
  INVXL U6533 ( .A(n14562), .Y(n6313) );
  INVX1 U6534 ( .A(n19776), .Y(n12327) );
  CLKINVX3 U6535 ( .A(n24665), .Y(n24640) );
  XOR2X1 U6536 ( .A(n6398), .B(n10081), .Y(U2_U0_z2[12]) );
  AND2X2 U6537 ( .A(n19537), .B(n19639), .Y(n6111) );
  XOR2XL U6538 ( .A(n9792), .B(n10039), .Y(U2_U0_z2[10]) );
  XOR2X1 U6539 ( .A(n13970), .B(n6692), .Y(n20047) );
  XOR2X1 U6540 ( .A(n13181), .B(n13177), .Y(n22965) );
  AOI21X2 U6541 ( .A0(n7622), .A1(n6484), .B0(n7663), .Y(n9546) );
  XOR2X1 U6542 ( .A(n7145), .B(n13958), .Y(n20050) );
  OAI21X2 U6543 ( .A0(n7142), .A1(n10880), .B0(n10879), .Y(n10883) );
  OAI21X1 U6544 ( .A0(n6712), .A1(n10541), .B0(n10540), .Y(n10546) );
  XOR2X2 U6545 ( .A(n10788), .B(n6918), .Y(U1_U2_z0[13]) );
  XOR2X1 U6546 ( .A(n13941), .B(n7153), .Y(n14956) );
  XOR2X2 U6547 ( .A(n10893), .B(n6962), .Y(U0_U2_z0[23]) );
  XNOR2X2 U6548 ( .A(n10745), .B(n10744), .Y(U1_U2_z0[19]) );
  XOR2X1 U6549 ( .A(n10083), .B(n10082), .Y(U2_U0_z1[12]) );
  XOR2X1 U6550 ( .A(n14477), .B(n14476), .Y(n25140) );
  XOR2X2 U6551 ( .A(n10793), .B(n6965), .Y(U1_U2_z0[12]) );
  XNOR2X2 U6552 ( .A(n10736), .B(n10735), .Y(U1_U2_z0[20]) );
  XNOR2X2 U6553 ( .A(n9569), .B(n9568), .Y(U1_U0_z0[24]) );
  XNOR2X2 U6554 ( .A(n10563), .B(n10562), .Y(U1_U0_z0[21]) );
  NAND2BX1 U6555 ( .AN(n10100), .B(n6180), .Y(n6179) );
  XOR2X2 U6556 ( .A(n7562), .B(n6976), .Y(U1_U1_z0[20]) );
  XOR2X2 U6557 ( .A(n14848), .B(n6094), .Y(n20041) );
  OAI21XL U6558 ( .A0(n7148), .A1(n10558), .B0(n10557), .Y(n10563) );
  INVX2 U6559 ( .A(n14053), .Y(n14133) );
  OAI21XL U6560 ( .A0(n10817), .A1(n10784), .B0(n10783), .Y(n10788) );
  OAI21XL U6561 ( .A0(n7197), .A1(n10875), .B0(n10874), .Y(n10878) );
  OAI21XL U6562 ( .A0(n11030), .A1(n10899), .B0(n10898), .Y(n10904) );
  CMPR32X1 U6563 ( .A(n23577), .B(n23576), .C(U2_A_i_d[9]), .CO(n23578), .S(
        n23527) );
  INVX1 U6564 ( .A(n20013), .Y(n14835) );
  OAI21XL U6565 ( .A0(n10477), .A1(n10440), .B0(n10439), .Y(n10445) );
  OAI21XL U6566 ( .A0(n10477), .A1(n10429), .B0(n10428), .Y(n10434) );
  OAI21XL U6567 ( .A0(n9792), .A1(n9789), .B0(n9790), .Y(n9772) );
  OR2X2 U6568 ( .A(n24662), .B(n24642), .Y(n8033) );
  OAI21XL U6569 ( .A0(n11348), .A1(n11315), .B0(n11314), .Y(n11320) );
  INVXL U6570 ( .A(n14945), .Y(n20006) );
  OAI21XL U6571 ( .A0(n10083), .A1(n10033), .B0(n10032), .Y(n10036) );
  XOR2X1 U6572 ( .A(n13082), .B(n7004), .Y(n14955) );
  XNOR2X1 U6573 ( .A(n11154), .B(n11153), .Y(U1_U1_z0[11]) );
  ADDFX2 U6574 ( .A(n17978), .B(n17977), .CI(U2_A_i_d[5]), .CO(n17979), .S(
        n17941) );
  AOI21X2 U6575 ( .A0(n6856), .A1(n5761), .B0(n6821), .Y(U1_U1_z1[16]) );
  OAI21XL U6576 ( .A0(n8892), .A1(n25111), .B0(n8891), .Y(n25093) );
  NOR2X1 U6577 ( .A(n22922), .B(n7565), .Y(n23068) );
  XOR2X1 U6578 ( .A(n13012), .B(n13011), .Y(n14953) );
  INVXL U6579 ( .A(n7696), .Y(n6190) );
  XOR2X1 U6580 ( .A(n6245), .B(n13165), .Y(n22959) );
  OAI21X1 U6581 ( .A0(n10522), .A1(n8228), .B0(n8227), .Y(n8231) );
  OAI21X2 U6582 ( .A0(n6982), .A1(n13908), .B0(n7459), .Y(n19993) );
  XNOR2X1 U6583 ( .A(n10057), .B(n10056), .Y(U2_U0_z1[9]) );
  NAND2X2 U6584 ( .A(n6642), .B(n6667), .Y(n6648) );
  XOR2X1 U6585 ( .A(n6668), .B(n8623), .Y(n19776) );
  OAI21X1 U6586 ( .A0(n10643), .A1(n8278), .B0(n8277), .Y(n8281) );
  XNOR2X1 U6587 ( .A(n13146), .B(n13145), .Y(n22957) );
  AOI21X2 U6588 ( .A0(n9196), .A1(n9180), .B0(n9195), .Y(n9214) );
  XOR2X2 U6589 ( .A(n8315), .B(n11585), .Y(U2_U0_z0[4]) );
  NAND2X1 U6590 ( .A(n7405), .B(n7404), .Y(n21524) );
  ADDFHX1 U6591 ( .A(n26760), .B(n26759), .CI(U2_A_r_d[18]), .CO(n26761), .S(
        n26705) );
  ADDFHX1 U6592 ( .A(n24041), .B(n24040), .CI(U2_A_i_d[17]), .CO(n24042), .S(
        n23984) );
  ADDFHX1 U6593 ( .A(n26461), .B(n26460), .CI(U2_A_r_d[13]), .CO(n26462), .S(
        n26406) );
  OAI21X2 U6594 ( .A0(n8006), .A1(n6898), .B0(n7764), .Y(n10187) );
  NOR2X1 U6595 ( .A(n6645), .B(n8626), .Y(n6644) );
  ADDFHX1 U6596 ( .A(n26516), .B(n26515), .CI(U2_A_r_d[14]), .CO(n26517), .S(
        n26463) );
  ADDFHX1 U6597 ( .A(n24098), .B(n24097), .CI(U2_A_i_d[18]), .CO(n24099), .S(
        n24043) );
  XNOR2X2 U6598 ( .A(n9525), .B(n9524), .Y(n13709) );
  ADDFHX1 U6599 ( .A(n18711), .B(n18710), .CI(U2_A_i_d[18]), .CO(n18712), .S(
        n18653) );
  ADDFHX1 U6600 ( .A(n5887), .B(n5888), .CI(U2_A_i_d[14]), .CO(n18496), .S(
        n18410) );
  ADDFHX1 U6601 ( .A(n18547), .B(n18546), .CI(U2_A_i_d[15]), .CO(n18548), .S(
        n18497) );
  ADDFHX1 U6602 ( .A(n18768), .B(n18767), .CI(U2_A_i_d[19]), .CO(n18769), .S(
        n18713) );
  INVX1 U6603 ( .A(n23981), .Y(n18595) );
  INVXL U6604 ( .A(n23937), .Y(n18547) );
  INVXL U6605 ( .A(n23871), .Y(n5887) );
  INVX1 U6606 ( .A(n23936), .Y(n18546) );
  INVX1 U6607 ( .A(n24098), .Y(n18711) );
  INVX1 U6608 ( .A(n24159), .Y(n18767) );
  INVX2 U6609 ( .A(n11557), .Y(n11582) );
  INVX1 U6610 ( .A(n14951), .Y(n5869) );
  OAI21XL U6611 ( .A0(n10477), .A1(n10447), .B0(n10446), .Y(n10451) );
  OAI21XL U6612 ( .A0(n7910), .A1(n13603), .B0(n7908), .Y(n7925) );
  INVX1 U6613 ( .A(n14031), .Y(n14076) );
  XOR2X1 U6614 ( .A(n10177), .B(n10176), .Y(U0_U0_z1[10]) );
  OAI21XL U6615 ( .A0(n10477), .A1(n10474), .B0(n10475), .Y(n10473) );
  CLKINVX3 U6616 ( .A(n14833), .Y(n7843) );
  INVXL U6617 ( .A(n9690), .Y(n13691) );
  INVXL U6618 ( .A(n19767), .Y(n6617) );
  OAI21XL U6619 ( .A0(n10097), .A1(n10096), .B0(n10095), .Y(n10098) );
  MXI2X1 U6620 ( .A(n7892), .B(n7160), .S0(n14800), .Y(n6104) );
  OAI2BB1XL U6621 ( .A0N(n11149), .A1N(n11107), .B0(n11148), .Y(n11154) );
  XOR2X1 U6622 ( .A(n13573), .B(n6972), .Y(n19272) );
  INVXL U6623 ( .A(n13082), .Y(n13585) );
  OAI2BB1X2 U6624 ( .A0N(n6297), .A1N(n6315), .B0(n6432), .Y(n9196) );
  XOR2X1 U6625 ( .A(n10489), .B(n10488), .Y(U0_U0_z0[6]) );
  NAND3X2 U6626 ( .A(n7683), .B(n7716), .C(n7682), .Y(n7696) );
  OAI21X1 U6627 ( .A0(W2[15]), .A1(n6943), .B0(n7234), .Y(n9931) );
  AOI21X2 U6628 ( .A0(n12264), .A1(n12259), .B0(n12263), .Y(n12273) );
  XNOR2X2 U6629 ( .A(n11599), .B(n11598), .Y(U2_U0_z0[2]) );
  INVXL U6630 ( .A(n13694), .Y(n9693) );
  NAND2X1 U6631 ( .A(n6424), .B(n8234), .Y(n10519) );
  XNOR2X2 U6632 ( .A(n10993), .B(n10992), .Y(U0_U2_z0[9]) );
  XOR2X1 U6633 ( .A(n13425), .B(n13424), .Y(n14040) );
  XOR2X2 U6634 ( .A(n10591), .B(n10590), .Y(U1_U0_z0[17]) );
  NAND2X1 U6635 ( .A(n7453), .B(n5993), .Y(n5992) );
  OAI21X1 U6636 ( .A0(n10817), .A1(n10767), .B0(n10766), .Y(n10771) );
  OAI2BB1X2 U6637 ( .A0N(n7773), .A1N(n7775), .B0(n7227), .Y(n24665) );
  OAI21X1 U6638 ( .A0(n11507), .A1(n11515), .B0(n11508), .Y(n7778) );
  NOR2X2 U6639 ( .A(n6643), .B(n8452), .Y(n6642) );
  XNOR2X2 U6640 ( .A(n7738), .B(n9089), .Y(n24661) );
  XOR2X2 U6641 ( .A(n6750), .B(n7953), .Y(n22932) );
  OAI22X2 U6642 ( .A0(n6063), .A1(n5991), .B0(n7900), .B1(n13940), .Y(n7899)
         );
  XOR2X2 U6643 ( .A(n6290), .B(n12643), .Y(n22931) );
  XOR2X2 U6644 ( .A(n6415), .B(n6970), .Y(n14086) );
  XOR2X2 U6645 ( .A(n6399), .B(n10046), .Y(U2_U0_z2[7]) );
  XOR2X2 U6646 ( .A(n13141), .B(n12633), .Y(n22933) );
  XOR2X2 U6647 ( .A(n7706), .B(n14428), .Y(n25162) );
  XOR2X2 U6648 ( .A(n13420), .B(n13419), .Y(n6228) );
  XOR2X1 U6649 ( .A(n7694), .B(n9467), .Y(n9694) );
  XOR2X2 U6650 ( .A(n6154), .B(n12991), .Y(n13037) );
  CLKINVX3 U6651 ( .A(n9504), .Y(n13694) );
  XNOR2X1 U6652 ( .A(n8208), .B(AOPB[26]), .Y(U0_U0_z0[0]) );
  INVX1 U6653 ( .A(n12963), .Y(n14932) );
  OAI21XL U6654 ( .A0(n13913), .A1(n6051), .B0(n6024), .Y(n6023) );
  INVX2 U6655 ( .A(n6597), .Y(n19751) );
  OAI21XL U6656 ( .A0(n10643), .A1(n10639), .B0(n10640), .Y(n10638) );
  INVX1 U6657 ( .A(n14826), .Y(n20003) );
  INVX1 U6658 ( .A(n14927), .Y(n19977) );
  OAI21XL U6659 ( .A0(n11348), .A1(n11344), .B0(n11345), .Y(n9650) );
  OAI21XL U6660 ( .A0(n10997), .A1(n10939), .B0(n10938), .Y(n10944) );
  OAI21XL U6661 ( .A0(n10086), .A1(n10072), .B0(n10071), .Y(n10075) );
  OAI21XL U6662 ( .A0(n12611), .A1(n12607), .B0(n12608), .Y(n12605) );
  XOR2X1 U6663 ( .A(n6844), .B(n9003), .Y(n24631) );
  XOR2X1 U6664 ( .A(n13019), .B(n13033), .Y(n19541) );
  XOR2X1 U6665 ( .A(n7186), .B(n6940), .Y(n7410) );
  OAI21XL U6666 ( .A0(n10997), .A1(n10982), .B0(n10981), .Y(n10986) );
  OAI21XL U6667 ( .A0(n9758), .A1(n9757), .B0(n9756), .Y(n9759) );
  NAND2X2 U6668 ( .A(n6053), .B(n6052), .Y(n13908) );
  XOR2X1 U6669 ( .A(n12193), .B(n12192), .Y(n14547) );
  NAND2BX2 U6670 ( .AN(n6048), .B(n7200), .Y(n7153) );
  NOR2X2 U6671 ( .A(n7440), .B(n7438), .Y(n14800) );
  INVX1 U6672 ( .A(n9118), .Y(n9130) );
  CMPR22X1 U6673 ( .A(U2_U0_y2[32]), .B(U2_U0_y0[32]), .CO(n24159), .S(n24098)
         );
  INVXL U6674 ( .A(U2_B_i[22]), .Y(n11452) );
  OAI21X2 U6675 ( .A0(n13413), .A1(n13409), .B0(n13410), .Y(n6415) );
  OAI21X2 U6676 ( .A0(n9107), .A1(n9106), .B0(n9105), .Y(n6274) );
  XOR2X1 U6677 ( .A(n9472), .B(n9478), .Y(n9690) );
  XOR2X1 U6678 ( .A(n14823), .B(n14822), .Y(n20001) );
  OAI2BB1X2 U6679 ( .A0N(n13152), .A1N(n6808), .B0(n6806), .Y(n13161) );
  CMPR22X1 U6680 ( .A(U2_U0_y2[23]), .B(U2_U0_y0[23]), .CO(n23633), .S(n23577)
         );
  CMPR22X1 U6681 ( .A(U2_U0_y2[22]), .B(U2_U0_y0[22]), .CO(n23576), .S(n23525)
         );
  AOI21X2 U6682 ( .A0(n8449), .A1(n8585), .B0(n6611), .Y(n6667) );
  CMPR22X1 U6683 ( .A(U2_U0_y2[24]), .B(U2_U0_y0[24]), .CO(n23690), .S(n23634)
         );
  CMPR22X1 U6684 ( .A(U2_U0_y2[25]), .B(U2_U0_y0[25]), .CO(n23742), .S(n23691)
         );
  OAI21X1 U6685 ( .A0(n13880), .A1(n13890), .B0(n13893), .Y(n6057) );
  XOR2X1 U6686 ( .A(n7697), .B(n6919), .Y(n7627) );
  OAI21X1 U6687 ( .A0(n11002), .A1(n10998), .B0(n10999), .Y(n6408) );
  NAND3X1 U6688 ( .A(n7591), .B(n14439), .C(n7590), .Y(n6729) );
  XNOR2X1 U6689 ( .A(n8978), .B(n8977), .Y(n24617) );
  NAND2X1 U6690 ( .A(n6105), .B(n7258), .Y(n7371) );
  CMPR22X1 U6691 ( .A(U2_U0_y2[27]), .B(U2_U0_y0[27]), .CO(n23870), .S(n23796)
         );
  INVX1 U6692 ( .A(n7117), .Y(n7118) );
  OAI21X1 U6693 ( .A0(n9114), .A1(n9113), .B0(n9112), .Y(n6275) );
  XOR2X1 U6694 ( .A(n14806), .B(n6010), .Y(n14833) );
  XNOR2X1 U6695 ( .A(n10802), .B(n10801), .Y(U1_U2_z0[11]) );
  AOI21X1 U6696 ( .A0(n6535), .A1(n6793), .B0(n6767), .Y(n6766) );
  XNOR2X2 U6697 ( .A(n10047), .B(n10046), .Y(U2_U0_z1[7]) );
  XNOR2X1 U6698 ( .A(n13030), .B(n13029), .Y(n13035) );
  XOR2X2 U6699 ( .A(n6372), .B(n8970), .Y(n24621) );
  XOR2X2 U6700 ( .A(n5945), .B(n13859), .Y(n19980) );
  XOR2X1 U6701 ( .A(n6006), .B(n14815), .Y(n20005) );
  XOR2X1 U6702 ( .A(n8569), .B(n8566), .Y(n12313) );
  ADDFHX1 U6703 ( .A(n21424), .B(n21423), .CI(U2_A_r_d[18]), .CO(n21425), .S(
        n21364) );
  ADDFHX1 U6704 ( .A(n21530), .B(n21529), .CI(U2_A_r_d[20]), .CO(n21531), .S(
        n21482) );
  XOR2X2 U6705 ( .A(n6386), .B(n12198), .Y(n14553) );
  ADDHXL U6706 ( .A(U0_pipe2[16]), .B(n28781), .CO(n26560), .S(n26478) );
  ADDHXL U6707 ( .A(U1_pipe11[17]), .B(U1_pipe10[17]), .CO(n18567), .S(n18538)
         );
  ADDHXL U6708 ( .A(U1_pipe1[17]), .B(U1_pipe0[17]), .CO(n21293), .S(n21238)
         );
  ADDHXL U6709 ( .A(U0_pipe5[17]), .B(U0_pipe4[17]), .CO(n23965), .S(n23908)
         );
  ADDHXL U6710 ( .A(U0_pipe11[17]), .B(U0_pipe10[17]), .CO(n23975), .S(n23916)
         );
  ADDHXL U6711 ( .A(U0_pipe1[17]), .B(U0_pipe0[17]), .CO(n26632), .S(n26565)
         );
  ADDHXL U6712 ( .A(U1_pipe7[17]), .B(U1_pipe6[17]), .CO(n18587), .S(n18522)
         );
  ADDHXL U6713 ( .A(U1_pipe5[17]), .B(U1_pipe4[17]), .CO(n18577), .S(n18530)
         );
  INVX1 U6714 ( .A(n26759), .Y(n21423) );
  INVX1 U6715 ( .A(n26819), .Y(n21479) );
  AND2X2 U6716 ( .A(n9750), .B(n9749), .Y(n10046) );
  OAI21XL U6717 ( .A0(n9999), .A1(n9998), .B0(n9997), .Y(n10000) );
  INVXL U6718 ( .A(n19744), .Y(n19736) );
  INVX1 U6719 ( .A(n10215), .Y(n7581) );
  AOI2BB1X1 U6720 ( .A0N(n6400), .A1N(n9746), .B0(n9747), .Y(n9802) );
  XOR2X1 U6721 ( .A(n12571), .B(n12570), .Y(n22918) );
  NOR2X2 U6722 ( .A(n6155), .B(n6074), .Y(n13012) );
  CLKBUFX8 U6723 ( .A(U0_U0_z1[1]), .Y(n6879) );
  XOR2X1 U6724 ( .A(n12166), .B(n12165), .Y(n14533) );
  XOR2X1 U6725 ( .A(n13392), .B(n13391), .Y(n14074) );
  AOI21X2 U6726 ( .A0(n9123), .A1(n9102), .B0(n9101), .Y(n9114) );
  OAI2BB1XL U6727 ( .A0N(n8828), .A1N(n7221), .B0(n8965), .Y(n6372) );
  NAND2BX2 U6728 ( .AN(n8225), .B(n6428), .Y(n10373) );
  XOR2X1 U6729 ( .A(n13873), .B(n13861), .Y(n19974) );
  XOR2X1 U6730 ( .A(n9448), .B(n9447), .Y(n13687) );
  OAI21X2 U6731 ( .A0(n10177), .A1(n10131), .B0(n10130), .Y(n10132) );
  NAND2BX1 U6732 ( .AN(n7506), .B(n13593), .Y(n6042) );
  OAI21X1 U6733 ( .A0(n6006), .A1(n14812), .B0(n14813), .Y(n6108) );
  AOI21X2 U6734 ( .A0(n6395), .A1(n9747), .B0(n6392), .Y(n6250) );
  NAND2BX1 U6735 ( .AN(n13582), .B(n6090), .Y(n6089) );
  OAI21X2 U6736 ( .A0(n7423), .A1(n11579), .B0(n11575), .Y(n11558) );
  NAND2X1 U6737 ( .A(U2_B_i[16]), .B(n6213), .Y(n11531) );
  XNOR2X1 U6738 ( .A(n13427), .B(n13372), .Y(n14071) );
  XOR2X1 U6739 ( .A(n12926), .B(n12925), .Y(n12963) );
  BUFX4 U6740 ( .A(n6048), .Y(n5991) );
  OAI2BB1X2 U6741 ( .A0N(n7356), .A1N(n5870), .B0(n7355), .Y(n7725) );
  OAI21X2 U6742 ( .A0(n8619), .A1(n8621), .B0(n8622), .Y(n6611) );
  NOR2X1 U6743 ( .A(n8222), .B(n10447), .Y(n8224) );
  OAI21X2 U6744 ( .A0(n7803), .A1(n7443), .B0(n7439), .Y(n7438) );
  INVX1 U6745 ( .A(n11437), .Y(n11536) );
  OAI21X1 U6746 ( .A0(n11284), .A1(n11289), .B0(n11285), .Y(n11277) );
  OAI21XL U6747 ( .A0(n6270), .A1(n11427), .B0(n11411), .Y(U2_B_i[23]) );
  XOR2X2 U6748 ( .A(n6502), .B(n14373), .Y(n25212) );
  XOR2X2 U6749 ( .A(n9426), .B(n9425), .Y(n13683) );
  AOI21X1 U6750 ( .A0(n9472), .A1(n7699), .B0(n7698), .Y(n7697) );
  XNOR2X2 U6751 ( .A(n6678), .B(n8573), .Y(n6597) );
  ADDFHX1 U6752 ( .A(n21017), .B(n21016), .CI(U2_A_r_d[11]), .CO(n21018), .S(
        n20962) );
  ADDFHX1 U6753 ( .A(n20960), .B(n20959), .CI(U2_A_r_d[10]), .CO(n20961), .S(
        n20905) );
  XOR2X2 U6754 ( .A(n7633), .B(n6958), .Y(n9504) );
  INVX1 U6755 ( .A(n26461), .Y(n21122) );
  INVXL U6756 ( .A(n26516), .Y(n21191) );
  INVXL U6757 ( .A(n26404), .Y(n21071) );
  XOR2X1 U6758 ( .A(n6831), .B(n10332), .Y(U1_U2_z2[10]) );
  OAI21XL U6759 ( .A0(n14360), .A1(n14359), .B0(n14358), .Y(n14365) );
  INVX1 U6760 ( .A(n10137), .Y(n10138) );
  OAI21XL U6761 ( .A0(n6835), .A1(n10044), .B0(n10018), .Y(n10019) );
  XOR2XL U6762 ( .A(n6235), .B(BOPA[48]), .Y(n6234) );
  INVX2 U6763 ( .A(n6633), .Y(n8620) );
  NAND2BX2 U6764 ( .AN(n9479), .B(n7680), .Y(n9491) );
  AOI21X2 U6765 ( .A0(n14816), .A1(n14808), .B0(n14807), .Y(n6006) );
  AOI21X2 U6766 ( .A0(n13019), .A1(n13040), .B0(n13045), .Y(n5951) );
  CMPR22X1 U6767 ( .A(U2_U0_y1[33]), .B(U2_U0_y0[33]), .CO(n26866), .S(n26820)
         );
  AOI21X2 U6768 ( .A0(n9472), .A1(n7329), .B0(n9463), .Y(n7633) );
  OAI2BB1X1 U6769 ( .A0N(n7615), .A1N(n7614), .B0(n7613), .Y(n9448) );
  XOR2X1 U6770 ( .A(n13307), .B(n7009), .Y(n14066) );
  XOR2X1 U6771 ( .A(n13327), .B(n13326), .Y(n14056) );
  XOR2X1 U6772 ( .A(n6946), .B(n7620), .Y(n13681) );
  CMPR22X1 U6773 ( .A(U2_U0_y1[34]), .B(U2_U0_y0[34]), .CO(n26908), .S(n26867)
         );
  INVX1 U6774 ( .A(n6158), .Y(n10731) );
  OAI2BB1XL U6775 ( .A0N(n5901), .A1N(n8825), .B0(n8823), .Y(n8752) );
  XNOR2X1 U6776 ( .A(n9429), .B(n7628), .Y(n13682) );
  NOR2X2 U6777 ( .A(n12252), .B(n12255), .Y(n6452) );
  NAND2X1 U6778 ( .A(n9188), .B(n9150), .Y(n7336) );
  OAI21X2 U6779 ( .A0(n9807), .A1(n9780), .B0(n9781), .Y(n9747) );
  NOR2X1 U6780 ( .A(n9519), .B(n9521), .Y(n7355) );
  NOR2X1 U6781 ( .A(n11297), .B(n11305), .Y(n8338) );
  ADDHX2 U6782 ( .A(U2_U0_y1[32]), .B(U2_U0_y0[32]), .CO(n26819), .S(n26760)
         );
  OAI21X1 U6783 ( .A0(n9748), .A1(n9800), .B0(n9749), .Y(n6392) );
  AOI21X1 U6784 ( .A0(n7830), .A1(n12915), .B0(n12896), .Y(n6148) );
  NAND3X1 U6785 ( .A(n7146), .B(n13960), .C(n13950), .Y(n6482) );
  XOR2X1 U6786 ( .A(n6716), .B(n9375), .Y(n9659) );
  OAI21X1 U6787 ( .A0(n10587), .A1(n10593), .B0(n10588), .Y(n10580) );
  NOR2X1 U6788 ( .A(n9626), .B(U2_B_r[6]), .Y(n11573) );
  OAI21XL U6789 ( .A0(n6403), .A1(n11427), .B0(n11404), .Y(U2_B_i[19]) );
  OAI21XL U6790 ( .A0(n28713), .A1(n11430), .B0(n9621), .Y(U2_B_r[12]) );
  AND2X2 U6791 ( .A(n9988), .B(n9987), .Y(n6999) );
  OAI21XL U6792 ( .A0(n28712), .A1(n11430), .B0(n11406), .Y(U2_B_r[16]) );
  NAND2X1 U6793 ( .A(W3[20]), .B(W3[4]), .Y(n9807) );
  INVX2 U6794 ( .A(U2_B_i[7]), .Y(n9627) );
  NOR2X1 U6795 ( .A(n8195), .B(AOPC[41]), .Y(n11297) );
  NAND2X1 U6796 ( .A(n8203), .B(AOPC[36]), .Y(n11340) );
  INVX1 U6797 ( .A(n10220), .Y(n10221) );
  OAI21XL U6798 ( .A0(n10441), .A1(n10448), .B0(n10442), .Y(n10426) );
  NOR2X1 U6799 ( .A(n9333), .B(n9334), .Y(n9521) );
  OAI21XL U6800 ( .A0(n7159), .A1(n14794), .B0(n14795), .Y(n7806) );
  NOR2X1 U6801 ( .A(n12249), .B(n12248), .Y(n12255) );
  INVX1 U6802 ( .A(n11072), .Y(n6273) );
  INVXL U6803 ( .A(U2_B_i[12]), .Y(n9638) );
  NAND3X2 U6804 ( .A(n6085), .B(n6084), .C(n6049), .Y(n13873) );
  CMPR22X1 U6805 ( .A(U2_U0_y1[23]), .B(U2_U0_y0[23]), .CO(n26290), .S(n26242)
         );
  CMPR22X1 U6806 ( .A(U2_U0_y1[24]), .B(U2_U0_y0[24]), .CO(n26355), .S(n26291)
         );
  OAI21X2 U6807 ( .A0(n9099), .A1(n9028), .B0(n9027), .Y(n9188) );
  XNOR2X1 U6808 ( .A(n10331), .B(n10330), .Y(U1_U2_z1[8]) );
  OAI21X1 U6809 ( .A0(n9904), .A1(n9901), .B0(n9902), .Y(n9900) );
  OAI21XL U6810 ( .A0(n28748), .A1(n11430), .B0(n9618), .Y(U2_B_r[10]) );
  NOR2XL U6811 ( .A(n13138), .B(n13134), .Y(n13140) );
  OAI21X2 U6812 ( .A0(n9764), .A1(n9794), .B0(n9765), .Y(n6396) );
  OAI21X1 U6813 ( .A0(n12626), .A1(n12627), .B0(n6811), .Y(n13153) );
  NOR2X1 U6814 ( .A(n14438), .B(n14434), .Y(n14424) );
  AOI21X1 U6815 ( .A0(n13048), .A1(n12917), .B0(n12909), .Y(n12914) );
  AND2X1 U6816 ( .A(n5839), .B(n9832), .Y(n10144) );
  NOR2X2 U6817 ( .A(W3[21]), .B(W3[5]), .Y(n9780) );
  NOR2X1 U6818 ( .A(n8022), .B(W3[21]), .Y(n10017) );
  NAND2X1 U6819 ( .A(n8030), .B(W3[20]), .Y(n10059) );
  NOR2X1 U6820 ( .A(n7955), .B(AOPB[38]), .Y(n10435) );
  NAND2X1 U6821 ( .A(n7972), .B(W1[28]), .Y(n10213) );
  INVX1 U6822 ( .A(n10261), .Y(n10262) );
  INVX1 U6823 ( .A(n10307), .Y(n10308) );
  NAND2X1 U6824 ( .A(n14250), .B(n14251), .Y(n14435) );
  NAND2X2 U6825 ( .A(n8438), .B(n8439), .Y(n8602) );
  OAI21XL U6826 ( .A0(n12077), .A1(n12078), .B0(n12080), .Y(n12074) );
  OAI21XL U6827 ( .A0(n9820), .A1(n9860), .B0(n9821), .Y(n9867) );
  OAI21XL U6828 ( .A0(n13922), .A1(n7184), .B0(n13921), .Y(n7155) );
  NOR2X1 U6829 ( .A(n13274), .B(n13273), .Y(n13446) );
  OAI21XL U6830 ( .A0(n9403), .A1(n9369), .B0(n9368), .Y(n9379) );
  NAND2X2 U6831 ( .A(n6595), .B(n8562), .Y(n8575) );
  NOR2X1 U6832 ( .A(n9066), .B(n9065), .Y(n9084) );
  NOR2X1 U6833 ( .A(n13067), .B(n13066), .Y(n13081) );
  NAND2X1 U6834 ( .A(W3[18]), .B(W3[2]), .Y(n9794) );
  OAI21X2 U6835 ( .A0(n6289), .A1(n10313), .B0(n10312), .Y(n10314) );
  NAND2X2 U6836 ( .A(n7156), .B(n13919), .Y(n7871) );
  NOR2X1 U6837 ( .A(n14666), .B(n14667), .Y(n14804) );
  NOR2X1 U6838 ( .A(n8589), .B(n8592), .Y(n8446) );
  INVX1 U6839 ( .A(n7802), .Y(n7887) );
  NOR2X2 U6840 ( .A(n7788), .B(n13058), .Y(n13589) );
  XNOR2X1 U6841 ( .A(n14992), .B(n9937), .Y(U1_U2_z2[1]) );
  NOR2X1 U6842 ( .A(n14670), .B(n14671), .Y(n14798) );
  NOR2X1 U6843 ( .A(n9986), .B(n6459), .Y(n9726) );
  NAND2X1 U6844 ( .A(n8442), .B(n8443), .Y(n6665) );
  NOR2X1 U6845 ( .A(n7901), .B(n13046), .Y(n7912) );
  AOI21X2 U6846 ( .A0(n9991), .A1(n9990), .B0(n9973), .Y(n6829) );
  NOR2X1 U6847 ( .A(n13083), .B(n13084), .Y(n13577) );
  NOR2X2 U6848 ( .A(n9462), .B(n9323), .Y(n9480) );
  AOI21X1 U6849 ( .A0(n10216), .A1(n7170), .B0(n10203), .Y(n10212) );
  OAI21X1 U6850 ( .A0(n13894), .A1(n13893), .B0(n13892), .Y(n7477) );
  OAI21X1 U6851 ( .A0(n7389), .A1(n11427), .B0(n8241), .Y(U2_B_i[15]) );
  OAI21X1 U6852 ( .A0(n13909), .A1(n13914), .B0(n13910), .Y(n13923) );
  AOI21X1 U6853 ( .A0(n9875), .A1(n6755), .B0(n9874), .Y(n9927) );
  NOR2X1 U6854 ( .A(n10954), .B(n10960), .Y(n10946) );
  NAND2X1 U6855 ( .A(n6296), .B(n6326), .Y(n6325) );
  OAI21X1 U6856 ( .A0(n6287), .A1(n11418), .B0(n8307), .Y(U2_B_i[4]) );
  OAI21X1 U6857 ( .A0(n9492), .A1(n9498), .B0(n9493), .Y(n9481) );
  XOR2X2 U6858 ( .A(n9979), .B(n10242), .Y(U1_U1_z2[3]) );
  OAI21XL U6859 ( .A0(n29102), .A1(n11430), .B0(n8306), .Y(U2_B_r[2]) );
  NOR2X2 U6860 ( .A(n8104), .B(AOPB[27]), .Y(n10524) );
  NAND2X1 U6861 ( .A(n8068), .B(AOPD[32]), .Y(n10999) );
  NAND2X1 U6862 ( .A(W0[28]), .B(W0[12]), .Y(n9860) );
  NOR2X1 U6863 ( .A(n7973), .B(W0[28]), .Y(n10172) );
  XOR2X1 U6864 ( .A(n7781), .B(BOPA[41]), .Y(n7389) );
  NOR2BX2 U6865 ( .AN(n9978), .B(n7276), .Y(n10242) );
  NOR2X1 U6866 ( .A(n9325), .B(n9324), .Y(n9497) );
  NOR2X1 U6867 ( .A(n8438), .B(n8439), .Y(n8601) );
  NAND2X1 U6868 ( .A(n12982), .B(n12983), .Y(n13027) );
  NAND2X1 U6869 ( .A(n12987), .B(n12986), .Y(n13060) );
  NOR2X1 U6870 ( .A(n9329), .B(n9328), .Y(n9486) );
  OAI21XL U6871 ( .A0(n9881), .A1(n9942), .B0(n9882), .Y(n9924) );
  NAND2X1 U6872 ( .A(n9328), .B(n9329), .Y(n9487) );
  NAND2X2 U6873 ( .A(n9975), .B(n6828), .Y(n10261) );
  INVX1 U6874 ( .A(n9484), .Y(n7636) );
  XOR2XL U6875 ( .A(U1_U1_y1[31]), .B(U1_U1_y0[31]), .Y(n14666) );
  AOI21X2 U6876 ( .A0(n9315), .A1(n9437), .B0(n7695), .Y(n9461) );
  NOR2X2 U6877 ( .A(n13922), .B(n13918), .Y(n7156) );
  INVXL U6878 ( .A(n11601), .Y(n6326) );
  NOR2X2 U6879 ( .A(n9619), .B(n7777), .Y(n6225) );
  INVX1 U6880 ( .A(n10410), .Y(n6425) );
  INVXL U6881 ( .A(U2_B_i[2]), .Y(n8311) );
  NAND2X1 U6882 ( .A(W1[10]), .B(W1[26]), .Y(n9987) );
  NOR2X2 U6883 ( .A(n7400), .B(n8563), .Y(n8586) );
  INVXL U6884 ( .A(n6459), .Y(n9959) );
  NOR2XL U6885 ( .A(n9886), .B(n9938), .Y(n9875) );
  NAND2X1 U6886 ( .A(n10161), .B(n10160), .Y(n12002) );
  NOR2X1 U6887 ( .A(n13909), .B(n13913), .Y(n13919) );
  NOR2X1 U6888 ( .A(n10119), .B(n10131), .Y(n10121) );
  NOR2X1 U6889 ( .A(n10202), .B(n10219), .Y(n7170) );
  OAI21X1 U6890 ( .A0(n13848), .A1(n7046), .B0(n13852), .Y(n13796) );
  CMPR22X1 U6891 ( .A(U0_U1_y2[33]), .B(U0_U1_y0[33]), .CO(n12645), .S(n12641)
         );
  CMPR22X1 U6892 ( .A(U0_U1_y2[32]), .B(U0_U1_y0[32]), .CO(n12642), .S(n12630)
         );
  OAI21X1 U6893 ( .A0(n9892), .A1(n9932), .B0(n9893), .Y(n6755) );
  XOR2X2 U6894 ( .A(n9619), .B(n28713), .Y(n6420) );
  CMPR22X1 U6895 ( .A(U0_U1_y1[32]), .B(U0_U1_y0[32]), .CO(n9068), .S(n9065)
         );
  CMPR22X1 U6896 ( .A(U1_U2_y2[31]), .B(U1_U2_y0[31]), .CO(n13927), .S(n13924)
         );
  CMPR22X1 U6897 ( .A(U0_U1_y1[33]), .B(U0_U1_y0[33]), .CO(n9070), .S(n9067)
         );
  NOR2X1 U6898 ( .A(n9890), .B(n9892), .Y(n9885) );
  CMPR22X1 U6899 ( .A(U0_U1_y1[31]), .B(U0_U1_y0[31]), .CO(n9066), .S(n9063)
         );
  NOR2X1 U6900 ( .A(n9826), .B(n9856), .Y(n9814) );
  XNOR2X1 U6901 ( .A(U1_U1_y1[32]), .B(n6136), .Y(n14668) );
  NOR2X1 U6902 ( .A(n10200), .B(n10223), .Y(n10217) );
  XOR2X1 U6903 ( .A(U1_U1_y0[32]), .B(U1_U1_y2[32]), .Y(n13066) );
  INVX1 U6904 ( .A(n8048), .Y(n6461) );
  NAND2X1 U6905 ( .A(n7998), .B(W0[24]), .Y(n10134) );
  NOR2X2 U6906 ( .A(n8127), .B(BOPC[31]), .Y(n11187) );
  NOR2X2 U6907 ( .A(W2[10]), .B(W2[26]), .Y(n9938) );
  NAND2X1 U6908 ( .A(W2[8]), .B(W2[24]), .Y(n9932) );
  NAND2X1 U6909 ( .A(n7951), .B(W0[26]), .Y(n10130) );
  NOR2X2 U6910 ( .A(W1[27]), .B(W1[11]), .Y(n6459) );
  NAND2X1 U6911 ( .A(n8102), .B(AOPC[27]), .Y(n11397) );
  NAND2X1 U6912 ( .A(n7952), .B(W1[26]), .Y(n10218) );
  NOR2X1 U6913 ( .A(n8119), .B(BOPB[34]), .Y(n10639) );
  NOR2X1 U6914 ( .A(n8185), .B(BOPC[38]), .Y(n11128) );
  NOR2X1 U6915 ( .A(n8036), .B(W3[18]), .Y(n10072) );
  NAND2X1 U6916 ( .A(n13049), .B(n13050), .Y(n13073) );
  NAND2X1 U6917 ( .A(n12940), .B(n12941), .Y(n12977) );
  OAI21X2 U6918 ( .A0(n8305), .A1(n29106), .B0(n8304), .Y(U2_B_i[2]) );
  NOR2X1 U6919 ( .A(n8996), .B(n8995), .Y(n9016) );
  NOR2X1 U6920 ( .A(n12546), .B(n12545), .Y(n12562) );
  NOR2X1 U6921 ( .A(n12567), .B(n12566), .Y(n12585) );
  INVX1 U6922 ( .A(n9845), .Y(n9853) );
  NOR2X1 U6923 ( .A(n9019), .B(n9018), .Y(n9131) );
  INVX1 U6924 ( .A(n9974), .Y(n6828) );
  AOI21X2 U6925 ( .A0(n13851), .A1(n7469), .B0(n6034), .Y(n6049) );
  NOR2X1 U6926 ( .A(n12589), .B(n12588), .Y(n12607) );
  NOR2X2 U6927 ( .A(n9439), .B(n9444), .Y(n9315) );
  AOI21X2 U6928 ( .A0(n6071), .A1(n13803), .B0(n5983), .Y(n13852) );
  AOI21X2 U6929 ( .A0(n7544), .A1(n7531), .B0(n6604), .Y(n6603) );
  NOR2X1 U6930 ( .A(n13044), .B(n13039), .Y(n6873) );
  NOR2X2 U6931 ( .A(n10970), .B(n10974), .Y(n8320) );
  NOR2X2 U6932 ( .A(n13364), .B(n13366), .Y(n13383) );
  NAND2X1 U6933 ( .A(n13262), .B(n6911), .Y(n13389) );
  INVX1 U6934 ( .A(n10975), .Y(n6560) );
  NAND2BX1 U6935 ( .AN(n9331), .B(n7684), .Y(n9484) );
  NOR2X1 U6936 ( .A(n12978), .B(n12974), .Y(n12981) );
  AOI21X1 U6937 ( .A0(n6368), .A1(n8894), .B0(n6367), .Y(n8952) );
  NOR2X1 U6938 ( .A(n13304), .B(n13308), .Y(n13314) );
  NOR2X1 U6939 ( .A(n11015), .B(n11037), .Y(n7207) );
  OAI2BB1X2 U6940 ( .A0N(n7468), .A1N(n12797), .B0(n6026), .Y(n7522) );
  OAI21X2 U6941 ( .A0(n9477), .A1(n9473), .B0(n9474), .Y(n9463) );
  CMPR22X1 U6942 ( .A(U1_U0_y2[33]), .B(U1_U0_y0[33]), .CO(n8445), .S(n8442)
         );
  CMPR22X1 U6943 ( .A(U1_U0_y2[31]), .B(U1_U0_y0[31]), .CO(n8441), .S(n8438)
         );
  OAI21X2 U6944 ( .A0(n13020), .A1(n13032), .B0(n13021), .Y(n13045) );
  NOR2BX1 U6945 ( .AN(n14810), .B(n6134), .Y(n6133) );
  NOR2X2 U6946 ( .A(n8207), .B(AOPD[26]), .Y(n11035) );
  NOR2X2 U6947 ( .A(n8201), .B(AOPD[37]), .Y(n10974) );
  NOR2X1 U6948 ( .A(W2[24]), .B(W2[8]), .Y(n9890) );
  AND2X2 U6949 ( .A(n13847), .B(n13851), .Y(n7867) );
  XNOR2X1 U6950 ( .A(BOPA[27]), .B(BOPA[26]), .Y(n8301) );
  NOR2X2 U6951 ( .A(n13002), .B(n13003), .Y(n13020) );
  INVX1 U6952 ( .A(n9825), .Y(n7266) );
  OAI21XL U6953 ( .A0(n8900), .A1(n8917), .B0(n8901), .Y(n6367) );
  NOR2X2 U6954 ( .A(n13256), .B(n13255), .Y(n13374) );
  NOR2X2 U6955 ( .A(n12985), .B(n12984), .Y(n13016) );
  NAND2X1 U6956 ( .A(n13256), .B(n13255), .Y(n13373) );
  NAND2X1 U6957 ( .A(n13000), .B(n13001), .Y(n13032) );
  NOR2X2 U6958 ( .A(n6486), .B(n13254), .Y(n13304) );
  OAI21XL U6959 ( .A0(n6524), .A1(n12552), .B0(n12555), .Y(n12534) );
  INVXL U6960 ( .A(n12218), .Y(n7241) );
  NOR2X1 U6961 ( .A(n8957), .B(n6741), .Y(n8993) );
  NAND2X1 U6962 ( .A(n9312), .B(n9313), .Y(n9445) );
  OAI21XL U6963 ( .A0(n8833), .A1(n8832), .B0(n8831), .Y(n8935) );
  NAND2BX1 U6964 ( .AN(n7604), .B(n13254), .Y(n13305) );
  NAND2X1 U6965 ( .A(n8080), .B(AOPD[29]), .Y(n11016) );
  OAI21X1 U6966 ( .A0(n28682), .A1(n11428), .B0(n8302), .Y(U2_B_r[1]) );
  NAND2X1 U6967 ( .A(n13004), .B(n13005), .Y(n13043) );
  NAND2X1 U6968 ( .A(n13252), .B(n13253), .Y(n13309) );
  NAND2X1 U6969 ( .A(n14701), .B(n7797), .Y(n7308) );
  NOR2X2 U6970 ( .A(n8576), .B(n8581), .Y(n8564) );
  NOR2X2 U6971 ( .A(n14817), .B(n14820), .Y(n14808) );
  NOR2X1 U6972 ( .A(n13848), .B(n7046), .Y(n7868) );
  OAI21X1 U6973 ( .A0(n9897), .A1(n9902), .B0(n9898), .Y(n6283) );
  OAI21X1 U6974 ( .A0(n8840), .A1(n8852), .B0(n8841), .Y(n8894) );
  CMPR22X1 U6975 ( .A(U0_U2_y1[29]), .B(U0_U2_y0[29]), .CO(n9025), .S(n9022)
         );
  CMPR22X1 U6976 ( .A(U1_U2_y2[30]), .B(U1_U2_y0[30]), .CO(n13925), .S(n13902)
         );
  CMPR22X1 U6977 ( .A(U1_U2_y2[29]), .B(U1_U2_y0[29]), .CO(n13903), .S(n13900)
         );
  CMPR22X1 U6978 ( .A(U0_U1_y0[25]), .B(U0_U1_y2[25]), .CO(n12567), .S(n12564)
         );
  CMPR22X1 U6979 ( .A(U0_U1_y2[26]), .B(U0_U1_y0[26]), .CO(n12589), .S(n12566)
         );
  CMPR22X1 U6980 ( .A(U1_U2_y2[27]), .B(U1_U2_y0[27]), .CO(n13899), .S(n13897)
         );
  NOR2X2 U6981 ( .A(n7980), .B(W2[20]), .Y(n10315) );
  NAND2X1 U6982 ( .A(W2[6]), .B(W2[22]), .Y(n9902) );
  NOR2X1 U6983 ( .A(W2[4]), .B(W2[20]), .Y(n9905) );
  NOR2X2 U6984 ( .A(n8432), .B(n8433), .Y(n8576) );
  NOR2X2 U6985 ( .A(n9052), .B(n9053), .Y(n9119) );
  CLKINVX2 U6986 ( .A(n9839), .Y(n5932) );
  INVX1 U6987 ( .A(n10227), .Y(n10228) );
  NOR2X2 U6988 ( .A(n14661), .B(n14660), .Y(n14817) );
  OAI21XL U6989 ( .A0(n13323), .A1(n13328), .B0(n13324), .Y(n7230) );
  OAI21XL U6990 ( .A0(n8874), .A1(n8799), .B0(n8798), .Y(n8938) );
  OAI21XL U6991 ( .A0(n14298), .A1(n14303), .B0(n14299), .Y(n6497) );
  OAI21XL U6992 ( .A0(n13332), .A1(n13243), .B0(n13242), .Y(n13301) );
  NOR2X2 U6993 ( .A(n14767), .B(n14769), .Y(n7797) );
  NOR2X1 U6994 ( .A(n14653), .B(n14652), .Y(n14760) );
  NOR2X2 U6995 ( .A(n12179), .B(n12176), .Y(n6210) );
  NOR2X2 U6996 ( .A(n6066), .B(n6064), .Y(n7046) );
  NOR2X2 U6997 ( .A(n13865), .B(n13863), .Y(n13851) );
  NOR2X2 U6998 ( .A(n10266), .B(n10341), .Y(n7196) );
  NOR2X2 U6999 ( .A(n12802), .B(n12800), .Y(n7468) );
  NOR2X1 U7000 ( .A(n12928), .B(n12930), .Y(n7448) );
  NOR2X1 U7001 ( .A(n8430), .B(n8431), .Y(n8581) );
  OAI21X2 U7002 ( .A0(n8464), .A1(n8469), .B0(n8465), .Y(n8473) );
  NAND3BX1 U7003 ( .AN(n14632), .B(n7852), .C(n7851), .Y(n14690) );
  OAI21X1 U7004 ( .A0(n9812), .A1(n9854), .B0(n9811), .Y(n9824) );
  NOR2X1 U7005 ( .A(n14296), .B(n14298), .Y(n14217) );
  NOR2X1 U7006 ( .A(n12818), .B(n12802), .Y(n6028) );
  OAI21X1 U7007 ( .A0(n14361), .A1(n14358), .B0(n14362), .Y(n6496) );
  CMPR22X1 U7008 ( .A(U1_U1_y2[29]), .B(U1_U1_y0[29]), .CO(n12989), .S(n12986)
         );
  CMPR22X1 U7009 ( .A(U1_U1_y2[28]), .B(U1_U1_y0[28]), .CO(n12987), .S(n12984)
         );
  CMPR22X1 U7010 ( .A(U0_U0_y0[21]), .B(U0_U0_y1[21]), .CO(n13258), .S(n13255)
         );
  CMPR22X1 U7011 ( .A(U0_U0_y1[30]), .B(U0_U0_y0[30]), .CO(n13274), .S(n13271)
         );
  XNOR2X1 U7012 ( .A(U0_U0_y1[19]), .B(n7605), .Y(n13252) );
  NAND2X1 U7013 ( .A(n10260), .B(n6216), .Y(n6215) );
  CMPR22X1 U7014 ( .A(U1_U2_y1[28]), .B(U1_U2_y0[28]), .CO(n13005), .S(n13002)
         );
  CMPR22X1 U7015 ( .A(U1_U0_y1[22]), .B(U1_U0_y0[22]), .CO(n9309), .S(n9306)
         );
  CMPR22X1 U7016 ( .A(U1_U2_y1[30]), .B(U1_U2_y0[30]), .CO(n13050), .S(n13006)
         );
  CMPR22X1 U7017 ( .A(U1_U2_y1[27]), .B(U1_U2_y0[27]), .CO(n13003), .S(n13000)
         );
  CMPR22X1 U7018 ( .A(U0_U2_y2[32]), .B(U0_U2_y0[32]), .CO(n12218), .S(n12215)
         );
  AOI21XL U7019 ( .A0(n6147), .A1(n6146), .B0(n6169), .Y(n6145) );
  NAND2X2 U7020 ( .A(n7947), .B(W2[18]), .Y(n10340) );
  NAND2X2 U7021 ( .A(W0[20]), .B(W0[4]), .Y(n9842) );
  NAND2X1 U7022 ( .A(W0[7]), .B(W0[23]), .Y(n9832) );
  NAND2X1 U7023 ( .A(W1[4]), .B(W1[20]), .Y(n9989) );
  NAND2X1 U7024 ( .A(W1[6]), .B(W1[22]), .Y(n9983) );
  AND2X1 U7025 ( .A(U1_U1_y0[21]), .B(U1_U1_y2[21]), .Y(n6709) );
  NOR2X2 U7026 ( .A(n13850), .B(n13849), .Y(n13865) );
  NOR2X2 U7027 ( .A(n12186), .B(n12185), .Y(n12205) );
  NOR2BX2 U7028 ( .AN(n8403), .B(n6679), .Y(n8514) );
  NOR2X1 U7029 ( .A(n12699), .B(n12698), .Y(n12800) );
  XOR2X1 U7030 ( .A(U1_U1_y0[21]), .B(U1_U1_y2[21]), .Y(n12782) );
  NAND2X1 U7031 ( .A(n8418), .B(n8417), .Y(n8533) );
  NOR2X2 U7032 ( .A(n9982), .B(n9968), .Y(n7393) );
  XOR2X1 U7033 ( .A(U1_U1_y1[25]), .B(U1_U1_y0[25]), .Y(n14654) );
  NOR2X2 U7034 ( .A(n12160), .B(n6752), .Y(n12176) );
  NOR2X2 U7035 ( .A(n13808), .B(n13806), .Y(n6071) );
  NOR2X1 U7036 ( .A(n8743), .B(n8742), .Y(n8898) );
  CMPR22X1 U7037 ( .A(U1_U1_y1[27]), .B(U1_U1_y0[27]), .CO(n14661), .S(n14658)
         );
  CMPR22X1 U7038 ( .A(U1_U1_y1[28]), .B(U1_U1_y0[28]), .CO(n14663), .S(n14660)
         );
  CMPR22X1 U7039 ( .A(U0_U1_y1[30]), .B(U0_U1_y0[30]), .CO(n9064), .S(n9056)
         );
  CMPR22X1 U7040 ( .A(U1_U1_y1[30]), .B(U1_U1_y0[30]), .CO(n14667), .S(n14664)
         );
  CMPR22X1 U7041 ( .A(U1_U1_y1[29]), .B(U1_U1_y0[29]), .CO(n14665), .S(n14662)
         );
  CMPR22X1 U7042 ( .A(U0_U1_y1[26]), .B(U0_U1_y0[26]), .CO(n9051), .S(n8985)
         );
  CMPR22X1 U7043 ( .A(U0_U1_y1[27]), .B(U0_U1_y0[27]), .CO(n9053), .S(n9050)
         );
  OAI21X1 U7044 ( .A0(n6070), .A1(n6069), .B0(n6067), .Y(n6066) );
  CMPR22X1 U7045 ( .A(U1_U1_y1[23]), .B(U1_U1_y0[23]), .CO(n14653), .S(n14650)
         );
  CMPR22X1 U7046 ( .A(U1_U1_y1[24]), .B(U1_U1_y0[24]), .CO(n14655), .S(n14652)
         );
  NOR2XL U7047 ( .A(n10232), .B(n6217), .Y(n6216) );
  NAND2X2 U7048 ( .A(W1[18]), .B(W1[2]), .Y(n10007) );
  NAND2X2 U7049 ( .A(W2[18]), .B(W2[2]), .Y(n9946) );
  NAND2X1 U7050 ( .A(W1[9]), .B(W1[25]), .Y(n9964) );
  NOR2X2 U7051 ( .A(W1[20]), .B(W1[4]), .Y(n9972) );
  INVX2 U7052 ( .A(n6547), .Y(n7276) );
  INVX1 U7053 ( .A(U1_U0_y0[29]), .Y(n6670) );
  NOR2X2 U7054 ( .A(n13782), .B(n13781), .Y(n13808) );
  OAI21XL U7055 ( .A0(n8484), .A1(n8489), .B0(n8485), .Y(n6581) );
  NOR2X1 U7056 ( .A(n13779), .B(n13780), .Y(n13806) );
  CLKINVX3 U7057 ( .A(n6875), .Y(n6876) );
  NAND2BXL U7058 ( .AN(n13826), .B(n13822), .Y(n6070) );
  AOI2BB1X1 U7059 ( .A0N(n13826), .A1N(n13823), .B0(n6068), .Y(n6067) );
  XNOR2X1 U7060 ( .A(U0_U2_y1[16]), .B(n6355), .Y(n8740) );
  CMPR22X1 U7061 ( .A(U1_U0_y2[22]), .B(U1_U0_y0[22]), .CO(n8422), .S(n8419)
         );
  OAI21X1 U7062 ( .A0(n12094), .A1(n12098), .B0(n12095), .Y(n12066) );
  CMPR22X1 U7063 ( .A(U0_U0_y1[18]), .B(U0_U0_y0[18]), .CO(n13253), .S(n13250)
         );
  CMPR22X1 U7064 ( .A(U0_U2_y2[26]), .B(U0_U2_y0[26]), .CO(n12182), .S(n12161)
         );
  NOR2X2 U7065 ( .A(W1[2]), .B(W1[18]), .Y(n10006) );
  NAND2X2 U7066 ( .A(W1[19]), .B(W1[3]), .Y(n6547) );
  NOR2X2 U7067 ( .A(n10241), .B(n6736), .Y(n6735) );
  OAI21X2 U7068 ( .A0(n6736), .A1(n10240), .B0(n10194), .Y(n6734) );
  CMPR22X1 U7069 ( .A(U1_U2_y2[18]), .B(U1_U2_y0[18]), .CO(n13784), .S(n13781)
         );
  NOR2X2 U7070 ( .A(n7949), .B(W1[21]), .Y(n10196) );
  NOR2X2 U7071 ( .A(n7950), .B(W1[23]), .Y(n10198) );
  NAND2X1 U7072 ( .A(n8020), .B(W1[20]), .Y(n10257) );
  NAND2X2 U7073 ( .A(n8041), .B(W1[18]), .Y(n10240) );
  OR2X2 U7074 ( .A(W1[3]), .B(n7083), .Y(n10194) );
  NAND2X1 U7075 ( .A(n8038), .B(W1[22]), .Y(n10233) );
  NOR2X2 U7076 ( .A(n8041), .B(W1[18]), .Y(n10241) );
  NOR2X1 U7077 ( .A(n8020), .B(W1[20]), .Y(n10256) );
  CMPR22X1 U7078 ( .A(U0_U2_y2[19]), .B(U0_U2_y0[19]), .CO(n12071), .S(n12068)
         );
  CMPR22X1 U7079 ( .A(U0_U2_y2[18]), .B(U0_U2_y0[18]), .CO(n12069), .S(n12064)
         );
  NAND2X2 U7080 ( .A(n9717), .B(n7076), .Y(n17178) );
  XNOR2X2 U7081 ( .A(n9534), .B(n6956), .Y(n9717) );
  NOR2X2 U7082 ( .A(n12598), .B(n12597), .Y(n12623) );
  NOR2X1 U7083 ( .A(n6835), .B(n10045), .Y(n6406) );
  NAND3X2 U7084 ( .A(n11599), .B(n11593), .C(n11597), .Y(n7762) );
  AOI21X2 U7085 ( .A0(n10042), .A1(n6406), .B0(n10019), .Y(n10020) );
  OAI21X2 U7086 ( .A0(n22975), .A1(n22970), .B0(n22969), .Y(n6246) );
  NOR2X1 U7087 ( .A(n5847), .B(n24693), .Y(n22970) );
  CMPR22X1 U7088 ( .A(U1_U2_y2[39]), .B(U1_U2_y0[39]), .CO(n13992), .S(n13984)
         );
  OAI21X1 U7089 ( .A0(n22186), .A1(n22171), .B0(n22170), .Y(n22172) );
  CMPR22X1 U7090 ( .A(U0_U2_y2[15]), .B(U0_U2_y0[15]), .CO(n12061), .S(n12058)
         );
  NOR2X1 U7091 ( .A(n22187), .B(n22171), .Y(n22173) );
  AOI21X2 U7092 ( .A0(n6277), .A1(n9211), .B0(n9210), .Y(n7284) );
  NOR2X1 U7093 ( .A(n24993), .B(n24714), .Y(n9211) );
  NOR2X1 U7094 ( .A(n12404), .B(n22968), .Y(n14581) );
  NOR2X1 U7095 ( .A(n6145), .B(n12693), .Y(n7827) );
  CMPR22X1 U7096 ( .A(U1_U2_y1[23]), .B(U1_U2_y0[23]), .CO(n12911), .S(n12907)
         );
  NAND2X2 U7097 ( .A(n9744), .B(n9743), .Y(n10067) );
  XOR2X1 U7098 ( .A(n9114), .B(n9104), .Y(n24652) );
  NAND2X1 U7099 ( .A(n9103), .B(n9112), .Y(n9104) );
  NOR2X1 U7100 ( .A(n8191), .B(BOPC[36]), .Y(n11146) );
  NOR2X1 U7101 ( .A(n7997), .B(W2[27]), .Y(n10272) );
  AOI21XL U7102 ( .A0(n8220), .A1(n10426), .B0(n8219), .Y(n8221) );
  NOR2X2 U7103 ( .A(n8081), .B(AOPB[29]), .Y(n10502) );
  NOR2X2 U7104 ( .A(n8135), .B(BOPB[29]), .Y(n10665) );
  NOR2X2 U7105 ( .A(W2[11]), .B(W2[27]), .Y(n9886) );
  NAND2X2 U7106 ( .A(n8226), .B(n10397), .Y(n6428) );
  NOR2X2 U7107 ( .A(W2[25]), .B(W2[9]), .Y(n9892) );
  NAND2X1 U7108 ( .A(W2[4]), .B(W2[20]), .Y(n9911) );
  NAND2X2 U7109 ( .A(W2[19]), .B(W2[3]), .Y(n9916) );
  NOR2X1 U7110 ( .A(n8050), .B(W1[25]), .Y(n10200) );
  OAI2BB1X2 U7111 ( .A0N(n9867), .A1N(n9866), .B0(n9865), .Y(n6335) );
  NOR2X1 U7112 ( .A(n12942), .B(n12943), .Y(n12978) );
  INVX1 U7113 ( .A(n7868), .Y(n6050) );
  AOI21XL U7114 ( .A0(n10519), .A1(n10518), .B0(n10517), .Y(n10520) );
  AOI21XL U7115 ( .A0(n10397), .A1(n10401), .B0(n10388), .Y(n10389) );
  OAI21XL U7116 ( .A0(n10477), .A1(n10464), .B0(n10463), .Y(n10468) );
  AOI21XL U7117 ( .A0(n10373), .A1(n10384), .B0(n10372), .Y(n10374) );
  NAND2X1 U7118 ( .A(n11536), .B(n11540), .Y(n11526) );
  AOI21XL U7119 ( .A0(n10839), .A1(n10819), .B0(n10818), .Y(n10829) );
  AND2X1 U7120 ( .A(n10792), .B(n10791), .Y(n6965) );
  NAND2X1 U7121 ( .A(n6223), .B(n6221), .Y(n11072) );
  XNOR2X1 U7122 ( .A(n10944), .B(n10943), .Y(U0_U2_z0[15]) );
  INVX1 U7123 ( .A(n6205), .Y(n11416) );
  NOR2X1 U7124 ( .A(n8030), .B(W3[20]), .Y(n10058) );
  NOR2X2 U7125 ( .A(n8040), .B(W1[17]), .Y(n6737) );
  AND2X1 U7126 ( .A(n24666), .B(n24640), .Y(n8034) );
  CMPR22X1 U7127 ( .A(U0_U0_y2[24]), .B(U0_U0_y0[24]), .CO(n14232), .S(n14229)
         );
  INVX1 U7128 ( .A(n13153), .Y(n6790) );
  CMPR22X1 U7129 ( .A(U0_U1_y1[21]), .B(U0_U1_y0[21]), .CO(n8933), .S(n8835)
         );
  AND2X1 U7130 ( .A(U1_U2_y2[23]), .B(U1_U2_y0[23]), .Y(n13857) );
  AOI21XL U7131 ( .A0(n8384), .A1(n8383), .B0(n8382), .Y(n8493) );
  OAI21X1 U7132 ( .A0(n13865), .A1(n13862), .B0(n13866), .Y(n6034) );
  CMPR22X1 U7133 ( .A(U1_U1_y2[23]), .B(U1_U1_y0[23]), .CO(n12898), .S(n12894)
         );
  CLKINVX2 U7134 ( .A(n9479), .Y(n5870) );
  CMPR22X1 U7135 ( .A(U1_U1_y1[26]), .B(U1_U1_y0[26]), .CO(n14659), .S(n14656)
         );
  AND2X1 U7136 ( .A(U1_U1_y1[31]), .B(U1_U1_y0[31]), .Y(n14669) );
  INVX1 U7137 ( .A(U2_B_i[23]), .Y(n11453) );
  AOI21XL U7138 ( .A0(n11599), .A1(n11597), .B0(n11591), .Y(n11595) );
  AND2X1 U7139 ( .A(n11077), .B(n11076), .Y(n11078) );
  AOI21XL U7140 ( .A0(n11253), .A1(n11243), .B0(n11242), .Y(n11244) );
  XOR2X1 U7141 ( .A(n6225), .B(BOPA[40]), .Y(n6224) );
  AND2X1 U7142 ( .A(n24662), .B(n24642), .Y(n8032) );
  OAI21X2 U7143 ( .A0(n14434), .A1(n14439), .B0(n14435), .Y(n14423) );
  NOR2X1 U7144 ( .A(n13252), .B(n13253), .Y(n13308) );
  OAI21X1 U7145 ( .A0(n12562), .A1(n12561), .B0(n12560), .Y(n12587) );
  OAI21X2 U7146 ( .A0(n13304), .A1(n13309), .B0(n13305), .Y(n13313) );
  OAI21X1 U7147 ( .A0(n12195), .A1(n12200), .B0(n12196), .Y(n12211) );
  AND2X1 U7148 ( .A(n19761), .B(U1_A_r_d0[16]), .Y(n19762) );
  NOR2X1 U7149 ( .A(n5934), .B(n13897), .Y(n13913) );
  NAND2X2 U7150 ( .A(n13589), .B(n7830), .Y(n7786) );
  NAND2X1 U7151 ( .A(n9316), .B(n9317), .Y(n9477) );
  AOI21XL U7152 ( .A0(n8399), .A1(n8398), .B0(n6691), .Y(n8499) );
  NOR2X1 U7153 ( .A(n6070), .B(n6065), .Y(n6064) );
  INVX1 U7154 ( .A(n9437), .Y(n7614) );
  XOR2XL U7155 ( .A(n10511), .B(n10510), .Y(U0_U0_z0[2]) );
  OAI21X1 U7156 ( .A0(n6712), .A1(n9567), .B0(n9566), .Y(n9569) );
  AND2X1 U7157 ( .A(n10892), .B(n10891), .Y(n6962) );
  XOR2XL U7158 ( .A(n11395), .B(n11394), .Y(U0_U1_z0[2]) );
  OAI21XL U7159 ( .A0(n28683), .A1(n11428), .B0(n11409), .Y(U2_B_r[14]) );
  CLKINVX2 U7160 ( .A(n8044), .Y(n29098) );
  NAND3X2 U7161 ( .A(n7161), .B(n7803), .C(n7887), .Y(n6010) );
  AND2X1 U7162 ( .A(n9537), .B(U1_A_i_d0[23]), .Y(n9538) );
  CMPR22X1 U7163 ( .A(U2_U0_y1[19]), .B(U2_U0_y0[19]), .CO(n26080), .S(n26036)
         );
  CMPR22X1 U7164 ( .A(U2_U0_y2[28]), .B(U2_U0_y0[28]), .CO(n23936), .S(n23871)
         );
  INVX1 U7165 ( .A(n26867), .Y(n21530) );
  INVX1 U7166 ( .A(n24207), .Y(n18818) );
  OAI21XL U7167 ( .A0(n22160), .A1(n22202), .B0(n22159), .Y(n22161) );
  NOR2X1 U7168 ( .A(n24669), .B(n24732), .Y(n24671) );
  INVX1 U7169 ( .A(n21949), .Y(n6758) );
  AOI21XL U7170 ( .A0(n12082), .A1(n12133), .B0(n12138), .Y(n12150) );
  INVX1 U7171 ( .A(n12139), .Y(n12122) );
  XOR2XL U7172 ( .A(U0_U2_y0[40]), .B(U0_U2_y2[40]), .Y(n12359) );
  AND2X1 U7173 ( .A(n9110), .B(n9109), .Y(n9111) );
  AOI21XL U7174 ( .A0(n8794), .A1(n8793), .B0(n8792), .Y(n8880) );
  AND2X1 U7175 ( .A(n13858), .B(n13870), .Y(n13859) );
  AND2X1 U7176 ( .A(n9341), .B(n9533), .Y(n6956) );
  AOI21XL U7177 ( .A0(n7005), .A1(n14885), .B0(n14884), .Y(n14886) );
  AND2X1 U7178 ( .A(n13877), .B(n13892), .Y(n6920) );
  AND2X1 U7179 ( .A(n13068), .B(n13079), .Y(n6894) );
  XOR2XL U7180 ( .A(n13977), .B(n7011), .Y(n14961) );
  AND2X1 U7181 ( .A(n13911), .B(n13910), .Y(n6905) );
  AND2X1 U7182 ( .A(n13085), .B(n13580), .Y(n6927) );
  OAI21XL U7183 ( .A0(n14837), .A1(n19256), .B0(n14836), .Y(n14838) );
  AOI21XL U7184 ( .A0(n13796), .A1(n13847), .B0(n7469), .Y(n13864) );
  AND2X1 U7185 ( .A(n14694), .B(n14693), .Y(n6930) );
  AND2X1 U7186 ( .A(n14845), .B(n14844), .Y(n7189) );
  XNOR2X2 U7187 ( .A(n10708), .B(n10707), .Y(U1_U2_z0[24]) );
  BUFX1 U7188 ( .A(U2_B_r[8]), .Y(n7130) );
  XOR2XL U7189 ( .A(U0_U2_y0[40]), .B(U0_U2_y1[40]), .Y(n12352) );
  ADDHXL U7190 ( .A(U0_pipe7[17]), .B(U0_pipe6[17]), .CO(n23955), .S(n23900)
         );
  ADDFX2 U7191 ( .A(n18408), .B(n18407), .CI(U2_A_i_d[13]), .CO(n18409), .S(
        n18363) );
  AND2X1 U7192 ( .A(n5872), .B(n5873), .Y(n6259) );
  OAI21XL U7193 ( .A0(n25049), .A1(n9010), .B0(n9009), .Y(n9011) );
  NOR2X1 U7194 ( .A(n22913), .B(n13114), .Y(n22044) );
  XOR2XL U7195 ( .A(n14302), .B(n14301), .Y(n25263) );
  XOR2X2 U7196 ( .A(n7306), .B(n13448), .Y(n14099) );
  XOR2X1 U7197 ( .A(n9196), .B(n7253), .Y(n24675) );
  XOR2X1 U7198 ( .A(n6768), .B(n12097), .Y(n13103) );
  XOR2X2 U7199 ( .A(n6275), .B(n6969), .Y(n24654) );
  XNOR2X1 U7200 ( .A(n12558), .B(n12557), .Y(n22915) );
  XOR2XL U7201 ( .A(n8904), .B(n8903), .Y(n24602) );
  NOR2X1 U7202 ( .A(n7233), .B(n7232), .Y(n14073) );
  XOR2XL U7203 ( .A(n12346), .B(n12345), .Y(n12347) );
  XOR2X1 U7204 ( .A(n9130), .B(n9129), .Y(n24647) );
  XNOR2XL U7205 ( .A(n8924), .B(n8923), .Y(n24587) );
  AOI21XL U7206 ( .A0(n19755), .A1(n19862), .B0(n19759), .Y(n19848) );
  INVX1 U7207 ( .A(n19974), .Y(n14934) );
  OAI21XL U7208 ( .A0(n17622), .A1(n14509), .B0(n14508), .Y(n17610) );
  XOR2X1 U7209 ( .A(n6689), .B(n8539), .Y(n19737) );
  XOR2X1 U7210 ( .A(n8552), .B(n8551), .Y(n19744) );
  XOR2X1 U7211 ( .A(n6584), .B(n8467), .Y(n19724) );
  OAI21XL U7212 ( .A0(n20254), .A1(n12307), .B0(n12306), .Y(n12308) );
  XOR2XL U7213 ( .A(n9403), .B(n9395), .Y(n13667) );
  XOR2XL U7214 ( .A(n8535), .B(n8477), .Y(n12296) );
  XOR2XL U7215 ( .A(n13812), .B(n13811), .Y(n19951) );
  XOR2XL U7216 ( .A(n7713), .B(n9356), .Y(n13675) );
  XOR2X2 U7217 ( .A(n9443), .B(n9442), .Y(n9681) );
  XOR2XL U7218 ( .A(n12817), .B(n12816), .Y(n19358) );
  XNOR2XL U7219 ( .A(n13048), .B(n12918), .Y(n19326) );
  XOR2XL U7220 ( .A(n7420), .B(n14782), .Y(n19984) );
  NAND2X1 U7221 ( .A(n6110), .B(n6109), .Y(n19594) );
  XOR2XL U7222 ( .A(n12352), .B(n12351), .Y(n12353) );
  OAI21X1 U7223 ( .A0(n21946), .A1(n7729), .B0(n6805), .Y(n7730) );
  XNOR2X1 U7224 ( .A(n9349), .B(n5791), .Y(n14974) );
  AOI21XL U7225 ( .A0(n23274), .A1(n23273), .B0(n23272), .Y(n23480) );
  OAI21XL U7226 ( .A0(n23689), .A1(n23924), .B0(n23932), .Y(n23741) );
  AOI21XL U7227 ( .A0(n25093), .A1(n8926), .B0(n8925), .Y(n25072) );
  AOI21XL U7228 ( .A0(n24509), .A1(n24922), .B0(n13511), .Y(n13512) );
  AND2X1 U7229 ( .A(n14088), .B(U2_A_r_d[13]), .Y(n24492) );
  AOI21XL U7230 ( .A0(n25517), .A1(n25516), .B0(n25515), .Y(n25537) );
  NOR2X1 U7231 ( .A(n21954), .B(n6447), .Y(n6446) );
  AOI21XL U7232 ( .A0(n21823), .A1(n21799), .B0(n21798), .Y(n21816) );
  AND2X1 U7233 ( .A(n5863), .B(U2_A_i_d[17]), .Y(n21852) );
  XOR2XL U7234 ( .A(n14321), .B(n14320), .Y(n25458) );
  AOI21XL U7235 ( .A0(n23049), .A1(n23001), .B0(n23000), .Y(n23014) );
  OAI21XL U7236 ( .A0(n13498), .A1(n13494), .B0(n13495), .Y(n13300) );
  AOI21XL U7237 ( .A0(n14083), .A1(n22810), .B0(n14082), .Y(n14084) );
  OAI21XL U7238 ( .A0(n25755), .A1(n12132), .B0(n12131), .Y(n6762) );
  XOR2XL U7239 ( .A(n13346), .B(n13345), .Y(n14016) );
  AND2X1 U7240 ( .A(n14441), .B(U2_A_r_d[13]), .Y(n25197) );
  AOI21XL U7241 ( .A0(n19766), .A1(n19836), .B0(n7039), .Y(n19824) );
  INVX1 U7242 ( .A(n19790), .Y(n5851) );
  AOI21XL U7243 ( .A0(n14877), .A1(n14876), .B0(n14875), .Y(n20389) );
  NOR2X1 U7244 ( .A(n20341), .B(n20327), .Y(n7842) );
  AOI21XL U7245 ( .A0(n9455), .A1(n9454), .B0(n9453), .Y(n17527) );
  AND2X1 U7246 ( .A(n9690), .B(U1_A_i_d0[13]), .Y(n17516) );
  AND2X1 U7247 ( .A(n19744), .B(U1_A_r_d0[11]), .Y(n19875) );
  AND2X1 U7248 ( .A(n19765), .B(U1_A_i_d0[17]), .Y(n6675) );
  AOI21XL U7249 ( .A0(n14920), .A1(n16909), .B0(n14919), .Y(n16889) );
  AOI21XL U7250 ( .A0(n9679), .A1(n9678), .B0(n9677), .Y(n19153) );
  AND2X1 U7251 ( .A(n9700), .B(U1_A_r_d0[17]), .Y(n19117) );
  OAI21XL U7252 ( .A0(n19393), .A1(n19085), .B0(n19086), .Y(n13714) );
  AOI21XL U7253 ( .A0(n24701), .A1(n5849), .B0(n6776), .Y(n6775) );
  OAI21XL U7254 ( .A0(n19254), .A1(n19242), .B0(n19241), .Y(n19246) );
  AOI21XL U7255 ( .A0(n24740), .A1(n24739), .B0(n24733), .Y(n24736) );
  INVX1 U7256 ( .A(n17455), .Y(n17476) );
  OAI21XL U7257 ( .A0(n17476), .A1(n17464), .B0(n17463), .Y(n17467) );
  AOI21X1 U7258 ( .A0(n17455), .A1(n7412), .B0(n7411), .Y(n17454) );
  OR2X2 U7259 ( .A(n28672), .B(n28678), .Y(n15967) );
  XOR2XL U7260 ( .A(n21693), .B(n21692), .Y(n7416) );
  OAI21XL U7261 ( .A0(n24742), .A1(n24732), .B0(n24731), .Y(n24740) );
  AOI21XL U7262 ( .A0(n24501), .A1(n24480), .B0(n24479), .Y(n24490) );
  INVX1 U7263 ( .A(n21952), .Y(n21976) );
  AOI21XL U7264 ( .A0(n22022), .A1(n22003), .B0(n22002), .Y(n22012) );
  XOR2XL U7265 ( .A(n12506), .B(n12505), .Y(n22727) );
  OAI21XL U7266 ( .A0(n21813), .A1(n21807), .B0(n21806), .Y(n21810) );
  CLKINVX2 U7267 ( .A(n6795), .Y(n22997) );
  NAND2BX2 U7268 ( .AN(n12579), .B(n6377), .Y(n22655) );
  XOR2XL U7269 ( .A(n8888), .B(n8887), .Y(n25448) );
  AOI21XL U7270 ( .A0(n25205), .A1(n25185), .B0(n25184), .Y(n25195) );
  NAND2BX1 U7271 ( .AN(n19991), .B(n5944), .Y(n20101) );
  AOI21XL U7272 ( .A0(n17347), .A1(n17327), .B0(n17326), .Y(n5955) );
  NAND2X1 U7273 ( .A(n7445), .B(n6054), .Y(n20361) );
  AOI21XL U7274 ( .A0(n17524), .A1(n17505), .B0(n17504), .Y(n17514) );
  AOI21XL U7275 ( .A0(n17664), .A1(n14500), .B0(n14505), .Y(n17632) );
  XOR2XL U7276 ( .A(n19568), .B(n14976), .Y(n7931) );
  OAI2BB1X1 U7277 ( .A0N(n14007), .A1N(n5966), .B0(n7821), .Y(n17081) );
  AOI21XL U7278 ( .A0(n16666), .A1(n16660), .B0(n16659), .Y(n16663) );
  OAI21XL U7279 ( .A0(n19116), .A1(n19105), .B0(n19104), .Y(n19114) );
  AOI21XL U7280 ( .A0(n16993), .A1(n16958), .B0(n16957), .Y(n16969) );
  XOR2XL U7281 ( .A(n12840), .B(n12839), .Y(n16932) );
  AOI21XL U7282 ( .A0(n7685), .A1(n19434), .B0(n19433), .Y(n19441) );
  BUFX4 U7283 ( .A(n5826), .Y(n27162) );
  BUFX4 U7284 ( .A(n5921), .Y(n28143) );
  CLKINVX3 U7285 ( .A(n27386), .Y(n5904) );
  AOI21XL U7286 ( .A0(n7166), .A1(n7000), .B0(n7164), .Y(n7163) );
  XNOR2XL U7287 ( .A(n19265), .B(n19264), .Y(n19266) );
  NOR2X1 U7288 ( .A(cs[1]), .B(cs[2]), .Y(n11636) );
  AOI21XL U7289 ( .A0(n6635), .A1(n6610), .B0(n6609), .Y(n8640) );
  XOR2XL U7290 ( .A(n25341), .B(n25340), .Y(n25342) );
  XOR2XL U7291 ( .A(n7733), .B(n7732), .Y(n12407) );
  XOR2XL U7292 ( .A(n17459), .B(n7616), .Y(n17460) );
  XNOR2XL U7293 ( .A(n26818), .B(n26610), .Y(n26611) );
  XNOR2XL U7294 ( .A(n23632), .B(n23580), .Y(n23581) );
  XOR2XL U7295 ( .A(n24103), .B(n24102), .Y(n24104) );
  XNOR2XL U7296 ( .A(n20818), .B(n20817), .Y(n20819) );
  XNOR2XL U7297 ( .A(n21614), .B(n21578), .Y(n21579) );
  XOR2XL U7298 ( .A(n18194), .B(n18193), .Y(n18195) );
  XNOR2XL U7299 ( .A(n24894), .B(n24893), .Y(n24895) );
  AOI21XL U7300 ( .A0(n6859), .A1(n7763), .B0(n6858), .Y(n24695) );
  XNOR2XL U7301 ( .A(n24788), .B(n24787), .Y(n24789) );
  XNOR2XL U7302 ( .A(n24437), .B(n24436), .Y(n24438) );
  AOI21XL U7303 ( .A0(n6528), .A1(n6527), .B0(n6526), .Y(n6525) );
  XOR2XL U7304 ( .A(n25534), .B(n25533), .Y(n25535) );
  XNOR2XL U7305 ( .A(n25614), .B(n25613), .Y(n25615) );
  XOR2XL U7306 ( .A(n21976), .B(n21975), .Y(n21977) );
  XOR2XL U7307 ( .A(n21837), .B(n21836), .Y(n21838) );
  XNOR2XL U7308 ( .A(n22344), .B(n22343), .Y(n22345) );
  XNOR2XL U7309 ( .A(n23012), .B(n23011), .Y(n23013) );
  XOR2XL U7310 ( .A(n22795), .B(n22794), .Y(n22796) );
  AOI2BB1X1 U7311 ( .A0N(n25658), .A1N(n25656), .B0(n6457), .Y(n25655) );
  XNOR2XL U7312 ( .A(n25735), .B(n25734), .Y(n25736) );
  XOR2XL U7313 ( .A(n22597), .B(n22979), .Y(n22598) );
  XOR2XL U7314 ( .A(n25366), .B(n25365), .Y(n25367) );
  XOR2XL U7315 ( .A(n20097), .B(n20096), .Y(n20098) );
  XOR2XL U7316 ( .A(n17392), .B(n17391), .Y(n17393) );
  XOR2XL U7317 ( .A(n20395), .B(n20394), .Y(n20396) );
  XNOR2XL U7318 ( .A(n17551), .B(n17550), .Y(n17552) );
  XNOR2XL U7319 ( .A(n17510), .B(n17509), .Y(n17511) );
  XNOR2XL U7320 ( .A(n17693), .B(n17692), .Y(n17694) );
  XNOR2XL U7321 ( .A(n19884), .B(n19883), .Y(n19885) );
  XNOR2XL U7322 ( .A(n17061), .B(n17060), .Y(n17062) );
  XNOR2XL U7323 ( .A(n16730), .B(n16729), .Y(n16731) );
  XNOR2XL U7324 ( .A(n16638), .B(n16637), .Y(n16639) );
  XOR2XL U7325 ( .A(n16863), .B(n16862), .Y(n16864) );
  XNOR2XL U7326 ( .A(n19180), .B(n19179), .Y(n19181) );
  XNOR2XL U7327 ( .A(n19361), .B(n19360), .Y(n19362) );
  XOR2XL U7328 ( .A(n6586), .B(n16965), .Y(n16966) );
  XOR2XL U7329 ( .A(n19420), .B(n19419), .Y(n19421) );
  XOR2XL U7330 ( .A(n19645), .B(n19644), .Y(n19646) );
  XOR2XL U7331 ( .A(n19591), .B(n19590), .Y(n19592) );
  AND2X1 U7332 ( .A(cs[0]), .B(cs[1]), .Y(n7305) );
  CLKINVX3 U7333 ( .A(n27496), .Y(n27686) );
  BUFX4 U7334 ( .A(n27379), .Y(n28068) );
  BUFX4 U7335 ( .A(n27431), .Y(n28179) );
  AOI21XL U7336 ( .A0(n27976), .A1(Q1[9]), .B0(n27852), .Y(n28352) );
  AOI21XL U7337 ( .A0(n27976), .A1(Q1[31]), .B0(n27947), .Y(n28483) );
  BUFX4 U7338 ( .A(n27772), .Y(n28295) );
  AND2X1 U7339 ( .A(n5693), .B(n5694), .Y(n29242) );
  BUFX3 U7340 ( .A(n11620), .Y(n29094) );
  BUFX3 U7341 ( .A(n11617), .Y(n29109) );
  AND2X1 U7342 ( .A(n9883), .B(n9882), .Y(n5759) );
  BUFX3 U7343 ( .A(n28322), .Y(n27631) );
  INVX1 U7344 ( .A(n28322), .Y(n11940) );
  OR2X2 U7345 ( .A(n7976), .B(W1[15]), .Y(n5761) );
  AND2X2 U7346 ( .A(n5761), .B(n10255), .Y(n5762) );
  AND2X1 U7347 ( .A(n9828), .B(n9827), .Y(n5763) );
  AND2X1 U7348 ( .A(U1_U0_y1[25]), .B(U1_U0_y0[25]), .Y(n5764) );
  INVX1 U7349 ( .A(n19758), .Y(n19754) );
  XOR2X1 U7350 ( .A(n6655), .B(n8579), .Y(n19758) );
  OR2X2 U7351 ( .A(n21532), .B(n21531), .Y(n5765) );
  XOR2X4 U7352 ( .A(n10263), .B(n10262), .Y(n5766) );
  OR2X2 U7353 ( .A(n14515), .B(n22892), .Y(n5767) );
  OR2X2 U7354 ( .A(n22892), .B(n13099), .Y(n5768) );
  AND2X1 U7355 ( .A(n9888), .B(n9887), .Y(n5769) );
  BUFX3 U7356 ( .A(W1[3]), .Y(n7143) );
  CLKINVX3 U7357 ( .A(n28054), .Y(n27205) );
  XNOR2X2 U7358 ( .A(n10073), .B(n6401), .Y(U2_U0_z2[3]) );
  AND2X2 U7359 ( .A(n9967), .B(n7393), .Y(n5770) );
  NOR2X2 U7360 ( .A(n8038), .B(W1[22]), .Y(n10232) );
  XOR2X4 U7361 ( .A(n9895), .B(n10307), .Y(n5771) );
  AND2X1 U7362 ( .A(n9726), .B(n9957), .Y(n5772) );
  BUFX3 U7363 ( .A(n5927), .Y(n7123) );
  CLKINVX2 U7364 ( .A(n11953), .Y(n11952) );
  CLKINVX2 U7365 ( .A(n11953), .Y(n11958) );
  BUFX3 U7366 ( .A(n5834), .Y(n11956) );
  INVX12 U7367 ( .A(n28997), .Y(n23239) );
  INVX12 U7368 ( .A(n28997), .Y(n24128) );
  CLKBUFX8 U7369 ( .A(OP2_done0), .Y(n27976) );
  CLKINVX3 U7370 ( .A(R7_valid), .Y(n5807) );
  CLKINVX2 U7371 ( .A(n5924), .Y(n6885) );
  CLKINVX2 U7372 ( .A(n5924), .Y(n6883) );
  CLKINVX2 U7373 ( .A(n5924), .Y(n6884) );
  CLKBUFX8 U7374 ( .A(n16496), .Y(n5924) );
  CLKINVX3 U7375 ( .A(R7_valid), .Y(n16496) );
  OR2X2 U7376 ( .A(n25125), .B(U2_A_r_d[25]), .Y(n5774) );
  OR2X2 U7377 ( .A(n25216), .B(U2_A_r_d[11]), .Y(n5775) );
  OR2X2 U7378 ( .A(n14018), .B(U2_A_r_d[1]), .Y(n5778) );
  OR2X2 U7379 ( .A(U0_U1_y1[11]), .B(U0_U1_y0[11]), .Y(n5779) );
  CLKINVX2 U7380 ( .A(n24696), .Y(n5815) );
  XOR2XL U7381 ( .A(n6436), .B(n12347), .Y(n24696) );
  INVX1 U7382 ( .A(U2_B_i[1]), .Y(n8308) );
  XNOR2XL U7383 ( .A(U2_U0_y2[39]), .B(U2_U0_y0[39]), .Y(n5784) );
  XNOR2XL U7384 ( .A(U2_U0_y1[39]), .B(U2_U0_y0[39]), .Y(n5785) );
  OR2X2 U7385 ( .A(n19758), .B(U1_A_i_d0[14]), .Y(n5786) );
  OR2X2 U7386 ( .A(n19986), .B(n19532), .Y(n5788) );
  XNOR2XL U7387 ( .A(n13993), .B(n13992), .Y(n5789) );
  INVX1 U7388 ( .A(n7814), .Y(n20026) );
  XOR2X2 U7389 ( .A(n5989), .B(n5789), .Y(n7814) );
  NAND2X1 U7390 ( .A(n14803), .B(n14802), .Y(n5790) );
  INVX1 U7391 ( .A(n16796), .Y(n5844) );
  XNOR2XL U7392 ( .A(n9348), .B(n9347), .Y(n5791) );
  AND2X1 U7393 ( .A(n8446), .B(n8588), .Y(n5792) );
  OR2X2 U7394 ( .A(n9029), .B(n9030), .Y(n5793) );
  OR2X2 U7395 ( .A(n24661), .B(n24660), .Y(n5794) );
  CLKINVX2 U7396 ( .A(n22884), .Y(n5814) );
  AND2X1 U7397 ( .A(n6796), .B(n22591), .Y(n5795) );
  OR2X2 U7398 ( .A(n14053), .B(U2_A_i_d[20]), .Y(n5796) );
  INVX1 U7399 ( .A(n9829), .Y(n9844) );
  AOI2BB1X2 U7400 ( .A0N(n9829), .A1N(n7556), .B0(n9830), .Y(n9836) );
  MXI2XL U7401 ( .A(n7511), .B(U1_pipe5[26]), .S0(n8053), .Y(n4923) );
  XNOR2X1 U7402 ( .A(n22312), .B(n22311), .Y(n22313) );
  MXI2X1 U7403 ( .A(n6003), .B(U1_pipe5[27]), .S0(n6002), .Y(n4924) );
  MXI2XL U7404 ( .A(n6613), .B(U1_pipe4[25]), .S0(n5835), .Y(n5093) );
  NAND3X1 U7405 ( .A(n7648), .B(n7625), .C(n7624), .Y(n9733) );
  MXI2X1 U7406 ( .A(n6300), .B(U0_pipe1[27]), .S0(n5835), .Y(n4404) );
  XNOR2X1 U7407 ( .A(n19401), .B(n19400), .Y(n19402) );
  XOR2X1 U7408 ( .A(n6082), .B(n20338), .Y(n6081) );
  MXI2XL U7409 ( .A(n7338), .B(U1_pipe9[25]), .S0(n5837), .Y(n4835) );
  AOI21XL U7410 ( .A0(n7503), .A1(n7178), .B0(n7212), .Y(n7505) );
  NAND2X1 U7411 ( .A(n6119), .B(n20039), .Y(n6118) );
  NAND2XL U7412 ( .A(n7487), .B(n7482), .Y(n7481) );
  MXI2XL U7413 ( .A(n7418), .B(U0_pipe15[25]), .S0(n5837), .Y(n4611) );
  INVXL U7414 ( .A(n7487), .Y(n6681) );
  NAND2XL U7415 ( .A(n6001), .B(n13994), .Y(n13995) );
  XOR2X1 U7416 ( .A(n5984), .B(n19575), .Y(n19576) );
  XOR2X1 U7417 ( .A(n16806), .B(n16805), .Y(n16807) );
  AOI21X1 U7418 ( .A0(n7178), .A1(n17297), .B0(n13651), .Y(n14109) );
  XOR2X1 U7419 ( .A(n5973), .B(n16803), .Y(n5972) );
  XOR2X1 U7420 ( .A(n16828), .B(n16827), .Y(n16829) );
  XNOR2X1 U7421 ( .A(n17090), .B(n17089), .Y(n17091) );
  MXI2XL U7422 ( .A(n7809), .B(U1_pipe3[25]), .S0(n5928), .Y(n5065) );
  AOI21X1 U7423 ( .A0(n7470), .A1(n7838), .B0(n5943), .Y(n5942) );
  NAND2XL U7424 ( .A(n6114), .B(n7855), .Y(n6113) );
  INVXL U7425 ( .A(n25526), .Y(n25527) );
  XOR2X1 U7426 ( .A(n16652), .B(n16651), .Y(n16653) );
  INVX1 U7427 ( .A(n7470), .Y(n16806) );
  MXI2X1 U7428 ( .A(U0_pipe10[21]), .B(n22768), .S0(n7095), .Y(n4556) );
  INVXL U7429 ( .A(n25656), .Y(n6458) );
  NAND2XL U7430 ( .A(n7491), .B(n20337), .Y(n7476) );
  AOI21X1 U7431 ( .A0(n7470), .A1(n7472), .B0(n7471), .Y(n5973) );
  XNOR2X1 U7432 ( .A(n16832), .B(n16831), .Y(n16833) );
  AOI21XL U7433 ( .A0(n21952), .A1(n6203), .B0(n6202), .Y(n6201) );
  XNOR2X1 U7434 ( .A(n25345), .B(n25344), .Y(n25346) );
  AOI21X1 U7435 ( .A0(n17455), .A1(n7618), .B0(n7617), .Y(n7616) );
  XOR2X1 U7436 ( .A(n19121), .B(n19120), .Y(n19122) );
  XNOR2X1 U7437 ( .A(n16821), .B(n16820), .Y(n16822) );
  XNOR2X1 U7438 ( .A(n17476), .B(n17475), .Y(n6914) );
  INVX1 U7439 ( .A(n20338), .Y(n6058) );
  INVXL U7440 ( .A(n12406), .Y(n6305) );
  XNOR2X1 U7441 ( .A(n23024), .B(n23023), .Y(n23025) );
  XNOR2X1 U7442 ( .A(n19125), .B(n19124), .Y(n19126) );
  INVXL U7443 ( .A(n17060), .Y(n16798) );
  INVX1 U7444 ( .A(n16823), .Y(n16832) );
  XNOR2X1 U7445 ( .A(n23034), .B(n23033), .Y(n23035) );
  AOI21XL U7446 ( .A0(n16633), .A1(n6518), .B0(n6602), .Y(n16631) );
  XOR2X1 U7447 ( .A(n21855), .B(n21854), .Y(n21856) );
  XNOR2X1 U7448 ( .A(n22640), .B(n22639), .Y(n22641) );
  XOR2X1 U7449 ( .A(n17101), .B(n17100), .Y(n17102) );
  XNOR2X1 U7450 ( .A(n20077), .B(n20076), .Y(n20078) );
  INVX1 U7451 ( .A(n6457), .Y(n25657) );
  XNOR2X1 U7452 ( .A(n22626), .B(n22625), .Y(n22627) );
  XOR2X1 U7453 ( .A(n25016), .B(n25015), .Y(n25017) );
  NAND2XL U7454 ( .A(n7219), .B(n20329), .Y(n6060) );
  XOR2X1 U7455 ( .A(n22619), .B(n22618), .Y(n22621) );
  INVX1 U7456 ( .A(n7491), .Y(n5986) );
  INVX1 U7457 ( .A(n6384), .Y(n6383) );
  INVXL U7458 ( .A(n12402), .Y(n6304) );
  XNOR2X1 U7459 ( .A(n22007), .B(n22006), .Y(n22008) );
  XNOR2X1 U7460 ( .A(n21988), .B(n21987), .Y(n21989) );
  NAND3X1 U7461 ( .A(n5964), .B(n5962), .C(n5961), .Y(n6156) );
  CLKINVX2 U7462 ( .A(n16944), .Y(n7535) );
  OAI21XL U7463 ( .A0(n25036), .A1(n25031), .B0(n25033), .Y(n6363) );
  NAND2XL U7464 ( .A(n6350), .B(n25018), .Y(n6349) );
  XOR2X1 U7465 ( .A(n17496), .B(n17495), .Y(n17497) );
  XOR2X1 U7466 ( .A(n7598), .B(n7597), .Y(n25529) );
  XOR2X1 U7467 ( .A(n17095), .B(n17094), .Y(n17096) );
  XNOR2X1 U7468 ( .A(n19114), .B(n19113), .Y(n19115) );
  XNOR2X1 U7469 ( .A(n25707), .B(n25706), .Y(n25708) );
  XNOR2X1 U7470 ( .A(n24750), .B(n24749), .Y(n24751) );
  XOR2X1 U7471 ( .A(n16663), .B(n16662), .Y(n16664) );
  INVXL U7472 ( .A(n7857), .Y(n6114) );
  MXI2X1 U7473 ( .A(U1_pipe8[16]), .B(n20241), .S0(n20240), .Y(n4997) );
  XNOR2X1 U7474 ( .A(n16840), .B(n16839), .Y(n16841) );
  INVX1 U7475 ( .A(n24742), .Y(n24750) );
  NOR2X1 U7476 ( .A(n16788), .B(n14970), .Y(n14971) );
  XNOR2X1 U7477 ( .A(n25180), .B(n25179), .Y(n25181) );
  XNOR2X1 U7478 ( .A(n17489), .B(n17488), .Y(n17490) );
  XOR2X1 U7479 ( .A(n24764), .B(n24763), .Y(n24765) );
  NAND2BX1 U7480 ( .AN(n20330), .B(n20332), .Y(n7873) );
  INVX1 U7481 ( .A(n16787), .Y(n5943) );
  NAND2X1 U7482 ( .A(n7753), .B(n7561), .Y(n6350) );
  NAND2X1 U7483 ( .A(n16791), .B(n16790), .Y(n17055) );
  XNOR2X1 U7484 ( .A(n14054), .B(n14104), .Y(n14055) );
  XNOR2X1 U7485 ( .A(n17500), .B(n17499), .Y(n17501) );
  XNOR2X1 U7486 ( .A(n16676), .B(n16675), .Y(n16677) );
  XOR2X1 U7487 ( .A(n24769), .B(n24768), .Y(n24770) );
  XOR2X1 U7488 ( .A(n25360), .B(n25359), .Y(n25361) );
  NAND3X1 U7489 ( .A(n19409), .B(n13708), .C(n7685), .Y(n7687) );
  XOR2X1 U7490 ( .A(n24458), .B(n24457), .Y(n24459) );
  BUFX2 U7491 ( .A(n25286), .Y(n7729) );
  XOR2X1 U7492 ( .A(n22651), .B(n22650), .Y(n22652) );
  XNOR2X1 U7493 ( .A(n21868), .B(n21867), .Y(n21869) );
  XOR2X1 U7494 ( .A(n24471), .B(n24470), .Y(n24472) );
  XOR2X1 U7495 ( .A(n22012), .B(n22011), .Y(n22013) );
  NAND3BX2 U7496 ( .AN(n14121), .B(n6243), .C(n6242), .Y(n22599) );
  XOR2X1 U7497 ( .A(n23039), .B(n23038), .Y(n23040) );
  XOR2X1 U7498 ( .A(n23045), .B(n23044), .Y(n23046) );
  AND2X2 U7499 ( .A(n7842), .B(n7337), .Y(n6061) );
  AND2X2 U7500 ( .A(n20331), .B(n20332), .Y(n20338) );
  AOI2BB1X2 U7501 ( .A0N(n22623), .A1N(n14112), .B0(n12636), .Y(n22619) );
  NAND2X1 U7502 ( .A(n19077), .B(n19076), .Y(n19390) );
  XNOR2X1 U7503 ( .A(n20087), .B(n20086), .Y(n20088) );
  MXI2X1 U7504 ( .A(U0_pipe6[21]), .B(n21838), .S0(n20240), .Y(n4469) );
  XOR2X1 U7505 ( .A(n19270), .B(n19269), .Y(n19271) );
  AOI21X1 U7506 ( .A0(n14009), .A1(n6046), .B0(n5963), .Y(n5962) );
  XOR2X1 U7507 ( .A(n22018), .B(n22017), .Y(n22019) );
  INVX1 U7508 ( .A(n16783), .Y(n16781) );
  XOR2X1 U7509 ( .A(n22645), .B(n22644), .Y(n22646) );
  XNOR2X1 U7510 ( .A(n21858), .B(n21857), .Y(n21859) );
  AOI21X1 U7511 ( .A0(n17630), .A1(n17628), .B0(n14502), .Y(n6153) );
  AOI21X1 U7512 ( .A0(n5966), .A1(n17086), .B0(n17085), .Y(n17095) );
  XNOR2X1 U7513 ( .A(n20370), .B(n20369), .Y(n20371) );
  INVX1 U7514 ( .A(n20069), .Y(n20077) );
  XOR2X1 U7515 ( .A(n22623), .B(n22630), .Y(n22631) );
  AOI21X1 U7516 ( .A0(n22655), .A1(n22635), .B0(n22634), .Y(n22645) );
  MXI2X1 U7517 ( .A(U1_pipe13[13]), .B(n20102), .S0(n20025), .Y(n4736) );
  XNOR2X1 U7518 ( .A(n24475), .B(n24474), .Y(n24476) );
  XNOR2X1 U7519 ( .A(n16686), .B(n16685), .Y(n16687) );
  MXI2X1 U7520 ( .A(U1_pipe8[14]), .B(n20249), .S0(n20240), .Y(n4995) );
  XOR2X1 U7521 ( .A(n20092), .B(n20091), .Y(n20093) );
  INVX1 U7522 ( .A(n5998), .Y(n16809) );
  INVX1 U7523 ( .A(n6032), .Y(n5963) );
  INVX1 U7524 ( .A(n21851), .Y(n21858) );
  XNOR2X1 U7525 ( .A(n24486), .B(n24485), .Y(n24487) );
  NAND2BX1 U7526 ( .AN(n25528), .B(U2_A_i_d[25]), .Y(n6699) );
  INVX1 U7527 ( .A(n17491), .Y(n17500) );
  XOR2X1 U7528 ( .A(n17655), .B(n17654), .Y(n17656) );
  XOR2X1 U7529 ( .A(n22048), .B(n22047), .Y(n22049) );
  MXI2X1 U7530 ( .A(U1_pipe8[15]), .B(n20244), .S0(n20240), .Y(n4996) );
  XOR2X1 U7531 ( .A(n17688), .B(n17687), .Y(n17689) );
  XOR2X1 U7532 ( .A(n17673), .B(n17672), .Y(n17674) );
  NAND2X1 U7533 ( .A(n20321), .B(n20344), .Y(n20349) );
  XOR2X1 U7534 ( .A(n22032), .B(n22031), .Y(n22033) );
  XNOR2X1 U7535 ( .A(n22655), .B(n22654), .Y(n22656) );
  NAND2XL U7536 ( .A(n7906), .B(n19566), .Y(n7875) );
  XNOR2X1 U7537 ( .A(n24463), .B(n24462), .Y(n24464) );
  XOR2X1 U7538 ( .A(n22777), .B(n22776), .Y(n22778) );
  XOR2X1 U7539 ( .A(n17366), .B(n17365), .Y(n17367) );
  XOR2X1 U7540 ( .A(n17660), .B(n17659), .Y(n17661) );
  XNOR2X1 U7541 ( .A(n19136), .B(n19135), .Y(n19137) );
  NOR2XL U7542 ( .A(n5815), .B(n22884), .Y(n6858) );
  XNOR2X1 U7543 ( .A(n24773), .B(n24772), .Y(n24774) );
  XNOR2X1 U7544 ( .A(n25581), .B(n25580), .Y(n25582) );
  XOR2X1 U7545 ( .A(n16879), .B(n16878), .Y(n16880) );
  XNOR2X1 U7546 ( .A(n25370), .B(n25369), .Y(n25371) );
  NAND2BXL U7547 ( .AN(n19075), .B(n14895), .Y(n7747) );
  NAND2XL U7548 ( .A(n14898), .B(n19385), .Y(n14899) );
  XNOR2X1 U7549 ( .A(n25569), .B(n25568), .Y(n25570) );
  XNOR2X1 U7550 ( .A(n19284), .B(n19283), .Y(n19285) );
  AND2X2 U7551 ( .A(n20060), .B(n6013), .Y(n6012) );
  XNOR2X1 U7552 ( .A(n19274), .B(n19273), .Y(n19275) );
  NAND2X2 U7553 ( .A(n6380), .B(n12392), .Y(n25321) );
  XNOR2X1 U7554 ( .A(n23049), .B(n23048), .Y(n23050) );
  NAND2XL U7555 ( .A(n17461), .B(n9539), .Y(n17457) );
  XOR2X1 U7556 ( .A(n16845), .B(n16844), .Y(n16846) );
  XOR2X1 U7557 ( .A(n16851), .B(n16850), .Y(n16852) );
  NAND2XL U7558 ( .A(n12342), .B(n6299), .Y(n6298) );
  AND2X2 U7559 ( .A(n21958), .B(n14576), .Y(n6445) );
  AOI21X1 U7560 ( .A0(n19265), .A1(n19263), .B0(n19258), .Y(n6005) );
  XOR2X1 U7561 ( .A(n22355), .B(n22354), .Y(n22356) );
  XNOR2X1 U7562 ( .A(n16883), .B(n16882), .Y(n16884) );
  NAND2X1 U7563 ( .A(n25315), .B(n25669), .Y(n25674) );
  MXI2X1 U7564 ( .A(U1_pipe2[13]), .B(n19151), .S0(n19215), .Y(n5025) );
  NOR2X1 U7565 ( .A(n16634), .B(n6519), .Y(n6518) );
  INVX1 U7566 ( .A(n24705), .Y(n6299) );
  NAND2X1 U7567 ( .A(n20061), .B(n6915), .Y(n6013) );
  NAND2BX1 U7568 ( .AN(n20041), .B(n5845), .Y(n20019) );
  NAND2BX1 U7569 ( .AN(n14944), .B(n5999), .Y(n5998) );
  NAND2BX1 U7570 ( .AN(n20345), .B(n20324), .Y(n20341) );
  XOR2X1 U7571 ( .A(n25393), .B(n25392), .Y(n25394) );
  XNOR2X1 U7572 ( .A(n22781), .B(n22780), .Y(n22782) );
  XNOR2X1 U7573 ( .A(n22791), .B(n22790), .Y(n22792) );
  XOR2X1 U7574 ( .A(n25379), .B(n25378), .Y(n25380) );
  INVX2 U7575 ( .A(n14577), .Y(n13178) );
  MXI2X1 U7576 ( .A(U1_pipe8[13]), .B(n20252), .S0(n20240), .Y(n4994) );
  XNOR2X1 U7577 ( .A(n17678), .B(n17677), .Y(n17679) );
  XNOR2X1 U7578 ( .A(n22052), .B(n22051), .Y(n22053) );
  MXI2X1 U7579 ( .A(U0_pipe2[13]), .B(n24502), .S0(n24784), .Y(n4390) );
  NAND2XL U7580 ( .A(n16804), .B(n17063), .Y(n17068) );
  XNOR2X1 U7581 ( .A(n22036), .B(n22035), .Y(n22037) );
  INVXL U7582 ( .A(n16800), .Y(n7472) );
  NAND2X1 U7583 ( .A(n14513), .B(n19233), .Y(n17597) );
  XNOR2X1 U7584 ( .A(n16867), .B(n16866), .Y(n16868) );
  MXI2X1 U7585 ( .A(U0_pipe4[13]), .B(n22237), .S0(n22543), .Y(n4334) );
  NAND2X1 U7586 ( .A(n6419), .B(n6256), .Y(n6255) );
  NAND2X1 U7587 ( .A(n19244), .B(n19561), .Y(n19581) );
  XOR2X1 U7588 ( .A(n7380), .B(n7027), .Y(n18910) );
  NAND2BXL U7589 ( .AN(n14575), .B(n5858), .Y(n14576) );
  XOR2X1 U7590 ( .A(n20110), .B(n20109), .Y(n20111) );
  XOR2X1 U7591 ( .A(n20125), .B(n20124), .Y(n20126) );
  XOR2X1 U7592 ( .A(n24511), .B(n24510), .Y(n24512) );
  INVX1 U7593 ( .A(n20319), .Y(n6054) );
  INVXL U7594 ( .A(n17664), .Y(n14506) );
  NAND2XL U7595 ( .A(n19822), .B(n19772), .Y(n6653) );
  NAND2X1 U7596 ( .A(n24716), .B(n24715), .Y(n24994) );
  NAND2X1 U7597 ( .A(n16819), .B(n6936), .Y(n13948) );
  NOR2X1 U7598 ( .A(n13716), .B(U1_A_r_d0[24]), .Y(n19075) );
  NAND2X1 U7599 ( .A(n13716), .B(U1_A_r_d0[24]), .Y(n19076) );
  NAND2X1 U7600 ( .A(n20029), .B(n19233), .Y(n19565) );
  OAI21X1 U7601 ( .A0(n13945), .A1(n17084), .B0(n13944), .Y(n14006) );
  NAND2XL U7602 ( .A(n24693), .B(n24692), .Y(n12341) );
  AOI21X1 U7603 ( .A0(n17230), .A1(n17214), .B0(n17213), .Y(n17222) );
  XOR2X1 U7604 ( .A(n17379), .B(n17378), .Y(n17380) );
  NAND2X1 U7605 ( .A(n17185), .B(n17184), .Y(n17465) );
  XOR2X1 U7606 ( .A(n19308), .B(n19307), .Y(n19309) );
  AND2X2 U7607 ( .A(n20016), .B(n14851), .Y(n20345) );
  MXI2X1 U7608 ( .A(U0_pipe13[8]), .B(n25403), .S0(n24784), .Y(n4684) );
  OR2X2 U7609 ( .A(n5851), .B(n29008), .Y(n6610) );
  XNOR2X1 U7610 ( .A(n25383), .B(n25382), .Y(n25384) );
  NAND2BX2 U7611 ( .AN(n13552), .B(n5950), .Y(n17370) );
  NAND2X1 U7612 ( .A(n6987), .B(n21969), .Y(n22311) );
  NAND2BX1 U7613 ( .AN(n20015), .B(n5817), .Y(n7025) );
  NOR2X1 U7614 ( .A(n16834), .B(n16836), .Y(n5999) );
  XNOR2X1 U7615 ( .A(n17383), .B(n17382), .Y(n17384) );
  INVXL U7616 ( .A(n13966), .Y(n16802) );
  NAND2X1 U7617 ( .A(n25133), .B(n25522), .Y(n25533) );
  NAND2X1 U7618 ( .A(n5853), .B(n5817), .Y(n6936) );
  NAND2BX2 U7619 ( .AN(n5817), .B(n5857), .Y(n20061) );
  MXI2X1 U7620 ( .A(U0_pipe14[13]), .B(n22520), .S0(n22543), .Y(n4651) );
  XNOR2X1 U7621 ( .A(n17397), .B(n17396), .Y(n17398) );
  NAND2XL U7622 ( .A(n14974), .B(U1_A_r_d0[25]), .Y(n14898) );
  NOR2X1 U7623 ( .A(n20363), .B(n14887), .Y(n20310) );
  NAND2X1 U7624 ( .A(n25339), .B(n25338), .Y(n25694) );
  XOR2X1 U7625 ( .A(n22663), .B(n22662), .Y(n22664) );
  INVX1 U7626 ( .A(n22773), .Y(n22781) );
  INVXL U7627 ( .A(n20029), .Y(n14863) );
  XOR2X1 U7628 ( .A(n17533), .B(n17532), .Y(n17534) );
  NAND2X1 U7629 ( .A(n20033), .B(n19237), .Y(n19563) );
  XOR2X1 U7630 ( .A(n22801), .B(n22800), .Y(n22802) );
  XNOR2X1 U7631 ( .A(n19856), .B(n19855), .Y(n19857) );
  NAND2X1 U7632 ( .A(n16819), .B(n16818), .Y(n17071) );
  NAND2XL U7633 ( .A(n14503), .B(n14501), .Y(n13095) );
  NOR2X1 U7634 ( .A(n20048), .B(n5850), .Y(n20018) );
  XOR2X1 U7635 ( .A(n19160), .B(n19159), .Y(n19161) );
  NAND2X1 U7636 ( .A(n19112), .B(n19414), .Y(n19419) );
  NAND2X1 U7637 ( .A(n24677), .B(n24687), .Y(n24705) );
  MXI2X1 U7638 ( .A(U0_pipe0[13]), .B(n24918), .S0(n5920), .Y(n4299) );
  XOR2X1 U7639 ( .A(n23058), .B(n23057), .Y(n23059) );
  MXI2X1 U7640 ( .A(U1_pipe13[8]), .B(n20135), .S0(n20025), .Y(n4731) );
  XNOR2X1 U7641 ( .A(n20130), .B(n20129), .Y(n20131) );
  NOR2X1 U7642 ( .A(n20016), .B(n20051), .Y(n20046) );
  XNOR2X1 U7643 ( .A(n20115), .B(n20114), .Y(n20116) );
  XOR2X1 U7644 ( .A(n19324), .B(n19323), .Y(n19325) );
  NAND2X1 U7645 ( .A(n25332), .B(n25683), .Y(n25688) );
  XNOR2X1 U7646 ( .A(n21484), .B(n21483), .Y(n21485) );
  XNOR2X1 U7647 ( .A(n24515), .B(n24514), .Y(n24516) );
  XOR2X1 U7648 ( .A(n25730), .B(n25729), .Y(n25731) );
  XOR2X1 U7649 ( .A(n25745), .B(n25744), .Y(n25746) );
  INVX1 U7650 ( .A(n21991), .Y(n13129) );
  XOR2X1 U7651 ( .A(n20409), .B(n20408), .Y(n20410) );
  XNOR2X1 U7652 ( .A(n21367), .B(n21366), .Y(n21368) );
  XOR2X1 U7653 ( .A(n24783), .B(n24782), .Y(n24785) );
  MXI2XL U7654 ( .A(n6268), .B(U2_pipe3[18]), .S0(n5929), .Y(n4235) );
  NAND2X1 U7655 ( .A(n20308), .B(n20311), .Y(n20352) );
  XNOR2X1 U7656 ( .A(n22667), .B(n22666), .Y(n22668) );
  XNOR2X1 U7657 ( .A(n19313), .B(n19312), .Y(n19314) );
  NAND2X1 U7658 ( .A(n22957), .B(n13166), .Y(n22309) );
  INVXL U7659 ( .A(n9142), .Y(n6343) );
  XOR2X1 U7660 ( .A(n19176), .B(n19175), .Y(n19177) );
  MXI2X1 U7661 ( .A(U1_pipe1[11]), .B(n19649), .S0(n20025), .Y(n5142) );
  NAND2X1 U7662 ( .A(n16650), .B(n16950), .Y(n16955) );
  NAND2BXL U7663 ( .AN(n14562), .B(n22932), .Y(n21991) );
  XOR2X1 U7664 ( .A(n24800), .B(n24799), .Y(n24801) );
  INVXL U7665 ( .A(n14972), .Y(n14513) );
  XOR2X1 U7666 ( .A(n22676), .B(n22675), .Y(n22677) );
  XNOR2X1 U7667 ( .A(n19164), .B(n19163), .Y(n19165) );
  NAND2X1 U7668 ( .A(n22470), .B(n22469), .Y(n22747) );
  XOR2X1 U7669 ( .A(n25214), .B(n25213), .Y(n25215) );
  MXI2X1 U7670 ( .A(U0_pipe5[8]), .B(n22385), .S0(n6888), .Y(n4311) );
  INVX1 U7671 ( .A(n22330), .Y(n21996) );
  INVX1 U7672 ( .A(n24724), .Y(n5849) );
  NAND2X1 U7673 ( .A(n22613), .B(n22612), .Y(n22995) );
  INVXL U7674 ( .A(n16825), .Y(n5969) );
  OR2X2 U7675 ( .A(n19617), .B(n19549), .Y(n6110) );
  OR2X2 U7676 ( .A(n12332), .B(U1_A_r_d0[24]), .Y(n19797) );
  INVX1 U7677 ( .A(n6062), .Y(n16826) );
  XOR2X1 U7678 ( .A(n21360), .B(n21313), .Y(n21314) );
  XOR2X1 U7679 ( .A(n6269), .B(n18655), .Y(n6268) );
  XOR2X1 U7680 ( .A(n21478), .B(n21427), .Y(n21428) );
  NAND2BX1 U7681 ( .AN(n14943), .B(n5975), .Y(n5977) );
  XOR2X1 U7682 ( .A(n21534), .B(n21533), .Y(n21535) );
  AND2X2 U7683 ( .A(n25716), .B(n25714), .Y(n6476) );
  XOR2X1 U7684 ( .A(n7541), .B(n7026), .Y(n26913) );
  XNOR2X1 U7685 ( .A(n20399), .B(n20398), .Y(n20400) );
  XOR2X1 U7686 ( .A(n26825), .B(n26824), .Y(n26826) );
  XOR2X1 U7687 ( .A(n22814), .B(n22813), .Y(n22815) );
  MXI2X1 U7688 ( .A(U0_pipe10[11]), .B(n22819), .S0(n22853), .Y(n4566) );
  XOR2X1 U7689 ( .A(n22828), .B(n22827), .Y(n22829) );
  MXI2X1 U7690 ( .A(U0_pipe10[9]), .B(n22833), .S0(n22853), .Y(n4568) );
  NAND2BX1 U7691 ( .AN(n14854), .B(n7275), .Y(n7274) );
  XNOR2X1 U7692 ( .A(n17537), .B(n17536), .Y(n17538) );
  XOR2X1 U7693 ( .A(n17547), .B(n17546), .Y(n17548) );
  NAND2X1 U7694 ( .A(n17341), .B(n17340), .Y(n17634) );
  XOR2X1 U7695 ( .A(n21271), .B(n21270), .Y(n21272) );
  NAND2X1 U7696 ( .A(n19763), .B(n19753), .Y(n19764) );
  XNOR2X1 U7697 ( .A(n20414), .B(n20413), .Y(n20415) );
  XOR2X1 U7698 ( .A(n24527), .B(n24526), .Y(n24528) );
  MXI2X1 U7699 ( .A(U1_pipe9[8]), .B(n20418), .S0(n21972), .Y(n4818) );
  XNOR2X1 U7700 ( .A(n23062), .B(n23061), .Y(n23063) );
  INVX1 U7701 ( .A(n25684), .Y(n25332) );
  NAND2X1 U7702 ( .A(n24426), .B(n24425), .Y(n24870) );
  NOR2X1 U7703 ( .A(n8609), .B(n16975), .Y(n16958) );
  XOR2X1 U7704 ( .A(n21888), .B(n21887), .Y(n21889) );
  XOR2X1 U7705 ( .A(n26651), .B(n26650), .Y(n26652) );
  XNOR2X1 U7706 ( .A(n19328), .B(n19327), .Y(n19329) );
  XOR2X1 U7707 ( .A(n26707), .B(n26706), .Y(n26708) );
  XOR2X1 U7708 ( .A(n23072), .B(n23071), .Y(n23073) );
  AOI21X1 U7709 ( .A0(n24917), .A1(n24902), .B0(n24901), .Y(n24909) );
  MXI2X1 U7710 ( .A(U0_pipe9[8]), .B(n25754), .S0(n6887), .Y(n4597) );
  XNOR2X1 U7711 ( .A(n25750), .B(n25749), .Y(n25751) );
  MXI2X1 U7712 ( .A(U0_pipe2[9]), .B(n24532), .S0(n22853), .Y(n4394) );
  NAND2X1 U7713 ( .A(n19094), .B(n19093), .Y(n19400) );
  XOR2X1 U7714 ( .A(n26765), .B(n26764), .Y(n26766) );
  XOR2X2 U7715 ( .A(n13654), .B(n13643), .Y(n14972) );
  INVX1 U7716 ( .A(n17372), .Y(n17401) );
  MXI2X1 U7717 ( .A(U1_pipe15[7]), .B(n17409), .S0(n6887), .Y(n4786) );
  NAND2X1 U7718 ( .A(n19552), .B(n19550), .Y(n19611) );
  MXI2X1 U7719 ( .A(U1_pipe15[6]), .B(n17417), .S0(n17187), .Y(n4785) );
  NAND2X1 U7720 ( .A(n24643), .B(n13128), .Y(n25691) );
  MXI2X1 U7721 ( .A(U0_pipe4[10]), .B(n22257), .S0(n22248), .Y(n4337) );
  MXI2X1 U7722 ( .A(U0_pipe4[11]), .B(n22249), .S0(n22248), .Y(n4336) );
  AND2XL U7723 ( .A(n14484), .B(U2_A_r_d[23]), .Y(n14485) );
  MXI2X1 U7724 ( .A(U0_pipe2[8]), .B(n24536), .S0(n22853), .Y(n4395) );
  MXI2X1 U7725 ( .A(U0_pipe1[8]), .B(n25071), .S0(n25091), .Y(n4276) );
  NOR2X1 U7726 ( .A(n5819), .B(n6344), .Y(n9142) );
  MXI2X1 U7727 ( .A(U0_pipe1[7]), .B(n25078), .S0(n25091), .Y(n4277) );
  NAND2X1 U7728 ( .A(n25516), .B(n25514), .Y(n25544) );
  XNOR2X1 U7729 ( .A(n23077), .B(n23076), .Y(n23078) );
  INVX1 U7730 ( .A(n20103), .Y(n20134) );
  MXI2X1 U7731 ( .A(U1_pipe12[9]), .B(n19901), .S0(n20025), .Y(n4903) );
  MXI2X1 U7732 ( .A(U1_pipe13[7]), .B(n20142), .S0(n20025), .Y(n4730) );
  MXI2X1 U7733 ( .A(U1_pipe13[6]), .B(n20150), .S0(n20025), .Y(n4729) );
  XOR2X1 U7734 ( .A(n19896), .B(n19895), .Y(n19897) );
  MXI2X1 U7735 ( .A(U1_pipe8[12]), .B(n20259), .S0(n20240), .Y(n4993) );
  MXI2X1 U7736 ( .A(U1_pipe12[11]), .B(n19885), .S0(n20025), .Y(n4905) );
  XOR2X1 U7737 ( .A(n19880), .B(n19879), .Y(n19881) );
  MXI2X1 U7738 ( .A(U1_pipe8[10]), .B(n20270), .S0(n20240), .Y(n4991) );
  XNOR2X1 U7739 ( .A(n25218), .B(n25217), .Y(n25219) );
  XOR2X1 U7740 ( .A(n25229), .B(n25228), .Y(n25230) );
  MXI2X1 U7741 ( .A(U1_pipe14[9]), .B(n17254), .S0(n22853), .Y(n4760) );
  INVX1 U7742 ( .A(n24640), .Y(n6783) );
  INVX1 U7743 ( .A(n20083), .Y(n20090) );
  MXI2X1 U7744 ( .A(U0_pipe13[7]), .B(n25410), .S0(n25611), .Y(n4685) );
  MXI2X1 U7745 ( .A(U0_pipe10[8]), .B(n22837), .S0(n22853), .Y(n4569) );
  MXI2X1 U7746 ( .A(U0_pipe13[6]), .B(n25418), .S0(n22853), .Y(n4686) );
  NAND2X1 U7747 ( .A(n5859), .B(n14954), .Y(n16837) );
  NAND2X1 U7748 ( .A(n5796), .B(n22435), .Y(n14104) );
  AOI21X1 U7749 ( .A0(n14541), .A1(n14540), .B0(n14539), .Y(n22025) );
  XNOR2X1 U7750 ( .A(n22542), .B(n22830), .Y(n22544) );
  AND2XL U7751 ( .A(n14484), .B(U2_A_i_d[23]), .Y(n21798) );
  XNOR2X1 U7752 ( .A(n21892), .B(n21891), .Y(n21893) );
  XOR2X1 U7753 ( .A(n21902), .B(n21901), .Y(n21903) );
  MXI2X1 U7754 ( .A(U1_pipe4[9]), .B(n17014), .S0(n24784), .Y(n5077) );
  XOR2X1 U7755 ( .A(n23987), .B(n23986), .Y(n23988) );
  XOR2X1 U7756 ( .A(n24045), .B(n24044), .Y(n24046) );
  AND2XL U7757 ( .A(n9501), .B(U1_A_i_d0[14]), .Y(n9502) );
  XOR2X1 U7758 ( .A(n16710), .B(n16709), .Y(n16711) );
  NAND2XL U7759 ( .A(n19998), .B(n20011), .Y(n20071) );
  MXI2X1 U7760 ( .A(U1_pipe2[8]), .B(n19185), .S0(n19215), .Y(n5020) );
  XNOR2X1 U7761 ( .A(n22681), .B(n22680), .Y(n22682) );
  XOR2X1 U7762 ( .A(n16726), .B(n16725), .Y(n16727) );
  XOR2X1 U7763 ( .A(n18552), .B(n18551), .Y(n18553) );
  INVX1 U7764 ( .A(n21832), .Y(n22168) );
  NOR2X1 U7765 ( .A(n5859), .B(n14954), .Y(n14944) );
  NAND2XL U7766 ( .A(n16836), .B(n16842), .Y(n7465) );
  XOR2X1 U7767 ( .A(n18822), .B(n18821), .Y(n18823) );
  CLKINVX3 U7768 ( .A(n19775), .Y(n19774) );
  INVX1 U7769 ( .A(n19252), .Y(n7275) );
  MXI2X1 U7770 ( .A(U0_pipe7[6]), .B(n22072), .S0(n21972), .Y(n4456) );
  NAND2X1 U7771 ( .A(n14957), .B(n19998), .Y(n16825) );
  MXI2X1 U7772 ( .A(U0_pipe0[8]), .B(n24942), .S0(n5920), .Y(n4304) );
  XOR2X1 U7773 ( .A(n24165), .B(n24164), .Y(n24166) );
  INVXL U7774 ( .A(n20041), .Y(n6123) );
  XOR2X1 U7775 ( .A(n24288), .B(n24252), .Y(n24253) );
  MXI2X1 U7776 ( .A(U0_pipe3[8]), .B(n24809), .S0(n24784), .Y(n4367) );
  XNOR2X1 U7777 ( .A(n24804), .B(n24803), .Y(n24805) );
  XNOR2X1 U7778 ( .A(n18406), .B(n18364), .Y(n18365) );
  MXI2X1 U7779 ( .A(U0_pipe1[6]), .B(n25086), .S0(n25091), .Y(n4278) );
  MXI2X1 U7780 ( .A(U0_pipe7[7]), .B(n22064), .S0(n21972), .Y(n4455) );
  NAND2X1 U7781 ( .A(n6511), .B(n22807), .Y(n6510) );
  NAND2X1 U7782 ( .A(n13694), .B(U1_A_i_d0[15]), .Y(n17220) );
  INVX1 U7783 ( .A(n14957), .Y(n13069) );
  MXI2X1 U7784 ( .A(U0_pipe6[8]), .B(n21909), .S0(n20438), .Y(n4482) );
  MXI2X1 U7785 ( .A(U0_pipe2[7]), .B(n24544), .S0(n22853), .Y(n4396) );
  XOR2X1 U7786 ( .A(n20908), .B(n20907), .Y(n20909) );
  MXI2X1 U7787 ( .A(U0_pipe13[5]), .B(n25423), .S0(n6887), .Y(n4687) );
  MXI2X1 U7788 ( .A(U0_pipe7[5]), .B(n22077), .S0(n21972), .Y(n4457) );
  XOR2X1 U7789 ( .A(n26409), .B(n26408), .Y(n26410) );
  INVX1 U7790 ( .A(n25140), .Y(n14484) );
  MXI2X1 U7791 ( .A(U1_pipe0[6]), .B(n19485), .S0(n19215), .Y(n5109) );
  MXI2X1 U7792 ( .A(U0_pipe10[7]), .B(n22845), .S0(n22853), .Y(n4570) );
  MXI2X1 U7793 ( .A(U0_pipe11[7]), .B(n23090), .S0(n24784), .Y(n4542) );
  MXI2X1 U7794 ( .A(U0_pipe11[6]), .B(n23098), .S0(n24784), .Y(n4543) );
  AOI21X1 U7795 ( .A0(n19293), .A1(n19291), .B0(n14827), .Y(n19277) );
  MXI2X1 U7796 ( .A(U1_pipe3[7]), .B(n19341), .S0(n19215), .Y(n5047) );
  MXI2X1 U7797 ( .A(U1_pipe9[7]), .B(n20425), .S0(n21972), .Y(n4817) );
  NAND2XL U7798 ( .A(n14939), .B(n14938), .Y(n5976) );
  OR2X2 U7799 ( .A(n17667), .B(n12973), .Y(n6029) );
  NAND2X1 U7800 ( .A(n12327), .B(U1_A_i_d0[21]), .Y(n16950) );
  NAND2X1 U7801 ( .A(n24679), .B(n22957), .Y(n22612) );
  MXI2X1 U7802 ( .A(U0_pipe6[6]), .B(n21923), .S0(n21972), .Y(n4484) );
  NAND2BX1 U7803 ( .AN(n22931), .B(n5819), .Y(n22617) );
  MXI2X1 U7804 ( .A(U1_pipe0[7]), .B(n19479), .S0(n19215), .Y(n5110) );
  MXI2X1 U7805 ( .A(U0_pipe6[7]), .B(n21915), .S0(n21972), .Y(n4483) );
  MXI2X1 U7806 ( .A(U0_pipe2[6]), .B(n24552), .S0(n22853), .Y(n4397) );
  MXI2X1 U7807 ( .A(U0_pipe9[6]), .B(n25769), .S0(n6887), .Y(n4599) );
  MXI2X1 U7808 ( .A(U0_pipe9[7]), .B(n25761), .S0(n6887), .Y(n4598) );
  MXI2X1 U7809 ( .A(U0_pipe3[7]), .B(n24816), .S0(n24784), .Y(n4368) );
  INVXL U7810 ( .A(n17364), .Y(n7519) );
  NAND2X1 U7811 ( .A(n7914), .B(n20011), .Y(n14834) );
  XOR2X1 U7812 ( .A(n21069), .B(n20963), .Y(n20964) );
  XOR2X1 U7813 ( .A(n21022), .B(n21021), .Y(n21024) );
  AOI21X1 U7814 ( .A0(n22521), .A1(n14039), .B0(n14038), .Y(n22446) );
  XOR2X1 U7815 ( .A(n18359), .B(n18257), .Y(n18258) );
  XOR2X1 U7816 ( .A(n18308), .B(n18307), .Y(n18309) );
  MXI2X1 U7817 ( .A(U1_pipe0[8]), .B(n19473), .S0(n19215), .Y(n5111) );
  MXI2X1 U7818 ( .A(U1_pipe9[6]), .B(n20433), .S0(n21972), .Y(n4816) );
  AND2X2 U7819 ( .A(n7492), .B(n6000), .Y(n7145) );
  XNOR2X1 U7820 ( .A(n21905), .B(n21904), .Y(n21906) );
  NAND2X1 U7821 ( .A(n24461), .B(n24460), .Y(n24887) );
  OR2X2 U7822 ( .A(n14956), .B(n14955), .Y(n14949) );
  XOR2X1 U7823 ( .A(n26459), .B(n26359), .Y(n26361) );
  MXI2X1 U7824 ( .A(U2_pipe3[8]), .B(n18099), .S0(n8054), .Y(n4215) );
  XOR2X1 U7825 ( .A(n26296), .B(n26295), .Y(n26297) );
  MXI2X1 U7826 ( .A(U0_pipe3[6]), .B(n24824), .S0(n24784), .Y(n4369) );
  XNOR2X1 U7827 ( .A(n19900), .B(n19899), .Y(n19901) );
  INVX1 U7828 ( .A(n20015), .Y(n5857) );
  NAND2X1 U7829 ( .A(n7914), .B(n7913), .Y(n19552) );
  NAND2X1 U7830 ( .A(n7018), .B(n13881), .Y(n13887) );
  MXI2X1 U7831 ( .A(U0_pipe15[5]), .B(n22706), .S0(n22620), .Y(n4631) );
  XNOR2X1 U7832 ( .A(n16714), .B(n16713), .Y(n16715) );
  MXI2X1 U7833 ( .A(U1_pipe14[6]), .B(n17272), .S0(n22853), .Y(n4757) );
  MXI2X1 U7834 ( .A(U1_pipe8[11]), .B(n20262), .S0(n20240), .Y(n4992) );
  MXI2X1 U7835 ( .A(U1_pipe14[7]), .B(n17265), .S0(n22853), .Y(n4758) );
  MXI2X1 U7836 ( .A(U1_pipe8[9]), .B(n20273), .S0(n20240), .Y(n4990) );
  NAND2X1 U7837 ( .A(n5867), .B(n19993), .Y(n20085) );
  MXI2X1 U7838 ( .A(U1_pipe14[8]), .B(n17258), .S0(n22853), .Y(n4759) );
  MXI2X1 U7839 ( .A(U0_pipe5[6]), .B(n22400), .S0(n22620), .Y(n4313) );
  XNOR2X1 U7840 ( .A(n25233), .B(n25232), .Y(n25234) );
  MXI2X1 U7841 ( .A(U1_pipe15[5]), .B(n17422), .S0(n6887), .Y(n4784) );
  MXI2X1 U7842 ( .A(U1_pipe2[6]), .B(n19202), .S0(n19215), .Y(n5018) );
  INVX1 U7843 ( .A(n20367), .Y(n20373) );
  OR2X2 U7844 ( .A(n24654), .B(n24644), .Y(n7014) );
  XNOR2X1 U7845 ( .A(n24158), .B(n23940), .Y(n23941) );
  MXI2X1 U7846 ( .A(U1_pipe3[6]), .B(n19349), .S0(n19405), .Y(n5046) );
  MXI2X1 U7847 ( .A(U0_pipe4[9]), .B(n22260), .S0(n22248), .Y(n4338) );
  INVX1 U7848 ( .A(n22476), .Y(n7612) );
  INVX1 U7849 ( .A(n20383), .Y(n20377) );
  MXI2X1 U7850 ( .A(U1_pipe2[7]), .B(n19192), .S0(n19215), .Y(n5019) );
  OR2X2 U7851 ( .A(n13037), .B(n19282), .Y(n13009) );
  AND2XL U7852 ( .A(n13037), .B(n19282), .Y(n8145) );
  OR2X2 U7853 ( .A(n5869), .B(n19542), .Y(n13025) );
  MXI2X1 U7854 ( .A(U1_pipe3[5]), .B(n19354), .S0(n19405), .Y(n5045) );
  NAND2X1 U7855 ( .A(n6991), .B(n17236), .Y(n17531) );
  MXI2X1 U7856 ( .A(U1_pipe3[4]), .B(n19362), .S0(n19405), .Y(n5044) );
  MXI2X1 U7857 ( .A(U0_pipe0[7]), .B(n24950), .S0(n5920), .Y(n4305) );
  MXI2X1 U7858 ( .A(U0_pipe0[6]), .B(n24958), .S0(n5920), .Y(n4306) );
  NAND2X1 U7859 ( .A(n24664), .B(n22931), .Y(n22616) );
  MXI2X1 U7860 ( .A(U1_pipe2[5]), .B(n19206), .S0(n19215), .Y(n5017) );
  NAND2X1 U7861 ( .A(n24661), .B(n22933), .Y(n22628) );
  MXI2X1 U7862 ( .A(U0_pipe4[8]), .B(n22263), .S0(n22248), .Y(n4339) );
  NOR2X1 U7863 ( .A(n19272), .B(n7843), .Y(n19610) );
  MXI2X1 U7864 ( .A(U0_pipe12[5]), .B(n25259), .S0(n25267), .Y(n4516) );
  XOR2X1 U7865 ( .A(n23639), .B(n23638), .Y(n23640) );
  NAND2X1 U7866 ( .A(n14950), .B(n14946), .Y(n17103) );
  CLKINVX3 U7867 ( .A(n20011), .Y(n7913) );
  CLKINVX3 U7868 ( .A(n7915), .Y(n7914) );
  NAND2X1 U7869 ( .A(n24484), .B(n24488), .Y(n13518) );
  NAND2X1 U7870 ( .A(n14955), .B(n5865), .Y(n17639) );
  XOR2X1 U7871 ( .A(n23794), .B(n23694), .Y(n23696) );
  NAND2X1 U7872 ( .A(n20108), .B(n20113), .Y(n19990) );
  NAND2XL U7873 ( .A(n6258), .B(n6259), .Y(n6253) );
  MXI2X1 U7874 ( .A(U2_pipe3[7]), .B(n18057), .S0(n8054), .Y(n4213) );
  XNOR2X1 U7875 ( .A(n18098), .B(n18097), .Y(n18099) );
  AOI21X1 U7876 ( .A0(n14385), .A1(n14384), .B0(n14383), .Y(n25208) );
  XNOR2X1 U7877 ( .A(n18187), .B(n18146), .Y(n18147) );
  MXI2X1 U7878 ( .A(U0_pipe9[5]), .B(n25774), .S0(n6887), .Y(n4600) );
  AOI21X1 U7879 ( .A0(n13451), .A1(n24492), .B0(n13450), .Y(n24478) );
  MXI2X1 U7880 ( .A(U0_pipe6[5]), .B(n21926), .S0(n21972), .Y(n4485) );
  NAND2BX1 U7881 ( .AN(n14945), .B(n14953), .Y(n16842) );
  MXI2X1 U7882 ( .A(U2_pipe0[8]), .B(n26159), .S0(n8054), .Y(n4059) );
  NAND2XL U7883 ( .A(n19751), .B(U1_A_i_d0[16]), .Y(n16684) );
  XNOR2X1 U7884 ( .A(n26194), .B(n26193), .Y(n26195) );
  INVX1 U7885 ( .A(n22807), .Y(n22836) );
  NAND2X1 U7886 ( .A(n19158), .B(n19157), .Y(n19454) );
  CLKINVX3 U7887 ( .A(n14553), .Y(n13123) );
  MXI2X1 U7888 ( .A(U0_pipe3[5]), .B(n24829), .S0(n24784), .Y(n4370) );
  OR2X2 U7889 ( .A(n19751), .B(U1_A_i_d0[16]), .Y(n8574) );
  XNOR2X1 U7890 ( .A(n26289), .B(n26245), .Y(n26246) );
  MXI2X1 U7891 ( .A(U0_pipe8[8]), .B(n25618), .S0(n6888), .Y(n4426) );
  MXI2X1 U7892 ( .A(U0_pipe11[5]), .B(n23103), .S0(n24784), .Y(n4544) );
  INVX1 U7893 ( .A(n14966), .Y(n5797) );
  MXI2X1 U7894 ( .A(U0_pipe11[4]), .B(n23110), .S0(n24784), .Y(n4545) );
  INVX1 U7895 ( .A(n19639), .Y(n19662) );
  XNOR2X1 U7896 ( .A(n20901), .B(n20858), .Y(n20859) );
  INVX1 U7897 ( .A(n20007), .Y(n5867) );
  AND2XL U7898 ( .A(n21774), .B(U2_A_r_d[14]), .Y(n14442) );
  AOI21XL U7899 ( .A0(n22526), .A1(n22524), .B0(n14035), .Y(n14036) );
  INVX1 U7900 ( .A(n22687), .Y(n22705) );
  INVX1 U7901 ( .A(n25207), .Y(n25237) );
  INVX1 U7902 ( .A(n19450), .Y(n19472) );
  INVX1 U7903 ( .A(n13114), .Y(n14536) );
  INVX1 U7904 ( .A(n21881), .Y(n21908) );
  NAND3BX2 U7905 ( .AN(n9183), .B(n6356), .C(n5889), .Y(n6348) );
  MXI2X1 U7906 ( .A(U1_pipe15[4]), .B(n17429), .S0(n6887), .Y(n4783) );
  AND2XL U7907 ( .A(n21774), .B(U2_A_i_d[14]), .Y(n21775) );
  NAND2X1 U7908 ( .A(n14791), .B(n14929), .Y(n20108) );
  MXI2X1 U7909 ( .A(U2_pipe2[4]), .B(n20610), .S0(n21023), .Y(n4155) );
  INVXL U7910 ( .A(n24904), .Y(n24488) );
  INVXL U7911 ( .A(n14950), .Y(n6033) );
  NOR2X1 U7912 ( .A(n18986), .B(n6259), .Y(n6256) );
  OR2X2 U7913 ( .A(n20002), .B(n14950), .Y(n14947) );
  AND2X1 U7914 ( .A(n12378), .B(n22918), .Y(n22027) );
  INVX1 U7915 ( .A(n19872), .Y(n19904) );
  MXI2X1 U7916 ( .A(U0_pipe4[7]), .B(n22269), .S0(n22248), .Y(n4340) );
  MXI2X1 U7917 ( .A(U2_pipe3[5]), .B(n17944), .S0(n8054), .Y(n4209) );
  AND2X1 U7918 ( .A(n19985), .B(n14940), .Y(n6952) );
  MXI2X1 U7919 ( .A(U0_pipe8[7]), .B(n25624), .S0(n6888), .Y(n4427) );
  INVX1 U7920 ( .A(n25072), .Y(n25090) );
  INVXL U7921 ( .A(n17680), .Y(n12967) );
  MXI2X1 U7922 ( .A(U0_pipe8[6]), .B(n25630), .S0(n6888), .Y(n4428) );
  NAND2X1 U7923 ( .A(n14828), .B(n19544), .Y(n19286) );
  MXI2X1 U7924 ( .A(U2_pipe3[4]), .B(n17894), .S0(n8054), .Y(n4207) );
  MXI2X1 U7925 ( .A(U0_pipe4[6]), .B(n22275), .S0(n22248), .Y(n4341) );
  XNOR2X1 U7926 ( .A(n17983), .B(n17982), .Y(n17984) );
  NAND2XL U7927 ( .A(n14083), .B(n22811), .Y(n14085) );
  MXI2X1 U7928 ( .A(U2_pipe3[3]), .B(n17849), .S0(n8054), .Y(n4205) );
  XOR2XL U7929 ( .A(n20167), .B(n20166), .Y(n20168) );
  INVX1 U7930 ( .A(n25199), .Y(n21774) );
  INVX1 U7931 ( .A(n18903), .Y(n18904) );
  OR2X2 U7932 ( .A(n12886), .B(n19520), .Y(n12795) );
  NOR2XL U7933 ( .A(n7549), .B(n26817), .Y(n7548) );
  MXI2X1 U7934 ( .A(U2_pipe1[4]), .B(n23280), .S0(n23695), .Y(n4103) );
  MXI2X1 U7935 ( .A(U2_pipe1[3]), .B(n23231), .S0(n23695), .Y(n4101) );
  MXI2X1 U7936 ( .A(U2_pipe0[5]), .B(n25992), .S0(n8054), .Y(n4053) );
  AND2X2 U7937 ( .A(n7225), .B(n22690), .Y(n7042) );
  MXI2X1 U7938 ( .A(U2_pipe2[3]), .B(n20559), .S0(n21023), .Y(n4153) );
  INVX1 U7939 ( .A(n7727), .Y(n9169) );
  INVX1 U7940 ( .A(n25755), .Y(n25773) );
  MXI2X1 U7941 ( .A(U2_pipe3[2]), .B(n17796), .S0(n8054), .Y(n4203) );
  NAND2BX1 U7942 ( .AN(n7245), .B(n5874), .Y(n6782) );
  XNOR2X1 U7943 ( .A(n17795), .B(n17794), .Y(n17796) );
  NAND2XL U7944 ( .A(n14073), .B(n7080), .Y(n14083) );
  OR2X2 U7945 ( .A(n21577), .B(n21576), .Y(n21575) );
  NAND2X1 U7946 ( .A(n21618), .B(n21617), .Y(n21656) );
  INVXL U7947 ( .A(n24287), .Y(n7383) );
  MXI2X1 U7948 ( .A(U2_pipe0[4]), .B(n25948), .S0(n8054), .Y(n4257) );
  NAND2BXL U7949 ( .AN(n13153), .B(n6809), .Y(n6808) );
  NAND2X1 U7950 ( .A(n18867), .B(n18866), .Y(n18903) );
  INVX1 U7951 ( .A(n20419), .Y(n20437) );
  OR2X2 U7952 ( .A(n19970), .B(n19969), .Y(n19950) );
  AND2X2 U7953 ( .A(n13604), .B(n13614), .Y(n7028) );
  OR2X2 U7954 ( .A(n19984), .B(n19311), .Y(n19310) );
  XNOR2X1 U7955 ( .A(n17155), .B(n17154), .Y(n17156) );
  INVXL U7956 ( .A(n12222), .Y(n5874) );
  INVX1 U7957 ( .A(n17403), .Y(n17421) );
  NOR2X1 U7958 ( .A(n5937), .B(n13949), .Y(n5936) );
  XOR2X1 U7959 ( .A(n14420), .B(n14419), .Y(n25203) );
  MXI2X1 U7960 ( .A(Q4[25]), .B(n19008), .S0(U1_valid[1]), .Y(n3961) );
  MXI2X1 U7961 ( .A(Q5[25]), .B(n19015), .S0(U1_valid[1]), .Y(n4013) );
  MXI2X1 U7962 ( .A(Q6[25]), .B(n19001), .S0(U1_valid[1]), .Y(n3882) );
  NAND2XL U7963 ( .A(n6548), .B(U2_A_i_d[6]), .Y(n22559) );
  NAND2X1 U7964 ( .A(n24621), .B(n22915), .Y(n22683) );
  INVX1 U7965 ( .A(n22888), .Y(n23087) );
  NAND2X1 U7966 ( .A(n21073), .B(n21072), .Y(n21179) );
  INVX1 U7967 ( .A(n6089), .Y(n13592) );
  INVX1 U7968 ( .A(n18050), .Y(n17937) );
  NOR2X1 U7969 ( .A(n18481), .B(n18486), .Y(n18489) );
  NAND2X1 U7970 ( .A(n9150), .B(n9155), .Y(n9183) );
  INVX2 U7971 ( .A(n14791), .Y(n19986) );
  NAND2XL U7972 ( .A(n12221), .B(n12243), .Y(n12222) );
  INVXL U7973 ( .A(n24289), .Y(n18906) );
  INVXL U7974 ( .A(n24249), .Y(n18864) );
  INVX2 U7975 ( .A(n13058), .Y(n5878) );
  OR2X2 U7976 ( .A(n13606), .B(n13605), .Y(n13604) );
  NOR2X1 U7977 ( .A(n13671), .B(U1_A_r_d0[4]), .Y(n19210) );
  NAND2X1 U7978 ( .A(n18363), .B(n18362), .Y(n18485) );
  NOR2X1 U7979 ( .A(n18363), .B(n18362), .Y(n18481) );
  NAND2X1 U7980 ( .A(n13575), .B(n13574), .Y(n13600) );
  AND2X2 U7981 ( .A(n5884), .B(n13590), .Y(n6994) );
  NOR2XL U7982 ( .A(n6931), .B(n13577), .Y(n7924) );
  NAND2X1 U7983 ( .A(n13904), .B(n13921), .Y(n13905) );
  INVX1 U7984 ( .A(n13674), .Y(n9664) );
  MXI2X1 U7985 ( .A(Q1[52]), .B(n27028), .S0(n24128), .Y(n3493) );
  MXI2X1 U7986 ( .A(Q0[24]), .B(n24361), .S0(n24128), .Y(n3519) );
  NOR2X1 U7987 ( .A(n20754), .B(n20753), .Y(n20848) );
  MXI2X1 U7988 ( .A(Q0[52]), .B(n27020), .S0(n24128), .Y(n3430) );
  NAND2X1 U7989 ( .A(n20754), .B(n20753), .Y(n20850) );
  MXI2X1 U7990 ( .A(Q1[24]), .B(n24353), .S0(n23239), .Y(n3467) );
  NOR2X1 U7991 ( .A(n13671), .B(U1_A_i_d0[4]), .Y(n17278) );
  MXI2X1 U7992 ( .A(Q2[52]), .B(n27012), .S0(n24128), .Y(n3624) );
  NOR2X1 U7993 ( .A(n23873), .B(n23872), .Y(n23927) );
  MXI2X1 U7994 ( .A(Q7[52]), .B(n21667), .S0(n24128), .Y(n3907) );
  XNOR2X1 U7995 ( .A(n19696), .B(n19695), .Y(n19697) );
  MXI2X1 U7996 ( .A(Q6[52]), .B(n21675), .S0(n24128), .Y(n3855) );
  MXI2X1 U7997 ( .A(Q3[24]), .B(n24345), .S0(n24128), .Y(n3546) );
  INVX1 U7998 ( .A(n6646), .Y(n6645) );
  MXI2X1 U7999 ( .A(Q3[52]), .B(n27004), .S0(n23239), .Y(n3572) );
  MXI2X1 U8000 ( .A(Q5[52]), .B(n21691), .S0(n24128), .Y(n3986) );
  INVX1 U8001 ( .A(n14409), .Y(n14420) );
  MXI2X1 U8002 ( .A(Q2[24]), .B(n24369), .S0(n23239), .Y(n3598) );
  INVX2 U8003 ( .A(n19737), .Y(n12301) );
  AOI2BB2XL U8004 ( .B0(n14797), .B1(n7159), .A0N(n14797), .A1N(n7049), .Y(
        n7158) );
  NOR2X1 U8005 ( .A(n26463), .B(n26462), .Y(n26591) );
  INVX1 U8006 ( .A(n12781), .Y(n12773) );
  NAND2X1 U8007 ( .A(n9071), .B(n9164), .Y(n9072) );
  NOR2X1 U8008 ( .A(n18054), .B(n18053), .Y(n18136) );
  NAND2X1 U8009 ( .A(n9168), .B(n9163), .Y(n9175) );
  NAND2X1 U8010 ( .A(n12220), .B(n12219), .Y(n12243) );
  INVX2 U8011 ( .A(n9659), .Y(n13671) );
  NAND2BX1 U8012 ( .AN(n8452), .B(n6647), .Y(n6646) );
  NAND2X1 U8013 ( .A(n18256), .B(n18255), .Y(n18355) );
  OAI21XL U8014 ( .A0(n5888), .A1(n5887), .B0(n6262), .Y(n23872) );
  NAND2X1 U8015 ( .A(n23798), .B(n23797), .Y(n23926) );
  INVXL U8016 ( .A(n26242), .Y(n20903) );
  XNOR2X1 U8017 ( .A(n17439), .B(n17438), .Y(n17440) );
  NAND2X1 U8018 ( .A(n12646), .B(n13136), .Y(n6923) );
  NAND2X1 U8019 ( .A(n12632), .B(n12638), .Y(n7953) );
  XNOR2X1 U8020 ( .A(n23174), .B(n16626), .Y(n16627) );
  AOI21X1 U8021 ( .A0(n11561), .A1(n11582), .B0(n11560), .Y(n11566) );
  INVX1 U8022 ( .A(n13590), .Y(n6088) );
  INVX1 U8023 ( .A(n9521), .Y(n9523) );
  INVX1 U8024 ( .A(n13923), .Y(n6076) );
  OR2X2 U8025 ( .A(n13923), .B(n13919), .Y(n6052) );
  NAND2XL U8026 ( .A(n7521), .B(n7522), .Y(n7831) );
  OAI21X2 U8027 ( .A0(n13063), .A1(n7524), .B0(n7523), .Y(n6155) );
  AND2X2 U8028 ( .A(n13094), .B(n13579), .Y(n6931) );
  INVX1 U8029 ( .A(n13939), .Y(n7900) );
  NAND2X2 U8030 ( .A(n12975), .B(n12981), .Y(n13058) );
  AND2X2 U8031 ( .A(n14843), .B(n14842), .Y(n6974) );
  NAND2X1 U8032 ( .A(n11455), .B(n11489), .Y(n11471) );
  INVX1 U8033 ( .A(n25263), .Y(n14338) );
  OR2X2 U8034 ( .A(n13049), .B(n13050), .Y(n13071) );
  INVX1 U8035 ( .A(n25256), .Y(n21747) );
  NAND2X1 U8036 ( .A(n8976), .B(n8975), .Y(n8977) );
  INVX1 U8037 ( .A(n12637), .Y(n5886) );
  NAND2X1 U8038 ( .A(n12146), .B(n12158), .Y(n12147) );
  NAND2X1 U8039 ( .A(n8944), .B(n8980), .Y(n8945) );
  AND2X2 U8040 ( .A(n12163), .B(n12177), .Y(n6893) );
  AND2X2 U8041 ( .A(n12568), .B(n12583), .Y(n6892) );
  INVX1 U8042 ( .A(n12639), .Y(n6789) );
  INVX1 U8043 ( .A(n13099), .Y(n14515) );
  INVX1 U8044 ( .A(n8149), .Y(n6647) );
  OAI21XL U8045 ( .A0(n23870), .A1(n23871), .B0(U2_A_i_d[14]), .Y(n6262) );
  NOR2BX2 U8046 ( .AN(n7929), .B(n12980), .Y(n5949) );
  NAND2X1 U8047 ( .A(n17941), .B(n17940), .Y(n18043) );
  NOR2X1 U8048 ( .A(n23368), .B(n23367), .Y(n23470) );
  NAND2X1 U8049 ( .A(n23368), .B(n23367), .Y(n23473) );
  AND2X2 U8050 ( .A(n13787), .B(n13793), .Y(n6993) );
  INVX1 U8051 ( .A(n12295), .Y(n19723) );
  INVX1 U8052 ( .A(n13670), .Y(n9658) );
  INVX1 U8053 ( .A(n9330), .Y(n7684) );
  NOR2X1 U8054 ( .A(n20606), .B(n20605), .Y(n20648) );
  NAND2X1 U8055 ( .A(n9331), .B(n9330), .Y(n9483) );
  NAND2X1 U8056 ( .A(n13587), .B(n13586), .Y(n13590) );
  NOR2X1 U8057 ( .A(n13641), .B(n13640), .Y(n13653) );
  NAND2X1 U8058 ( .A(n13630), .B(n13629), .Y(n13637) );
  NAND2X1 U8059 ( .A(n14683), .B(n14682), .Y(n14849) );
  NOR2X1 U8060 ( .A(n14686), .B(n14685), .Y(n14858) );
  INVX1 U8061 ( .A(n8568), .Y(n8565) );
  XOR2X1 U8062 ( .A(U1_U1_y0[40]), .B(U1_U1_y2[40]), .Y(n13656) );
  NAND2XL U8063 ( .A(n9205), .B(n9204), .Y(n9219) );
  INVX1 U8064 ( .A(n9128), .Y(n6322) );
  NAND2X1 U8065 ( .A(n5899), .B(n8531), .Y(n8532) );
  INVX1 U8066 ( .A(n13031), .Y(n5896) );
  OR2X2 U8067 ( .A(n9192), .B(n9191), .Y(n9190) );
  INVX1 U8068 ( .A(n25269), .Y(n21742) );
  NAND2X1 U8069 ( .A(n13386), .B(n13385), .Y(n13387) );
  NAND2X1 U8070 ( .A(n13143), .B(n13142), .Y(n13149) );
  NAND2X1 U8071 ( .A(n13067), .B(n13066), .Y(n13079) );
  INVX1 U8072 ( .A(n25275), .Y(n21739) );
  INVXL U8073 ( .A(U2_U0_y2[36]), .Y(n6411) );
  NOR2X2 U8074 ( .A(n14673), .B(n14672), .Y(n14794) );
  OR2XL U8075 ( .A(n14908), .B(n14907), .Y(n14906) );
  NAND2X1 U8076 ( .A(n14669), .B(n14668), .Y(n14802) );
  OR2XL U8077 ( .A(n19711), .B(U1_A_r_d0[1]), .Y(n19710) );
  NOR2X1 U8078 ( .A(n12891), .B(n7827), .Y(n7825) );
  NOR2X1 U8079 ( .A(n23324), .B(n23323), .Y(n23363) );
  NOR2X1 U8080 ( .A(n17792), .B(n17791), .Y(n17840) );
  NAND2BX2 U8081 ( .AN(n13853), .B(n6056), .Y(n13860) );
  NOR2X1 U8082 ( .A(n13183), .B(n13182), .Y(n13187) );
  NAND2X1 U8083 ( .A(n11492), .B(n11491), .Y(n11493) );
  INVX1 U8084 ( .A(n12344), .Y(n5893) );
  NAND2X1 U8085 ( .A(n5900), .B(n8582), .Y(n8583) );
  XOR2X1 U8086 ( .A(U1_U1_y0[40]), .B(U1_U1_y1[40]), .Y(n14688) );
  OR2XL U8087 ( .A(n14908), .B(n19954), .Y(n19953) );
  INVX1 U8088 ( .A(n12291), .Y(n19717) );
  NAND2X1 U8089 ( .A(n13285), .B(n13474), .Y(n13475) );
  NAND2X1 U8090 ( .A(n14676), .B(n14675), .Y(n14842) );
  NOR2X1 U8091 ( .A(n9069), .B(n9070), .Y(n9166) );
  NAND2X1 U8092 ( .A(n9070), .B(n9069), .Y(n9164) );
  NOR2X1 U8093 ( .A(n25988), .B(n25987), .Y(n26033) );
  OR2X2 U8094 ( .A(n12861), .B(n19373), .Y(n12860) );
  NAND2X1 U8095 ( .A(n9171), .B(n9170), .Y(n9177) );
  INVX1 U8096 ( .A(n23634), .Y(n18254) );
  NAND2X1 U8097 ( .A(n13897), .B(n5934), .Y(n13914) );
  NOR2X1 U8098 ( .A(n20510), .B(n20509), .Y(n20550) );
  NAND2X1 U8099 ( .A(n9229), .B(n9228), .Y(n12343) );
  INVX1 U8100 ( .A(n8536), .Y(n8538) );
  AND2X2 U8101 ( .A(n14764), .B(n14763), .Y(n14765) );
  NAND2X1 U8102 ( .A(n14353), .B(n14352), .Y(n14354) );
  NOR2X2 U8103 ( .A(n8943), .B(n8942), .Y(n8982) );
  NAND2X1 U8104 ( .A(n8933), .B(n8932), .Y(n8975) );
  NOR2X1 U8105 ( .A(n25890), .B(n25889), .Y(n25939) );
  AND2X2 U8106 ( .A(U1_U0_y1[29]), .B(U1_U0_y0[29]), .Y(n7029) );
  NOR2X2 U8107 ( .A(n12920), .B(n12922), .Y(n7930) );
  INVX1 U8108 ( .A(n12938), .Y(n12896) );
  INVX1 U8109 ( .A(n12939), .Y(n7933) );
  NOR2X1 U8110 ( .A(n12472), .B(n12475), .Y(n12530) );
  NAND2X1 U8111 ( .A(n8996), .B(n8995), .Y(n9014) );
  INVX1 U8112 ( .A(n8821), .Y(n5901) );
  INVX1 U8113 ( .A(n13409), .Y(n13411) );
  OAI21XL U8114 ( .A0(n12813), .A1(n12822), .B0(n12814), .Y(n7173) );
  INVX1 U8115 ( .A(n14758), .Y(n14764) );
  INVX1 U8116 ( .A(U1_U1_y0[32]), .Y(n6136) );
  INVX2 U8117 ( .A(n9350), .Y(n9403) );
  NOR2X2 U8118 ( .A(n12892), .B(n6709), .Y(n12922) );
  NOR2X1 U8119 ( .A(n12895), .B(n12894), .Y(n12936) );
  NAND2X2 U8120 ( .A(n12895), .B(n12894), .Y(n12938) );
  NAND2X1 U8121 ( .A(n13268), .B(n13267), .Y(n13417) );
  NAND2X1 U8122 ( .A(n11452), .B(n7118), .Y(n11491) );
  NAND2X1 U8123 ( .A(n11451), .B(U2_B_r[21]), .Y(n11498) );
  BUFX4 U8124 ( .A(n11623), .Y(n29093) );
  BUFX4 U8125 ( .A(n11615), .Y(n29108) );
  NOR2X2 U8126 ( .A(n12467), .B(n12466), .Y(n12475) );
  NAND2X1 U8127 ( .A(n8893), .B(n6368), .Y(n8948) );
  INVX1 U8128 ( .A(n12092), .Y(n12099) );
  BUFX12 U8129 ( .A(n27560), .Y(n28579) );
  BUFX4 U8130 ( .A(n11635), .Y(n29096) );
  INVX1 U8131 ( .A(n11579), .Y(n11574) );
  NOR2X1 U8132 ( .A(n8840), .B(n8851), .Y(n8893) );
  BUFX12 U8133 ( .A(n28168), .Y(n28125) );
  NAND2X1 U8134 ( .A(n8478), .B(n6592), .Y(n8463) );
  INVX1 U8135 ( .A(U0_U2_y0[24]), .Y(n6742) );
  INVX1 U8136 ( .A(n8898), .Y(n8918) );
  INVX1 U8137 ( .A(n11531), .Y(n11519) );
  NOR2X1 U8138 ( .A(n12465), .B(n12464), .Y(n12472) );
  NAND2X1 U8139 ( .A(n8314), .B(n11583), .Y(n8315) );
  BUFX8 U8140 ( .A(n28186), .Y(n28237) );
  NAND2X1 U8141 ( .A(n14649), .B(n14648), .Y(n14770) );
  INVX1 U8142 ( .A(n18722), .Y(n18660) );
  AOI2BB1X1 U8143 ( .A0N(n9385), .A1N(n9389), .B0(n6514), .Y(n6513) );
  NAND2BXL U8144 ( .AN(n9289), .B(n5919), .Y(n6512) );
  INVX1 U8145 ( .A(n9367), .Y(n9368) );
  NAND2X1 U8146 ( .A(n12758), .B(n12757), .Y(n12875) );
  INVX1 U8147 ( .A(n26785), .Y(n26746) );
  INVX1 U8148 ( .A(n26773), .Y(n26713) );
  INVX1 U8149 ( .A(n21471), .Y(n21406) );
  INVX1 U8150 ( .A(n24111), .Y(n24051) );
  NAND2X4 U8151 ( .A(n5826), .B(n28675), .Y(n27379) );
  INVX1 U8152 ( .A(n6371), .Y(n6370) );
  INVX1 U8153 ( .A(n21435), .Y(n21373) );
  INVX1 U8154 ( .A(n21447), .Y(n21384) );
  BUFX4 U8155 ( .A(n11627), .Y(n29095) );
  INVX1 U8156 ( .A(n26809), .Y(n26724) );
  NAND2X2 U8157 ( .A(C_sel_reg[1]), .B(n28252), .Y(n28054) );
  CLKINVX3 U8158 ( .A(n5829), .Y(n12000) );
  NAND2X1 U8159 ( .A(n8805), .B(n8804), .Y(n8921) );
  INVX1 U8160 ( .A(n23892), .Y(n23649) );
  BUFX12 U8161 ( .A(U1_U1_z2[3]), .Y(n6877) );
  NAND2X1 U8162 ( .A(n12457), .B(n12456), .Y(n12483) );
  AOI21X1 U8163 ( .A0(n8734), .A1(n8733), .B0(n7970), .Y(n8865) );
  NAND2X1 U8164 ( .A(n12459), .B(n12458), .Y(n12523) );
  NOR2X1 U8165 ( .A(n12459), .B(n12458), .Y(n12516) );
  CLKINVX3 U8166 ( .A(U2_B_i[5]), .Y(n9623) );
  INVX1 U8167 ( .A(U2_U0_y1[13]), .Y(n20468) );
  CLKINVX2 U8168 ( .A(n11940), .Y(n5918) );
  INVX1 U8169 ( .A(n18514), .Y(n18267) );
  BUFX12 U8170 ( .A(n27686), .Y(n28353) );
  INVX8 U8171 ( .A(n15003), .Y(n5826) );
  NAND2X1 U8172 ( .A(n12697), .B(n12696), .Y(n12867) );
  AOI21X1 U8173 ( .A0(n27976), .A1(Q1[10]), .B0(n27856), .Y(n28360) );
  CLKINVX2 U8174 ( .A(n11940), .Y(n5798) );
  OR2X2 U8175 ( .A(n12831), .B(n12836), .Y(n6169) );
  INVX2 U8176 ( .A(n11612), .Y(n11998) );
  NOR2X1 U8177 ( .A(n14978), .B(n7305), .Y(n11908) );
  OAI21XL U8178 ( .A0(n7300), .A1(n28673), .B0(n7298), .Y(n11911) );
  NOR2X1 U8179 ( .A(n14721), .B(n14726), .Y(n14633) );
  INVXL U8180 ( .A(n25101), .Y(n6532) );
  AND2X2 U8181 ( .A(B_sel_reg[0]), .B(n28322), .Y(n11891) );
  AOI21X1 U8182 ( .A0(n10782), .A1(n10792), .B0(n10781), .Y(n10783) );
  CLKINVX8 U8183 ( .A(n16375), .Y(n5799) );
  NAND2X1 U8184 ( .A(n9852), .B(n9851), .Y(n10191) );
  INVX4 U8185 ( .A(n5924), .Y(n5800) );
  NOR2X1 U8186 ( .A(n12750), .B(U1_U2_y1[13]), .Y(n12851) );
  BUFX3 U8187 ( .A(n10126), .Y(n10127) );
  BUFX2 U8188 ( .A(n10055), .Y(n10056) );
  NAND2X1 U8189 ( .A(n9287), .B(U1_U0_y1[13]), .Y(n9390) );
  INVX8 U8190 ( .A(n11719), .Y(n5801) );
  INVX1 U8191 ( .A(n9927), .Y(n9876) );
  CLKINVX3 U8192 ( .A(n9869), .Y(n5923) );
  INVX8 U8193 ( .A(n11677), .Y(n5802) );
  INVX8 U8194 ( .A(n11679), .Y(n5803) );
  INVXL U8195 ( .A(n6394), .Y(n6400) );
  NAND2X1 U8196 ( .A(n6395), .B(n6394), .Y(n6393) );
  CLKINVX8 U8197 ( .A(n7096), .Y(n5804) );
  INVX1 U8198 ( .A(n10905), .Y(n10897) );
  INVX1 U8199 ( .A(n11261), .Y(n11253) );
  NOR2X1 U8200 ( .A(n11080), .B(n8294), .Y(n11208) );
  NAND2X2 U8201 ( .A(n10405), .B(n6429), .Y(n10397) );
  INVX4 U8202 ( .A(n5837), .Y(n5920) );
  NAND2X1 U8203 ( .A(n6654), .B(U1_U0_y2[13]), .Y(n8399) );
  NAND2X1 U8204 ( .A(n28960), .B(n5840), .Y(n27143) );
  NAND2X1 U8205 ( .A(n28961), .B(n5927), .Y(n27147) );
  NAND2X1 U8206 ( .A(n28962), .B(n5927), .Y(n27151) );
  NAND2X1 U8207 ( .A(n28965), .B(n5840), .Y(n27164) );
  NAND2X1 U8208 ( .A(n28966), .B(n5840), .Y(n27168) );
  NAND2X1 U8209 ( .A(n28970), .B(n5840), .Y(n27220) );
  NAND2X1 U8210 ( .A(n28971), .B(n5840), .Y(n27224) );
  NAND2X1 U8211 ( .A(n28972), .B(n5840), .Y(n27228) );
  NAND2X1 U8212 ( .A(n28958), .B(n5840), .Y(n27135) );
  NAND2X1 U8213 ( .A(n28959), .B(n5840), .Y(n27139) );
  INVX4 U8214 ( .A(n5837), .Y(n5805) );
  INVX1 U8215 ( .A(n22248), .Y(n5838) );
  NAND2X1 U8216 ( .A(n28974), .B(n5927), .Y(n27237) );
  NAND2X1 U8217 ( .A(n28975), .B(n5927), .Y(n27241) );
  NAND2X1 U8218 ( .A(n28977), .B(n5840), .Y(n27249) );
  NAND2X1 U8219 ( .A(n28978), .B(n5840), .Y(n27253) );
  NAND2X1 U8220 ( .A(n28979), .B(n5840), .Y(n27257) );
  NAND2X1 U8221 ( .A(n28980), .B(n5840), .Y(n27261) );
  NAND2X1 U8222 ( .A(n28981), .B(n5840), .Y(n27266) );
  NAND2X1 U8223 ( .A(n28982), .B(n5840), .Y(n27270) );
  NAND2X1 U8224 ( .A(n11354), .B(n11353), .Y(n11355) );
  NAND2X1 U8225 ( .A(n10579), .B(n9561), .Y(n10565) );
  NAND2X1 U8226 ( .A(n10443), .B(n10442), .Y(n10444) );
  NAND2X1 U8227 ( .A(n10449), .B(n10448), .Y(n10450) );
  NAND2X1 U8228 ( .A(n10423), .B(n10422), .Y(n10424) );
  AND2X2 U8229 ( .A(n9239), .B(n10754), .Y(n7002) );
  NAND2X1 U8230 ( .A(BOPA[24]), .B(n11430), .Y(n11424) );
  OAI32X1 U8231 ( .A0(n7305), .A1(C_sel_reg[8]), .A2(A_sel_reg[4]), .B0(n14994), .B1(n11633), .Y(n16416) );
  NAND2X1 U8232 ( .A(n11276), .B(n8345), .Y(n11262) );
  NAND2X1 U8233 ( .A(n10247), .B(n10252), .Y(n10208) );
  NAND2X1 U8234 ( .A(n10951), .B(n10950), .Y(n10952) );
  INVX4 U8235 ( .A(n15633), .Y(n5926) );
  CLKBUFX8 U8236 ( .A(n15969), .Y(n5925) );
  INVX8 U8237 ( .A(n15179), .Y(n5836) );
  CLKINVX3 U8238 ( .A(n15495), .Y(n16161) );
  NAND2X1 U8239 ( .A(n10355), .B(n8233), .Y(n8235) );
  NAND2X1 U8240 ( .A(n10406), .B(n10405), .Y(n10407) );
  NAND2X1 U8241 ( .A(n9791), .B(n9790), .Y(n10039) );
  NAND2X1 U8242 ( .A(n9940), .B(n9939), .Y(n10332) );
  AND2X1 U8243 ( .A(n10701), .B(n10848), .Y(n10702) );
  NAND2BX2 U8244 ( .AN(n10404), .B(n6425), .Y(n6429) );
  INVX1 U8245 ( .A(n9763), .Y(n9796) );
  NAND2X1 U8246 ( .A(n10466), .B(n10465), .Y(n10467) );
  INVX1 U8247 ( .A(n10779), .Y(n10792) );
  OR2XL U8248 ( .A(n18696), .B(n18695), .Y(n18694) );
  OR2XL U8249 ( .A(n21438), .B(n21437), .Y(n21436) );
  INVX1 U8250 ( .A(n10370), .Y(n10384) );
  AOI21X1 U8251 ( .A0(n14603), .A1(n14602), .B0(n14601), .Y(n14609) );
  OR2XL U8252 ( .A(n18587), .B(n18586), .Y(n18585) );
  OR2XL U8253 ( .A(n21541), .B(n21540), .Y(n21539) );
  OR2XL U8254 ( .A(n21627), .B(n21626), .Y(n21625) );
  OR2XL U8255 ( .A(n26738), .B(n26737), .Y(n26736) );
  OR2XL U8256 ( .A(n18663), .B(n18662), .Y(n18661) );
  OR2XL U8257 ( .A(n26983), .B(n26982), .Y(n26981) );
  NOR2X1 U8258 ( .A(n10691), .B(n10693), .Y(n10722) );
  INVX8 U8259 ( .A(n15967), .Y(n15982) );
  OR2XL U8260 ( .A(n18940), .B(n18939), .Y(n18938) );
  OR2XL U8261 ( .A(n26885), .B(n26884), .Y(n26883) );
  NAND2X1 U8262 ( .A(n11418), .B(BOPA[14]), .Y(n9240) );
  INVX8 U8263 ( .A(n5931), .Y(n5806) );
  INVXL U8264 ( .A(n9799), .Y(n9801) );
  OR2XL U8265 ( .A(n18762), .B(n18761), .Y(n18760) );
  INVX1 U8266 ( .A(n10387), .Y(n10401) );
  OR2XL U8267 ( .A(n26632), .B(n26631), .Y(n26630) );
  OR2XL U8268 ( .A(n18853), .B(n18852), .Y(n18851) );
  INVX1 U8269 ( .A(n9856), .Y(n9858) );
  CLKINVX3 U8270 ( .A(n15218), .Y(n15179) );
  INVX2 U8271 ( .A(n15214), .Y(n15948) );
  INVX1 U8272 ( .A(n27942), .Y(n27943) );
  NOR2X1 U8273 ( .A(n10553), .B(n10559), .Y(n10548) );
  BUFX12 U8274 ( .A(n25330), .Y(n20240) );
  OR2XL U8275 ( .A(n26975), .B(n26974), .Y(n26973) );
  OR2XL U8276 ( .A(n18829), .B(n18828), .Y(n18827) );
  OR2XL U8277 ( .A(n24308), .B(n24307), .Y(n24306) );
  OR2XL U8278 ( .A(n21635), .B(n21634), .Y(n21633) );
  INVX1 U8279 ( .A(n9764), .Y(n9766) );
  INVX1 U8280 ( .A(n9742), .Y(n9744) );
  OR2XL U8281 ( .A(n18725), .B(n18724), .Y(n18723) );
  OR2XL U8282 ( .A(n18557), .B(n18556), .Y(n18555) );
  OR2XL U8283 ( .A(n18517), .B(n18516), .Y(n18515) );
  OR2XL U8284 ( .A(n21300), .B(n21299), .Y(n21298) );
  OR2XL U8285 ( .A(n21233), .B(n21232), .Y(n21231) );
  OR2XL U8286 ( .A(n18916), .B(n18915), .Y(n18914) );
  OR2XL U8287 ( .A(n23975), .B(n23974), .Y(n23973) );
  OR2XL U8288 ( .A(n18845), .B(n18844), .Y(n18843) );
  OR2XL U8289 ( .A(n21213), .B(n21212), .Y(n21211) );
  OR2XL U8290 ( .A(n21276), .B(n21275), .Y(n21274) );
  OR2XL U8291 ( .A(n18932), .B(n18931), .Y(n18930) );
  OR2XL U8292 ( .A(n21376), .B(n21375), .Y(n21374) );
  OR2XL U8293 ( .A(n26800), .B(n26799), .Y(n26798) );
  CLKBUFX8 U8294 ( .A(n25330), .Y(n22248) );
  OR2XL U8295 ( .A(n18577), .B(n18576), .Y(n18575) );
  OR2XL U8296 ( .A(n24241), .B(n24240), .Y(n24239) );
  OR2XL U8297 ( .A(n21565), .B(n21564), .Y(n21563) );
  CLKINVX8 U8298 ( .A(n11628), .Y(n5808) );
  OR2XL U8299 ( .A(n18685), .B(n18684), .Y(n18683) );
  INVX1 U8300 ( .A(n10737), .Y(n10751) );
  OR2XL U8301 ( .A(n21450), .B(n21449), .Y(n21448) );
  OR2XL U8302 ( .A(n24126), .B(n24125), .Y(n24124) );
  OR2XL U8303 ( .A(n21387), .B(n21386), .Y(n21385) );
  OR2XL U8304 ( .A(n26893), .B(n26892), .Y(n26891) );
  CLKINVX8 U8305 ( .A(n17249), .Y(n5809) );
  OR2XL U8306 ( .A(n18750), .B(n18749), .Y(n18748) );
  OR2XL U8307 ( .A(n24087), .B(n24086), .Y(n24085) );
  NOR2X1 U8308 ( .A(n10911), .B(n10915), .Y(n8328) );
  OR2XL U8309 ( .A(n26812), .B(n26811), .Y(n26810) );
  OR2XL U8310 ( .A(n21293), .B(n21292), .Y(n21291) );
  OR2XL U8311 ( .A(n26727), .B(n26726), .Y(n26725) );
  OR2XL U8312 ( .A(n26639), .B(n26638), .Y(n26637) );
  OR2XL U8313 ( .A(n21398), .B(n21397), .Y(n21396) );
  OR2XL U8314 ( .A(n26560), .B(n26559), .Y(n26558) );
  OR2XL U8315 ( .A(n21462), .B(n21461), .Y(n21460) );
  INVX1 U8316 ( .A(n10621), .Y(n10631) );
  CLKINVX3 U8317 ( .A(n25330), .Y(n17032) );
  OR2XL U8318 ( .A(n26967), .B(n26966), .Y(n26965) );
  OR2XL U8319 ( .A(n26901), .B(n26900), .Y(n26899) );
  OR2XL U8320 ( .A(n24139), .B(n24138), .Y(n24137) );
  OR2XL U8321 ( .A(n24233), .B(n24232), .Y(n24231) );
  AOI21XL U8322 ( .A0(n8362), .A1(n8361), .B0(n8360), .Y(n8369) );
  OR2XL U8323 ( .A(n24316), .B(n24315), .Y(n24314) );
  INVXL U8324 ( .A(U1_U0_y0[13]), .Y(n6654) );
  OR2XL U8325 ( .A(n21557), .B(n21556), .Y(n21555) );
  OR2XL U8326 ( .A(n21643), .B(n21642), .Y(n21641) );
  INVX1 U8327 ( .A(n10146), .Y(n10149) );
  OR2XL U8328 ( .A(n23965), .B(n23964), .Y(n23963) );
  OR2XL U8329 ( .A(n24076), .B(n24075), .Y(n24074) );
  OR2XL U8330 ( .A(n21651), .B(n21650), .Y(n21649) );
  OR2XL U8331 ( .A(n18924), .B(n18923), .Y(n18922) );
  INVX1 U8332 ( .A(n10670), .Y(n10530) );
  OR2XL U8333 ( .A(n18837), .B(n18836), .Y(n18835) );
  OR2XL U8334 ( .A(n18737), .B(n18736), .Y(n18735) );
  OR2XL U8335 ( .A(n18674), .B(n18673), .Y(n18672) );
  OR2XL U8336 ( .A(n26776), .B(n26775), .Y(n26774) );
  OR2XL U8337 ( .A(n26716), .B(n26715), .Y(n26714) );
  OR2XL U8338 ( .A(n26877), .B(n26876), .Y(n26875) );
  NOR2X1 U8339 ( .A(n11087), .B(n11096), .Y(n6222) );
  OR2XL U8340 ( .A(n26615), .B(n26614), .Y(n26613) );
  OR2XL U8341 ( .A(n26540), .B(n26539), .Y(n26538) );
  OR2XL U8342 ( .A(n26959), .B(n26958), .Y(n26957) );
  INVX8 U8343 ( .A(n27211), .Y(n5840) );
  INVX1 U8344 ( .A(n11083), .Y(n11097) );
  INVX1 U8345 ( .A(n11379), .Y(n11237) );
  OR2XL U8346 ( .A(n24054), .B(n24053), .Y(n24052) );
  OR2XL U8347 ( .A(n24114), .B(n24113), .Y(n24112) );
  OR2XL U8348 ( .A(n24151), .B(n24150), .Y(n24149) );
  OR2XL U8349 ( .A(n24065), .B(n24064), .Y(n24063) );
  OR2XL U8350 ( .A(n23955), .B(n23954), .Y(n23953) );
  OR2XL U8351 ( .A(n24217), .B(n24216), .Y(n24215) );
  OR2XL U8352 ( .A(n24300), .B(n24299), .Y(n24298) );
  INVX1 U8353 ( .A(n10553), .Y(n10567) );
  OR2XL U8354 ( .A(n18567), .B(n18566), .Y(n18565) );
  OR2XL U8355 ( .A(n24324), .B(n24323), .Y(n24322) );
  OR2XL U8356 ( .A(n23895), .B(n23894), .Y(n23893) );
  OR2XL U8357 ( .A(n23945), .B(n23944), .Y(n23943) );
  OR2XL U8358 ( .A(n24225), .B(n24224), .Y(n24223) );
  INVX1 U8359 ( .A(n11020), .Y(n10881) );
  OR2XL U8360 ( .A(n26588), .B(n26587), .Y(n26586) );
  OR2XL U8361 ( .A(n21283), .B(n21282), .Y(n21281) );
  OR2XL U8362 ( .A(n21261), .B(n21260), .Y(n21259) );
  BUFX12 U8363 ( .A(n25330), .Y(n24784) );
  INVX8 U8364 ( .A(n5928), .Y(n5810) );
  INVX1 U8365 ( .A(n10866), .Y(n10908) );
  INVX1 U8366 ( .A(n9778), .Y(n9808) );
  OR2XL U8367 ( .A(n26622), .B(n26621), .Y(n26620) );
  OR2XL U8368 ( .A(n26749), .B(n26748), .Y(n26747) );
  OR2XL U8369 ( .A(n26788), .B(n26787), .Y(n26786) );
  NOR2X1 U8370 ( .A(n9780), .B(n9778), .Y(n6394) );
  INVX1 U8371 ( .A(n20025), .Y(n5811) );
  OR2XL U8372 ( .A(n21409), .B(n21408), .Y(n21407) );
  INVX1 U8373 ( .A(n9807), .Y(n9779) );
  OR2XL U8374 ( .A(n21474), .B(n21473), .Y(n21472) );
  OR2XL U8375 ( .A(n21549), .B(n21548), .Y(n21547) );
  INVX4 U8376 ( .A(OP_done1), .Y(n27211) );
  NAND2X1 U8377 ( .A(n8178), .B(BOPD[42]), .Y(n10754) );
  ADDHXL U8378 ( .A(U0_pipe12[20]), .B(n28793), .CO(n26776), .S(n26715) );
  NOR2X1 U8379 ( .A(n8154), .B(BOPC[49]), .Y(n11055) );
  INVX1 U8380 ( .A(B0_q[25]), .Y(n16468) );
  ADDHXL U8381 ( .A(U1_pipe2[16]), .B(n28845), .CO(n21233), .S(n21169) );
  ADDHXL U8382 ( .A(U1_pipe11[19]), .B(U1_pipe10[19]), .CO(n18674), .S(n18643)
         );
  ADDHXL U8383 ( .A(U0_pipe11[24]), .B(U0_pipe10[24]), .CO(n24308), .S(n24281)
         );
  OR2XL U8384 ( .A(U1_U1_y1[5]), .B(U1_U1_y0[5]), .Y(n14603) );
  OR2XL U8385 ( .A(U0_U2_y1[10]), .B(U0_U2_y0[10]), .Y(n8721) );
  ADDHXL U8386 ( .A(U0_pipe12[22]), .B(n28934), .CO(n26877), .S(n26830) );
  ADDHXL U8387 ( .A(U0_pipe12[19]), .B(n28794), .CO(n26716), .S(n26658) );
  ADDHXL U8388 ( .A(U1_pipe11[22]), .B(U1_pipe10[22]), .CO(n18837), .S(n18801)
         );
  OR2XL U8389 ( .A(U0_U0_y1[8]), .B(U0_U0_y0[8]), .Y(n13222) );
  ADDHXL U8390 ( .A(U1_pipe11[24]), .B(U1_pipe10[24]), .CO(n18924), .S(n18881)
         );
  ADDHXL U8391 ( .A(U1_pipe11[20]), .B(U1_pipe10[20]), .CO(n18737), .S(n18673)
         );
  ADDHXL U8392 ( .A(U1_pipe1[19]), .B(U1_pipe0[19]), .CO(n21398), .S(n21343)
         );
  OR2X2 U8393 ( .A(U1_U2_y2[11]), .B(U1_U2_y0[11]), .Y(n13762) );
  ADDHXL U8394 ( .A(U0_pipe12[17]), .B(n28796), .CO(n26615), .S(n26539) );
  BUFX12 U8395 ( .A(n25330), .Y(n5812) );
  INVX8 U8396 ( .A(n15747), .Y(n5813) );
  ADDHXL U8397 ( .A(U0_pipe12[16]), .B(n28797), .CO(n26540), .S(n26469) );
  ADDHXL U8398 ( .A(U0_pipe12[24]), .B(n28932), .CO(n26959), .S(n26917) );
  NOR2X1 U8399 ( .A(n8155), .B(BOPD[49]), .Y(n10715) );
  NAND2X1 U8400 ( .A(n8201), .B(AOPD[37]), .Y(n10975) );
  OR2XL U8401 ( .A(U1_U0_y2[12]), .B(U1_U0_y0[12]), .Y(n8385) );
  ADDHXL U8402 ( .A(U1_pipe5[24]), .B(U1_pipe4[24]), .CO(n18932), .S(n18889)
         );
  ADDHXL U8403 ( .A(U0_pipe2[19]), .B(n28778), .CO(n26727), .S(n26692) );
  NOR2X1 U8404 ( .A(n8100), .B(AOPD[46]), .Y(n10866) );
  ADDHXL U8405 ( .A(U0_pipe2[20]), .B(n28777), .CO(n26812), .S(n26726) );
  NOR2X1 U8406 ( .A(n7054), .B(AOPD[40]), .Y(n10949) );
  ADDHXL U8407 ( .A(U0_pipe2[22]), .B(n28930), .CO(n26901), .S(n26854) );
  NOR2X1 U8408 ( .A(n8091), .B(AOPD[49]), .Y(n10890) );
  ADDHXL U8409 ( .A(U0_pipe2[24]), .B(n28928), .CO(n26967), .S(n26941) );
  ADDHXL U8410 ( .A(U0_pipe2[17]), .B(n28780), .CO(n26639), .S(n26559) );
  ADDHXL U8411 ( .A(U1_pipe5[19]), .B(U1_pipe4[19]), .CO(n18685), .S(n18631)
         );
  OR2XL U8412 ( .A(U1_U1_y1[8]), .B(U1_U1_y0[8]), .Y(n14614) );
  NAND2X1 U8413 ( .A(W0[14]), .B(W0[30]), .Y(n9865) );
  NAND2X1 U8414 ( .A(n8169), .B(BOPB[45]), .Y(n10575) );
  ADDHXL U8415 ( .A(U0_pipe1[24]), .B(U0_pipe0[24]), .CO(n26975), .S(n26933)
         );
  ADDHXL U8416 ( .A(U0_pipe7[22]), .B(U0_pipe6[22]), .CO(n24225), .S(n24178)
         );
  ADDHXL U8417 ( .A(U0_pipe7[20]), .B(U0_pipe6[20]), .CO(n24151), .S(n24064)
         );
  ADDHXL U8418 ( .A(U0_pipe7[19]), .B(U0_pipe6[19]), .CO(n24065), .S(n24030)
         );
  ADDHXL U8419 ( .A(U0_pipe1[19]), .B(U0_pipe0[19]), .CO(n26738), .S(n26681)
         );
  ADDHXL U8420 ( .A(U1_pipe5[20]), .B(U1_pipe4[20]), .CO(n18750), .S(n18684)
         );
  INVX1 U8421 ( .A(B0_q[35]), .Y(n16427) );
  ADDHXL U8422 ( .A(U0_pipe1[20]), .B(U0_pipe0[20]), .CO(n26800), .S(n26737)
         );
  OR2X2 U8423 ( .A(U1_U1_y2[11]), .B(U1_U1_y0[11]), .Y(n12682) );
  OR2XL U8424 ( .A(U1_U1_y2[10]), .B(U1_U1_y0[10]), .Y(n7979) );
  ADDHXL U8425 ( .A(U0_pipe1[22]), .B(U0_pipe0[22]), .CO(n26893), .S(n26846)
         );
  OR2X2 U8426 ( .A(U1_U1_y2[9]), .B(U1_U1_y0[9]), .Y(n12681) );
  NAND2X2 U8427 ( .A(W3[0]), .B(W3[16]), .Y(n9777) );
  ADDHXL U8428 ( .A(U0_pipe7[24]), .B(U0_pipe6[24]), .CO(n24324), .S(n24265)
         );
  OR2XL U8429 ( .A(U1_U1_y2[8]), .B(U1_U1_y0[8]), .Y(n12680) );
  ADDHXL U8430 ( .A(U1_pipe5[22]), .B(U1_pipe4[22]), .CO(n18845), .S(n18793)
         );
  NAND2X1 U8431 ( .A(n7054), .B(AOPD[40]), .Y(n10950) );
  ADDHXL U8432 ( .A(U1_pipe7[19]), .B(U1_pipe6[19]), .CO(n18696), .S(n18619)
         );
  ADDHXL U8433 ( .A(U1_pipe12[17]), .B(n28860), .CO(n21276), .S(n21212) );
  ADDHXL U8434 ( .A(U1_pipe12[19]), .B(n28858), .CO(n21376), .S(n21320) );
  ADDHXL U8435 ( .A(U1_pipe8[17]), .B(n28828), .CO(n21283), .S(n21260) );
  ADDHXL U8436 ( .A(U1_pipe7[22]), .B(U1_pipe6[22]), .CO(n18853), .S(n18785)
         );
  ADDHXL U8437 ( .A(U1_pipe14[22]), .B(n28954), .CO(n18829), .S(n18777) );
  ADDHXL U8438 ( .A(U1_pipe7[20]), .B(U1_pipe6[20]), .CO(n18762), .S(n18695)
         );
  ADDHXL U8439 ( .A(U1_pipe12[16]), .B(n28861), .CO(n21213), .S(n21132) );
  ADDHXL U8440 ( .A(U1_pipe12[24]), .B(n28948), .CO(n21627), .S(n21583) );
  ADDHXL U8441 ( .A(U0_pipe14[22]), .B(n28938), .CO(n24217), .S(n24170) );
  ADDHXL U8442 ( .A(U1_pipe12[20]), .B(n28857), .CO(n21438), .S(n21375) );
  NAND2X1 U8443 ( .A(n7056), .B(AOPC[33]), .Y(n11353) );
  NAND2X1 U8444 ( .A(n8113), .B(AOPB[43]), .Y(n10405) );
  NOR2X1 U8445 ( .A(n8090), .B(AOPC[49]), .Y(n11246) );
  ADDHXL U8446 ( .A(U1_pipe14[24]), .B(n28952), .CO(n18916), .S(n18873) );
  ADDHXL U8447 ( .A(U1_pipe12[22]), .B(n28950), .CO(n21541), .S(n21489) );
  ADDHXL U8448 ( .A(U0_pipe14[24]), .B(n28936), .CO(n24300), .S(n24257) );
  AND2X2 U8449 ( .A(n7975), .B(W0[30]), .Y(n7981) );
  ADDHXL U8450 ( .A(U1_pipe14[16]), .B(n28877), .CO(n18517), .S(n18418) );
  ADDHXL U8451 ( .A(U0_pipe8[20]), .B(n28761), .CO(n26788), .S(n26748) );
  ADDHXL U8452 ( .A(U0_pipe8[17]), .B(n28764), .CO(n26622), .S(n26587) );
  ADDHXL U8453 ( .A(U0_pipe8[16]), .B(n28765), .CO(n26588), .S(n26506) );
  ADDHXL U8454 ( .A(U1_pipe8[20]), .B(n28825), .CO(n21474), .S(n21408) );
  ADDHXL U8455 ( .A(U0_pipe5[19]), .B(U0_pipe4[19]), .CO(n24076), .S(n24018)
         );
  ADDHXL U8456 ( .A(U0_pipe8[19]), .B(n28762), .CO(n26749), .S(n26669) );
  ADDHXL U8457 ( .A(U1_pipe14[20]), .B(n28873), .CO(n18725), .S(n18662) );
  ADDHXL U8458 ( .A(U1_pipe8[19]), .B(n28826), .CO(n21409), .S(n21354) );
  ADDHXL U8459 ( .A(U0_pipe5[24]), .B(U0_pipe4[24]), .CO(n24316), .S(n24273)
         );
  ADDHXL U8460 ( .A(U1_pipe7[24]), .B(U1_pipe6[24]), .CO(n18940), .S(n18898)
         );
  ADDHXL U8461 ( .A(U1_pipe14[17]), .B(n28876), .CO(n18557), .S(n18516) );
  ADDHXL U8462 ( .A(U0_pipe5[20]), .B(U0_pipe4[20]), .CO(n24139), .S(n24075)
         );
  NOR2X1 U8463 ( .A(n8101), .B(AOPB[46]), .Y(n10370) );
  ADDHXL U8464 ( .A(U1_pipe14[19]), .B(n28874), .CO(n18663), .S(n18607) );
  ADDHXL U8465 ( .A(U0_pipe8[22]), .B(n28926), .CO(n26885), .S(n26838) );
  NOR2X1 U8466 ( .A(ram_sel_reg[9]), .B(n28759), .Y(n14996) );
  ADDHXL U8467 ( .A(U0_pipe5[22]), .B(U0_pipe4[22]), .CO(n24233), .S(n24186)
         );
  ADDHXL U8468 ( .A(U0_pipe8[24]), .B(n28924), .CO(n26983), .S(n26925) );
  NAND2X1 U8469 ( .A(AOPC[25]), .B(n8055), .Y(n11381) );
  ADDHXL U8470 ( .A(U1_pipe8[24]), .B(n28940), .CO(n21651), .S(n21591) );
  NAND2X1 U8471 ( .A(W2[11]), .B(W2[27]), .Y(n9887) );
  ADDHXL U8472 ( .A(U1_pipe2[22]), .B(n28946), .CO(n21565), .S(n21513) );
  INVX8 U8473 ( .A(n28697), .Y(n27042) );
  NOR2X1 U8474 ( .A(n8153), .B(BOPB[49]), .Y(n10542) );
  NAND2X1 U8475 ( .A(BOPC[25]), .B(n8130), .Y(n11209) );
  ADDHXL U8476 ( .A(U1_pipe1[22]), .B(U1_pipe0[22]), .CO(n21557), .S(n21505)
         );
  ADDHXL U8477 ( .A(U1_pipe2[24]), .B(n28944), .CO(n21635), .S(n21607) );
  OR2XL U8478 ( .A(U0_U0_y2[10]), .B(U0_U0_y0[10]), .Y(n14164) );
  ADDHXL U8479 ( .A(U0_pipe11[19]), .B(U0_pipe10[19]), .CO(n24087), .S(n24006)
         );
  ADDHXL U8480 ( .A(U1_pipe8[22]), .B(n28942), .CO(n21549), .S(n21497) );
  ADDHXL U8481 ( .A(U1_pipe1[20]), .B(U1_pipe0[20]), .CO(n21462), .S(n21397)
         );
  ADDHXL U8482 ( .A(U0_pipe11[20]), .B(U0_pipe10[20]), .CO(n24126), .S(n24086)
         );
  ADDHXL U8483 ( .A(U0_pipe14[19]), .B(n28810), .CO(n24054), .S(n23994) );
  ADDHXL U8484 ( .A(U0_pipe14[20]), .B(n28809), .CO(n24114), .S(n24053) );
  ADDHXL U8485 ( .A(U0_pipe11[22]), .B(U0_pipe10[22]), .CO(n24241), .S(n24194)
         );
  ADDHXL U8486 ( .A(U1_pipe8[16]), .B(n28829), .CO(n21261), .S(n21141) );
  ADDHXL U8487 ( .A(U1_pipe2[17]), .B(n28844), .CO(n21300), .S(n21232) );
  ADDHXL U8488 ( .A(U1_pipe2[19]), .B(n28842), .CO(n21387), .S(n21331) );
  ADDHXL U8489 ( .A(U1_pipe2[20]), .B(n28841), .CO(n21450), .S(n21386) );
  ADDHXL U8490 ( .A(U1_pipe1[24]), .B(U1_pipe0[24]), .CO(n21643), .S(n21599)
         );
  ADDHXL U8491 ( .A(U0_pipe14[16]), .B(n28813), .CO(n23895), .S(n23804) );
  ADDHXL U8492 ( .A(U0_pipe14[17]), .B(n28812), .CO(n23945), .S(n23894) );
  MXI2X1 U8493 ( .A(U0_pipe5[22]), .B(n22313), .S0(n22248), .Y(n4496) );
  MXI2X1 U8494 ( .A(U0_pipe5[23]), .B(n22308), .S0(n22248), .Y(n4495) );
  MXI2X1 U8495 ( .A(U0_pipe5[25]), .B(n22299), .S0(n22248), .Y(n4493) );
  MXI2X1 U8496 ( .A(U0_pipe5[24]), .B(n22302), .S0(n22248), .Y(n4494) );
  MXI2X1 U8497 ( .A(U1_pipe14[26]), .B(n9606), .S0(n17187), .Y(n4777) );
  MXI2X1 U8498 ( .A(U0_pipe5[21]), .B(n22316), .S0(n22248), .Y(n4497) );
  MXI2X1 U8499 ( .A(U0_pipe13[22]), .B(n25314), .S0(n25318), .Y(n4670) );
  MXI2X1 U8500 ( .A(U1_pipe13[21]), .B(n20054), .S0(n20025), .Y(n4744) );
  MXI2X1 U8501 ( .A(U1_pipe2[24]), .B(n19080), .S0(n24784), .Y(n5036) );
  MXI2X1 U8502 ( .A(U0_pipe7[23]), .B(n21966), .S0(n22248), .Y(n4439) );
  MXI2X1 U8503 ( .A(U1_pipe2[25]), .B(n19071), .S0(n24784), .Y(n5037) );
  MXI2X1 U8504 ( .A(U1_pipe0[22]), .B(n19402), .S0(n19405), .Y(n5125) );
  MXI2X1 U8505 ( .A(U0_pipe9[25]), .B(n12285), .S0(n6887), .Y(n4580) );
  MXI2X1 U8506 ( .A(U0_pipe13[21]), .B(n25319), .S0(n25318), .Y(n4671) );
  XOR2X1 U8507 ( .A(n19387), .B(n14899), .Y(n6191) );
  MXI2X1 U8508 ( .A(U1_pipe0[25]), .B(n13718), .S0(n6888), .Y(n5128) );
  NAND2XL U8509 ( .A(n6078), .B(n5812), .Y(n6077) );
  MXI2X1 U8510 ( .A(U0_pipe7[22]), .B(n21973), .S0(n21972), .Y(n4440) );
  MXI2X1 U8511 ( .A(U1_pipe0[23]), .B(n19397), .S0(n19405), .Y(n5126) );
  MXI2X1 U8512 ( .A(U0_pipe1[23]), .B(n24996), .S0(n25101), .Y(n4261) );
  NAND2X1 U8513 ( .A(n24989), .B(n6360), .Y(n6529) );
  XNOR2X1 U8514 ( .A(n20043), .B(n6118), .Y(n20044) );
  NAND2XL U8515 ( .A(n6681), .B(n6682), .Y(n7030) );
  XOR2X1 U8516 ( .A(n14109), .B(n7862), .Y(n14110) );
  MXI2X1 U8517 ( .A(U1_pipe12[25]), .B(n19794), .S0(n19405), .Y(n4720) );
  NOR2XL U8518 ( .A(n7484), .B(n7485), .Y(n7483) );
  MXI2X1 U8519 ( .A(U0_pipe3[24]), .B(n24709), .S0(n25273), .Y(n4351) );
  MXI2X1 U8520 ( .A(U1_pipe5[24]), .B(n17057), .S0(n5804), .Y(n4921) );
  MXI2X1 U8521 ( .A(U0_pipe7[25]), .B(n21951), .S0(n22248), .Y(n4437) );
  MXI2X1 U8522 ( .A(U0_pipe1[21]), .B(n25005), .S0(n25101), .Y(n4263) );
  MXI2XL U8523 ( .A(n5941), .B(U1_pipe7[24]), .S0(n5940), .Y(n4977) );
  XOR2X1 U8524 ( .A(n6079), .B(n16798), .Y(n6078) );
  INVX1 U8525 ( .A(n6528), .Y(n24989) );
  MXI2X1 U8526 ( .A(U1_pipe14[21]), .B(n17197), .S0(n5809), .Y(n4772) );
  MXI2XL U8527 ( .A(n5972), .B(U1_pipe7[22]), .S0(n5971), .Y(n4975) );
  MXI2X1 U8528 ( .A(U1_pipe7[21]), .B(n16807), .S0(n5812), .Y(n4974) );
  MXI2X1 U8529 ( .A(U0_pipe1[24]), .B(n24991), .S0(n25101), .Y(n4407) );
  MXI2X1 U8530 ( .A(U1_pipe4[20]), .B(n16964), .S0(n5812), .Y(n5088) );
  MXI2X1 U8531 ( .A(U1_pipe9[20]), .B(n14892), .S0(n6888), .Y(n4830) );
  MXI2X1 U8532 ( .A(U1_pipe12[22]), .B(n19817), .S0(n19405), .Y(n4717) );
  MXI2X1 U8533 ( .A(U1_pipe12[23]), .B(n19810), .S0(n19405), .Y(n4718) );
  MXI2X1 U8534 ( .A(U1_pipe14[24]), .B(n17179), .S0(n17187), .Y(n4775) );
  MXI2X1 U8535 ( .A(U0_pipe3[23]), .B(n24719), .S0(n25273), .Y(n4352) );
  MXI2X1 U8536 ( .A(U1_pipe9[21]), .B(n20351), .S0(n20240), .Y(n4831) );
  MXI2X1 U8537 ( .A(U1_pipe4[22]), .B(n16954), .S0(n5812), .Y(n5090) );
  MXI2X1 U8538 ( .A(U0_pipe1[18]), .B(n25023), .S0(n25101), .Y(n4266) );
  MXI2X1 U8539 ( .A(U1_pipe0[21]), .B(n19406), .S0(n19405), .Y(n5124) );
  MXI2X1 U8540 ( .A(U1_pipe2[21]), .B(n19101), .S0(n24784), .Y(n5033) );
  MXI2X1 U8541 ( .A(U1_pipe4[23]), .B(n16949), .S0(n5805), .Y(n5091) );
  MXI2X1 U8542 ( .A(U1_pipe0[24]), .B(n19391), .S0(n19405), .Y(n5127) );
  MXI2X1 U8543 ( .A(U1_pipe5[21]), .B(n17070), .S0(n25267), .Y(n4918) );
  MXI2X1 U8544 ( .A(U1_pipe10[24]), .B(n17460), .S0(n17641), .Y(n4862) );
  MXI2X1 U8545 ( .A(U0_pipe7[21]), .B(n21977), .S0(n21972), .Y(n4441) );
  NAND3XL U8546 ( .A(n7872), .B(n5986), .C(n5920), .Y(n6098) );
  MXI2X1 U8547 ( .A(U0_pipe13[17]), .B(n25346), .S0(n6887), .Y(n4675) );
  MXI2X1 U8548 ( .A(U1_pipe8[23]), .B(n20199), .S0(n20438), .Y(n5004) );
  MXI2X1 U8549 ( .A(U1_pipe4[24]), .B(n16943), .S0(n6888), .Y(n5092) );
  XOR2XL U8550 ( .A(n17069), .B(n17068), .Y(n17070) );
  MXI2X1 U8551 ( .A(U1_pipe9[18]), .B(n20359), .S0(n20025), .Y(n4828) );
  MXI2X1 U8552 ( .A(U1_pipe11[21]), .B(n17626), .S0(n5812), .Y(n4887) );
  NAND2XL U8553 ( .A(n19793), .B(n6625), .Y(n6624) );
  MXI2X1 U8554 ( .A(U1_pipe4[21]), .B(n16956), .S0(n5812), .Y(n5089) );
  MXI2X1 U8555 ( .A(U0_pipe1[17]), .B(n25026), .S0(n25101), .Y(n4267) );
  MXI2X1 U8556 ( .A(U0_pipe3[21]), .B(n24728), .S0(n25273), .Y(n4354) );
  NOR2XL U8557 ( .A(n7479), .B(n7480), .Y(n6682) );
  MXI2X1 U8558 ( .A(U1_pipe8[25]), .B(n20191), .S0(n20240), .Y(n5006) );
  MXI2X1 U8559 ( .A(U0_pipe13[19]), .B(n25335), .S0(n6887), .Y(n4673) );
  NAND2BXL U8560 ( .AN(n7853), .B(n6113), .Y(n6112) );
  INVX1 U8561 ( .A(n6004), .Y(n6001) );
  MXI2X1 U8562 ( .A(U1_pipe12[21]), .B(n19821), .S0(n19405), .Y(n4716) );
  XOR2X1 U8563 ( .A(n16792), .B(n5942), .Y(n5941) );
  MXI2X1 U8564 ( .A(U1_pipe9[19]), .B(n20354), .S0(n20240), .Y(n4829) );
  MXI2X1 U8565 ( .A(U1_pipe5[16]), .B(n17091), .S0(n17187), .Y(n4913) );
  MXI2X1 U8566 ( .A(U1_pipe12[20]), .B(n19832), .S0(n19405), .Y(n4715) );
  NAND2X1 U8567 ( .A(n6080), .B(n16795), .Y(n6079) );
  MXI2X1 U8568 ( .A(U1_pipe2[18]), .B(n19122), .S0(n17641), .Y(n5030) );
  MXI2X1 U8569 ( .A(U0_pipe11[23]), .B(n22988), .S0(n22853), .Y(n4526) );
  MXI2X1 U8570 ( .A(U1_pipe0[18]), .B(n19427), .S0(n19405), .Y(n5121) );
  MXI2X1 U8571 ( .A(U0_pipe11[21]), .B(n22998), .S0(n22620), .Y(n4528) );
  MXI2X1 U8572 ( .A(U1_pipe5[19]), .B(n17073), .S0(n17187), .Y(n4916) );
  MXI2X1 U8573 ( .A(U1_pipe14[18]), .B(n17206), .S0(n5809), .Y(n4769) );
  MXI2X1 U8574 ( .A(U1_pipe13[18]), .B(n20075), .S0(n20025), .Y(n4741) );
  MXI2X1 U8575 ( .A(U0_pipe15[21]), .B(n22615), .S0(n22620), .Y(n4615) );
  NAND2X1 U8576 ( .A(n6458), .B(n25657), .Y(n6456) );
  MXI2X1 U8577 ( .A(U1_pipe0[20]), .B(n19418), .S0(n19405), .Y(n5123) );
  XOR2X1 U8578 ( .A(n6059), .B(n6058), .Y(n7338) );
  MXI2X1 U8579 ( .A(U0_pipe7[18]), .B(n21995), .S0(n21972), .Y(n4444) );
  MXI2X1 U8580 ( .A(U0_pipe3[20]), .B(n24737), .S0(n25273), .Y(n4355) );
  NOR3X1 U8581 ( .A(n20335), .B(n7799), .C(n7873), .Y(n6135) );
  MXI2X1 U8582 ( .A(U1_pipe15[21]), .B(n17321), .S0(n25267), .Y(n4800) );
  INVX2 U8583 ( .A(n25289), .Y(n25317) );
  MXI2X1 U8584 ( .A(U0_pipe1[20]), .B(n25013), .S0(n25101), .Y(n4264) );
  MXI2X1 U8585 ( .A(U0_pipe7[20]), .B(n21986), .S0(n21972), .Y(n4442) );
  MXI2X1 U8586 ( .A(U0_pipe9[20]), .B(n25687), .S0(n6887), .Y(n4585) );
  MXI2X1 U8587 ( .A(U1_pipe15[19]), .B(n17337), .S0(n25267), .Y(n4798) );
  MXI2X1 U8588 ( .A(U0_pipe3[22]), .B(n24723), .S0(n25273), .Y(n4353) );
  MXI2X1 U8589 ( .A(U1_pipe8[22]), .B(n20204), .S0(n20438), .Y(n5003) );
  NAND2XL U8590 ( .A(n20336), .B(n7476), .Y(n7475) );
  MXI2X1 U8591 ( .A(U0_pipe15[24]), .B(n22598), .S0(n22620), .Y(n4612) );
  NAND2XL U8592 ( .A(n7214), .B(n13651), .Y(n7213) );
  MXI2X1 U8593 ( .A(U0_pipe6[18]), .B(n21856), .S0(n20438), .Y(n4472) );
  MXI2X1 U8594 ( .A(U1_pipe8[21]), .B(n20207), .S0(n20438), .Y(n5002) );
  NAND3X2 U8595 ( .A(n6470), .B(n6383), .C(n6379), .Y(n25289) );
  NAND2X1 U8596 ( .A(n20333), .B(n7814), .Y(n20336) );
  MXI2X1 U8597 ( .A(U0_pipe4[22]), .B(n22195), .S0(n22248), .Y(n4325) );
  AOI21X1 U8598 ( .A0(n7157), .A1(n6061), .B0(n6060), .Y(n6059) );
  MXI2X1 U8599 ( .A(U0_pipe4[23]), .B(n22190), .S0(n22248), .Y(n4324) );
  MXI2X1 U8600 ( .A(U0_pipe1[14]), .B(n25043), .S0(n25091), .Y(n4270) );
  MXI2X1 U8601 ( .A(U0_pipe7[17]), .B(n21999), .S0(n21972), .Y(n4445) );
  MXI2X1 U8602 ( .A(U0_pipe14[21]), .B(n22487), .S0(n25318), .Y(n4643) );
  MXI2X1 U8603 ( .A(U0_pipe12[18]), .B(n25177), .S0(n5810), .Y(n4702) );
  MXI2X1 U8604 ( .A(U0_pipe9[16]), .B(n25708), .S0(n6887), .Y(n4589) );
  MXI2X1 U8605 ( .A(U0_pipe1[19]), .B(n25017), .S0(n25101), .Y(n4265) );
  MXI2X1 U8606 ( .A(U1_pipe10[18]), .B(n17497), .S0(n17641), .Y(n4856) );
  MXI2X1 U8607 ( .A(U0_pipe7[19]), .B(n21989), .S0(n21972), .Y(n4443) );
  MXI2X1 U8608 ( .A(U0_pipe9[18]), .B(n25696), .S0(n6887), .Y(n4587) );
  MXI2X1 U8609 ( .A(U0_pipe13[16]), .B(n25356), .S0(n6887), .Y(n4676) );
  MXI2X1 U8610 ( .A(U0_pipe15[19]), .B(n22621), .S0(n22620), .Y(n4617) );
  MXI2X1 U8611 ( .A(U1_pipe13[19]), .B(n20068), .S0(n20025), .Y(n4742) );
  NAND2XL U8612 ( .A(n5843), .B(n7814), .Y(n6719) );
  MXI2X1 U8613 ( .A(U0_pipe10[25]), .B(n22743), .S0(n24784), .Y(n4552) );
  MXI2X1 U8614 ( .A(U1_pipe13[17]), .B(n20078), .S0(n20025), .Y(n4740) );
  MXI2X1 U8615 ( .A(U0_pipe3[17]), .B(n24751), .S0(n25273), .Y(n4358) );
  MXI2X1 U8616 ( .A(U1_pipe0[19]), .B(n19421), .S0(n19405), .Y(n5122) );
  MXI2X1 U8617 ( .A(U1_pipe10[20]), .B(n17486), .S0(n17641), .Y(n4858) );
  MXI2X1 U8618 ( .A(U0_pipe7[16]), .B(n22008), .S0(n21972), .Y(n4446) );
  MXI2X1 U8619 ( .A(U1_pipe8[24]), .B(n20193), .S0(n20438), .Y(n5005) );
  NAND2XL U8620 ( .A(n6349), .B(n25024), .Y(n25022) );
  MXI2X1 U8621 ( .A(U1_pipe14[19]), .B(n17201), .S0(n5809), .Y(n4770) );
  MXI2X1 U8622 ( .A(U0_pipe9[19]), .B(n25690), .S0(n6887), .Y(n4586) );
  NOR2X1 U8623 ( .A(n7863), .B(n7814), .Y(n17050) );
  MXI2X1 U8624 ( .A(U0_pipe14[24]), .B(n22472), .S0(n5805), .Y(n4640) );
  MXI2X1 U8625 ( .A(U0_pipe5[19]), .B(n22328), .S0(n22248), .Y(n4499) );
  MXI2X1 U8626 ( .A(U1_pipe6[18]), .B(n16673), .S0(n17187), .Y(n4943) );
  MXI2X1 U8627 ( .A(U1_pipe15[17]), .B(n17348), .S0(n25267), .Y(n4796) );
  AOI2BB1XL U8628 ( .A0N(n5842), .A1N(n24987), .B0(n6532), .Y(n6360) );
  MXI2X1 U8629 ( .A(U0_pipe11[17]), .B(n23025), .S0(n22620), .Y(n4532) );
  MXI2X1 U8630 ( .A(U1_pipe5[17]), .B(n17082), .S0(n17187), .Y(n4914) );
  MXI2X1 U8631 ( .A(U1_pipe2[19]), .B(n19115), .S0(n24784), .Y(n5031) );
  MXI2X1 U8632 ( .A(U0_pipe3[19]), .B(n24741), .S0(n25273), .Y(n4356) );
  MXI2X1 U8633 ( .A(U1_pipe8[20]), .B(n20219), .S0(n20438), .Y(n5001) );
  MXI2X1 U8634 ( .A(U0_pipe11[19]), .B(n23013), .S0(n22620), .Y(n4530) );
  MXI2X1 U8635 ( .A(U0_pipe1[15]), .B(n25037), .S0(n25091), .Y(n4269) );
  MXI2X1 U8636 ( .A(U0_pipe11[16]), .B(n23035), .S0(n22620), .Y(n4533) );
  MXI2X1 U8637 ( .A(U1_pipe5[14]), .B(n17102), .S0(n17187), .Y(n4911) );
  MXI2X1 U8638 ( .A(U1_pipe2[17]), .B(n19126), .S0(n19215), .Y(n5029) );
  MXI2X1 U8639 ( .A(U1_pipe5[15]), .B(n17096), .S0(n17187), .Y(n4912) );
  MXI2X1 U8640 ( .A(U0_pipe15[16]), .B(n22641), .S0(n22620), .Y(n4620) );
  INVX1 U8641 ( .A(n6156), .Y(n17069) );
  MXI2X1 U8642 ( .A(U0_pipe15[18]), .B(n22627), .S0(n22620), .Y(n4618) );
  MXI2X1 U8643 ( .A(U0_pipe6[20]), .B(n21847), .S0(n20438), .Y(n4470) );
  NAND2XL U8644 ( .A(n6601), .B(n16642), .Y(n6600) );
  MXI2X1 U8645 ( .A(U1_pipe4[19]), .B(n16966), .S0(n5812), .Y(n5087) );
  MXI2X1 U8646 ( .A(U0_pipe14[20]), .B(n14055), .S0(n6887), .Y(n4644) );
  MXI2X1 U8647 ( .A(U0_pipe6[24]), .B(n21821), .S0(n20438), .Y(n4466) );
  MXI2X1 U8648 ( .A(U0_pipe6[25]), .B(n21814), .S0(n20438), .Y(n4465) );
  MXI2X1 U8649 ( .A(U1_pipe9[17]), .B(n20362), .S0(n22853), .Y(n4827) );
  MXI2X1 U8650 ( .A(U1_pipe8[19]), .B(n20222), .S0(n20438), .Y(n5000) );
  MXI2X1 U8651 ( .A(U1_pipe5[13]), .B(n17106), .S0(n17187), .Y(n4910) );
  MXI2X1 U8652 ( .A(U0_pipe12[17]), .B(n25181), .S0(n5810), .Y(n4703) );
  MXI2X1 U8653 ( .A(U0_pipe6[23]), .B(n21829), .S0(n20438), .Y(n4467) );
  MXI2X1 U8654 ( .A(U1_pipe10[16]), .B(n17511), .S0(n17641), .Y(n4854) );
  MXI2X1 U8655 ( .A(U1_pipe10[19]), .B(n17490), .S0(n17641), .Y(n4857) );
  MXI2X1 U8656 ( .A(U0_pipe2[21]), .B(n24448), .S0(n6888), .Y(n4382) );
  INVX1 U8657 ( .A(n25336), .Y(n25345) );
  MXI2X1 U8658 ( .A(U0_pipe15[14]), .B(n22652), .S0(n22620), .Y(n4622) );
  NAND2XL U8659 ( .A(n6815), .B(n22884), .Y(n6813) );
  NAND2X1 U8660 ( .A(n19578), .B(n6868), .Y(n5954) );
  MXI2X1 U8661 ( .A(U0_pipe14[18]), .B(n22496), .S0(n25318), .Y(n4646) );
  MXI2X1 U8662 ( .A(U0_pipe4[24]), .B(n22184), .S0(n22248), .Y(n4323) );
  MXI2X1 U8663 ( .A(U0_pipe1[13]), .B(n25047), .S0(n25091), .Y(n4271) );
  MXI2X1 U8664 ( .A(U0_pipe6[16]), .B(n21869), .S0(n20438), .Y(n4474) );
  MXI2X1 U8665 ( .A(U1_pipe1[17]), .B(n19615), .S0(n20025), .Y(n5148) );
  MXI2X1 U8666 ( .A(U0_pipe6[17]), .B(n21859), .S0(n20438), .Y(n4473) );
  INVXL U8667 ( .A(n6350), .Y(n25019) );
  MXI2X1 U8668 ( .A(U1_pipe10[17]), .B(n17501), .S0(n17641), .Y(n4855) );
  MXI2X1 U8669 ( .A(U0_pipe11[14]), .B(n23046), .S0(n22620), .Y(n4535) );
  MXI2X1 U8670 ( .A(U0_pipe6[19]), .B(n21850), .S0(n20438), .Y(n4471) );
  NAND2BXL U8671 ( .AN(n22592), .B(n22591), .Y(n7208) );
  NAND2XL U8672 ( .A(n6586), .B(n16665), .Y(n6585) );
  MXI2X1 U8673 ( .A(U0_pipe15[15]), .B(n22646), .S0(n22620), .Y(n4621) );
  MXI2X1 U8674 ( .A(U0_pipe11[15]), .B(n23040), .S0(n22620), .Y(n4534) );
  MXI2X1 U8675 ( .A(U0_pipe13[15]), .B(n25361), .S0(n6887), .Y(n4677) );
  MXI2X1 U8676 ( .A(U1_pipe9[16]), .B(n20371), .S0(n22853), .Y(n4826) );
  MXI2X1 U8677 ( .A(U0_pipe2[20]), .B(n24459), .S0(n6888), .Y(n4383) );
  MXI2X1 U8678 ( .A(U0_pipe4[21]), .B(n22198), .S0(n22248), .Y(n4326) );
  MXI2X1 U8679 ( .A(U0_pipe2[18]), .B(n24472), .S0(n6888), .Y(n4385) );
  MXI2X1 U8680 ( .A(U0_pipe6[22]), .B(n21835), .S0(n20438), .Y(n4468) );
  MXI2X1 U8681 ( .A(U0_pipe8[23]), .B(n25541), .S0(n6888), .Y(n4411) );
  MXI2X1 U8682 ( .A(U1_pipe0[16]), .B(n19439), .S0(n19405), .Y(n5119) );
  MXI2X1 U8683 ( .A(U1_pipe3[20]), .B(n19261), .S0(n19215), .Y(n5060) );
  MXI2X1 U8684 ( .A(U0_pipe8[25]), .B(n25532), .S0(n6888), .Y(n4409) );
  MXI2X1 U8685 ( .A(U0_pipe5[16]), .B(n22345), .S0(n22248), .Y(n4502) );
  MXI2X1 U8686 ( .A(U0_pipe7[14]), .B(n22019), .S0(n21972), .Y(n4448) );
  INVX1 U8687 ( .A(n7006), .Y(n6306) );
  INVXL U8688 ( .A(n22300), .Y(n6200) );
  MXI2X1 U8689 ( .A(U1_pipe14[16]), .B(n17219), .S0(n5809), .Y(n4767) );
  MXI2X1 U8690 ( .A(U0_pipe3[15]), .B(n24765), .S0(n25273), .Y(n4360) );
  XOR2X1 U8691 ( .A(n6153), .B(n13095), .Y(n13096) );
  MXI2X1 U8692 ( .A(U1_pipe6[19]), .B(n16667), .S0(n17187), .Y(n4944) );
  MXI2X1 U8693 ( .A(U1_pipe0[17]), .B(n19430), .S0(n19405), .Y(n5120) );
  MXI2X1 U8694 ( .A(U1_pipe3[18]), .B(n19271), .S0(n20438), .Y(n5058) );
  MXI2X1 U8695 ( .A(U0_pipe9[15]), .B(n25713), .S0(n6887), .Y(n4590) );
  NAND3BX2 U8696 ( .AN(n13707), .B(n7686), .C(n7687), .Y(n19392) );
  AND2X2 U8697 ( .A(n21948), .B(n21949), .Y(n22298) );
  MXI2X1 U8698 ( .A(U0_pipe7[15]), .B(n22013), .S0(n21972), .Y(n4447) );
  MXI2X1 U8699 ( .A(U0_pipe0[24]), .B(n24872), .S0(n24784), .Y(n4288) );
  MXI2X1 U8700 ( .A(U0_pipe12[16]), .B(n25192), .S0(n5810), .Y(n4704) );
  MXI2X1 U8701 ( .A(U0_pipe9[17]), .B(n25698), .S0(n6887), .Y(n4588) );
  MXI2X1 U8702 ( .A(U1_pipe7[16]), .B(n16841), .S0(n24784), .Y(n4969) );
  MXI2X1 U8703 ( .A(U1_pipe13[16]), .B(n20088), .S0(n20025), .Y(n4739) );
  MXI2X1 U8704 ( .A(U1_pipe14[17]), .B(n17210), .S0(n5809), .Y(n4768) );
  MXI2X1 U8705 ( .A(U0_pipe3[14]), .B(n24770), .S0(n25273), .Y(n4361) );
  MXI2X1 U8706 ( .A(U0_pipe0[18]), .B(n24895), .S0(n24784), .Y(n4294) );
  MXI2X1 U8707 ( .A(U0_pipe8[19]), .B(n25564), .S0(n25611), .Y(n4415) );
  MXI2X1 U8708 ( .A(U0_pipe13[14]), .B(n25367), .S0(n6887), .Y(n4678) );
  MXI2X1 U8709 ( .A(U0_pipe5[18]), .B(n22334), .S0(n22248), .Y(n4500) );
  MXI2X1 U8710 ( .A(U1_pipe6[17]), .B(n16677), .S0(n5812), .Y(n4942) );
  MXI2X1 U8711 ( .A(U0_pipe2[25]), .B(n24420), .S0(n24784), .Y(n4378) );
  MXI2X1 U8712 ( .A(U2_pipe2[24]), .B(n21659), .S0(n21700), .Y(n4195) );
  MXI2X1 U8713 ( .A(U0_pipe3[13]), .B(n24774), .S0(n25091), .Y(n4362) );
  INVX1 U8714 ( .A(n25286), .Y(n25654) );
  INVXL U8715 ( .A(n25685), .Y(n25329) );
  MXI2X1 U8716 ( .A(U1_pipe15[15]), .B(n17361), .S0(n22853), .Y(n4794) );
  NAND2XL U8717 ( .A(n7854), .B(n7855), .Y(n6116) );
  MXI2X1 U8718 ( .A(U1_pipe9[15]), .B(n20376), .S0(n22853), .Y(n4825) );
  MXI2X1 U8719 ( .A(U1_pipe6[16]), .B(n16687), .S0(n17641), .Y(n4941) );
  MXI2X1 U8720 ( .A(U0_pipe12[15]), .B(n25196), .S0(n5810), .Y(n4705) );
  MXI2X1 U8721 ( .A(U1_pipe9[14]), .B(n20382), .S0(n22853), .Y(n4824) );
  MXI2X1 U8722 ( .A(U1_pipe15[14]), .B(n17367), .S0(n22853), .Y(n4793) );
  MXI2X1 U8723 ( .A(U0_pipe4[19]), .B(n22209), .S0(n22248), .Y(n4328) );
  MXI2X1 U8724 ( .A(U0_pipe12[14]), .B(n25202), .S0(n5810), .Y(n4706) );
  MXI2X1 U8725 ( .A(U0_pipe2[19]), .B(n24464), .S0(n6888), .Y(n4384) );
  MXI2X1 U8726 ( .A(U0_pipe9[14]), .B(n25719), .S0(n6887), .Y(n4591) );
  NAND2X1 U8727 ( .A(n7903), .B(n7254), .Y(n7857) );
  NAND2BXL U8728 ( .AN(n25293), .B(n25652), .Y(n6474) );
  MXI2X1 U8729 ( .A(U0_pipe4[18]), .B(n22215), .S0(n22248), .Y(n4329) );
  MXI2X1 U8730 ( .A(U0_pipe4[16]), .B(n22226), .S0(n22543), .Y(n4331) );
  MXI2X1 U8731 ( .A(U1_pipe11[14]), .B(n17661), .S0(n17641), .Y(n4880) );
  MXI2X1 U8732 ( .A(U0_pipe2[16]), .B(n24487), .S0(n6888), .Y(n4387) );
  OAI21X1 U8733 ( .A0(n19599), .A1(n19598), .B0(n6230), .Y(n19607) );
  MXI2X1 U8734 ( .A(U1_pipe11[15]), .B(n17656), .S0(n5812), .Y(n4881) );
  MXI2X1 U8735 ( .A(U1_pipe7[10]), .B(n16880), .S0(n5812), .Y(n4963) );
  MXI2X1 U8736 ( .A(U1_pipe10[15]), .B(n17515), .S0(n5812), .Y(n4853) );
  MXI2X1 U8737 ( .A(U0_pipe7[10]), .B(n22049), .S0(n21972), .Y(n4452) );
  MXI2X1 U8738 ( .A(U1_pipe11[17]), .B(n17642), .S0(n17641), .Y(n4883) );
  MXI2X1 U8739 ( .A(U0_pipe7[12]), .B(n22033), .S0(n21972), .Y(n4450) );
  INVXL U8740 ( .A(n6663), .Y(n6659) );
  MXI2X1 U8741 ( .A(U0_pipe7[13]), .B(n22023), .S0(n21972), .Y(n4449) );
  MXI2X1 U8742 ( .A(U1_pipe7[12]), .B(n16864), .S0(n5812), .Y(n4965) );
  MXI2X1 U8743 ( .A(U0_pipe8[21]), .B(n25549), .S0(n25611), .Y(n4413) );
  MXI2X1 U8744 ( .A(U1_pipe2[16]), .B(n19137), .S0(n19215), .Y(n5028) );
  MXI2X1 U8745 ( .A(U1_pipe14[15]), .B(n17223), .S0(n5809), .Y(n4766) );
  MXI2X1 U8746 ( .A(U0_pipe8[18]), .B(n25570), .S0(n25611), .Y(n4416) );
  MXI2X1 U8747 ( .A(U1_pipe7[14]), .B(n16852), .S0(n5812), .Y(n4967) );
  MXI2X1 U8748 ( .A(U1_pipe10[14]), .B(n17521), .S0(n5812), .Y(n4852) );
  NAND2X1 U8749 ( .A(n20042), .B(n20326), .Y(n20342) );
  NAND2X1 U8750 ( .A(n5844), .B(n16797), .Y(n17060) );
  MXI2X1 U8751 ( .A(U1_pipe7[15]), .B(n16846), .S0(n24784), .Y(n4968) );
  MXI2X1 U8752 ( .A(U1_pipe8[17]), .B(n20231), .S0(n20438), .Y(n4998) );
  MXI2X1 U8753 ( .A(U0_pipe8[17]), .B(n25573), .S0(n25611), .Y(n4417) );
  NAND2X1 U8754 ( .A(n7337), .B(n20329), .Y(n20339) );
  MXI2X1 U8755 ( .A(U0_pipe8[16]), .B(n25582), .S0(n25611), .Y(n4418) );
  NAND2X1 U8756 ( .A(n20333), .B(n19568), .Y(n19572) );
  MXI2X1 U8757 ( .A(U1_pipe8[18]), .B(n20228), .S0(n20438), .Y(n4999) );
  INVX1 U8758 ( .A(n21990), .Y(n21998) );
  MXI2X1 U8759 ( .A(U0_pipe5[17]), .B(n22336), .S0(n22248), .Y(n4501) );
  MXI2X1 U8760 ( .A(U0_pipe11[13]), .B(n23050), .S0(n22620), .Y(n4536) );
  MXI2X1 U8761 ( .A(U0_pipe15[13]), .B(n22656), .S0(n22620), .Y(n4623) );
  MXI2X1 U8762 ( .A(U0_pipe0[21]), .B(n24886), .S0(n24784), .Y(n4291) );
  NAND2X1 U8763 ( .A(n12404), .B(n22968), .Y(n14580) );
  MXI2X1 U8764 ( .A(U0_pipe0[19]), .B(n24889), .S0(n24784), .Y(n4293) );
  MXI2X1 U8765 ( .A(U1_pipe13[14]), .B(n20098), .S0(n20025), .Y(n4737) );
  NAND3X1 U8766 ( .A(n20194), .B(n19797), .C(n12331), .Y(n6630) );
  MXI2X1 U8767 ( .A(U0_pipe2[17]), .B(n24476), .S0(n6888), .Y(n4386) );
  MXI2X1 U8768 ( .A(U1_pipe13[15]), .B(n20093), .S0(n20025), .Y(n4738) );
  INVXL U8769 ( .A(n19429), .Y(n19424) );
  MXI2X1 U8770 ( .A(U1_pipe3[16]), .B(n19285), .S0(n20438), .Y(n5056) );
  MXI2X1 U8771 ( .A(U0_pipe14[19]), .B(n22491), .S0(n25318), .Y(n4645) );
  MXI2X1 U8772 ( .A(U1_pipe3[19]), .B(n19266), .S0(n20438), .Y(n5059) );
  NAND2X2 U8773 ( .A(n6676), .B(n7402), .Y(n16633) );
  INVX1 U8774 ( .A(n20316), .Y(n14888) );
  MXI2X1 U8775 ( .A(U0_pipe10[18]), .B(n22778), .S0(n22853), .Y(n4559) );
  MXI2X1 U8776 ( .A(U1_pipe3[17]), .B(n19275), .S0(n20438), .Y(n5057) );
  MXI2X1 U8777 ( .A(U0_pipe6[15]), .B(n21872), .S0(n20438), .Y(n4475) );
  MXI2X1 U8778 ( .A(U0_pipe5[14]), .B(n22356), .S0(n22248), .Y(n4504) );
  MXI2X1 U8779 ( .A(U0_pipe6[14]), .B(n21877), .S0(n20438), .Y(n4476) );
  MXI2X1 U8780 ( .A(U1_pipe1[14]), .B(n19634), .S0(n20025), .Y(n5145) );
  MXI2X1 U8781 ( .A(U0_pipe5[15]), .B(n22350), .S0(n22248), .Y(n4503) );
  MXI2X1 U8782 ( .A(U0_pipe10[20]), .B(n14106), .S0(n6888), .Y(n4557) );
  MXI2X1 U8783 ( .A(U1_pipe1[15]), .B(n19628), .S0(n20025), .Y(n5146) );
  MXI2X1 U8784 ( .A(U1_pipe0[15]), .B(n19442), .S0(n19405), .Y(n5118) );
  MXI2X1 U8785 ( .A(U1_pipe11[12]), .B(n17674), .S0(n5812), .Y(n4878) );
  MXI2X1 U8786 ( .A(U1_pipe11[10]), .B(n17689), .S0(n17641), .Y(n4876) );
  NOR2BXL U8787 ( .AN(n13624), .B(n17299), .Y(n7860) );
  MXI2X1 U8788 ( .A(U1_pipe7[13]), .B(n16856), .S0(n5812), .Y(n4966) );
  MXI2X1 U8789 ( .A(U1_pipe2[14]), .B(n19147), .S0(n19215), .Y(n5026) );
  MXI2X1 U8790 ( .A(U1_pipe2[15]), .B(n19141), .S0(n19215), .Y(n5027) );
  MXI2X1 U8791 ( .A(U0_pipe10[17]), .B(n22782), .S0(n22853), .Y(n4560) );
  MXI2X1 U8792 ( .A(U1_pipe15[12]), .B(n17380), .S0(n22853), .Y(n4791) );
  NOR2X1 U8793 ( .A(n13178), .B(n22960), .Y(n21955) );
  MXI2X1 U8794 ( .A(U0_pipe10[16]), .B(n22792), .S0(n22853), .Y(n4561) );
  NAND2X1 U8795 ( .A(n22960), .B(n13178), .Y(n21956) );
  MXI2X1 U8796 ( .A(U0_pipe2[12]), .B(n24512), .S0(n24784), .Y(n4391) );
  MXI2X1 U8797 ( .A(U1_pipe15[10]), .B(n17393), .S0(n24784), .Y(n4789) );
  NAND2X1 U8798 ( .A(n24677), .B(n13178), .Y(n25293) );
  MXI2X1 U8799 ( .A(U0_pipe12[13]), .B(n25206), .S0(n5810), .Y(n4707) );
  NAND2BX1 U8800 ( .AN(n17176), .B(n17175), .Y(n7751) );
  MXI2X1 U8801 ( .A(U1_pipe11[11]), .B(n17679), .S0(n5812), .Y(n4877) );
  MXI2X1 U8802 ( .A(U0_pipe10[19]), .B(n22772), .S0(n22853), .Y(n4558) );
  MXI2X1 U8803 ( .A(U2_pipe3[24]), .B(n18946), .S0(n18987), .Y(n4247) );
  MXI2X1 U8804 ( .A(U0_pipe6[13]), .B(n21880), .S0(n20438), .Y(n4477) );
  OR2X2 U8805 ( .A(n14972), .B(n20028), .Y(n13987) );
  MXI2X1 U8806 ( .A(U1_pipe11[13]), .B(n17665), .S0(n17187), .Y(n4879) );
  MXI2X1 U8807 ( .A(U0_pipe14[17]), .B(n22499), .S0(n25318), .Y(n4647) );
  NAND3BXL U8808 ( .AN(n7653), .B(n7647), .C(n7644), .Y(n7643) );
  MXI2X1 U8809 ( .A(U2_pipe3[23]), .B(n18910), .S0(n18987), .Y(n4245) );
  NAND3X1 U8810 ( .A(n6257), .B(n6255), .C(n6251), .Y(n6260) );
  MXI2X1 U8811 ( .A(U1_pipe11[9]), .B(n17694), .S0(n24784), .Y(n4875) );
  MXI2X1 U8812 ( .A(U1_pipe1[13]), .B(n19638), .S0(n20025), .Y(n5144) );
  MXI2X1 U8813 ( .A(U0_pipe7[9]), .B(n22053), .S0(n21972), .Y(n4453) );
  MXI2X1 U8814 ( .A(U1_pipe9[13]), .B(n20387), .S0(n22853), .Y(n4823) );
  MXI2X1 U8815 ( .A(U1_pipe7[9]), .B(n16884), .S0(n5804), .Y(n4962) );
  INVX1 U8816 ( .A(n25006), .Y(n25046) );
  INVX1 U8817 ( .A(n14579), .Y(n12404) );
  MXI2X1 U8818 ( .A(U0_pipe7[11]), .B(n22037), .S0(n21972), .Y(n4451) );
  MXI2X1 U8819 ( .A(U1_pipe5[12]), .B(n17113), .S0(n17187), .Y(n4909) );
  MXI2X1 U8820 ( .A(U1_pipe7[11]), .B(n16868), .S0(n24784), .Y(n4964) );
  MXI2X1 U8821 ( .A(U0_pipe14[16]), .B(n22508), .S0(n22248), .Y(n4648) );
  MXI2X1 U8822 ( .A(U0_pipe2[15]), .B(n24491), .S0(n6888), .Y(n4388) );
  MXI2X1 U8823 ( .A(U1_pipe3[14]), .B(n19296), .S0(n19215), .Y(n5054) );
  MXI2X1 U8824 ( .A(U0_pipe2[14]), .B(n24498), .S0(n6888), .Y(n4389) );
  MXI2X1 U8825 ( .A(U1_pipe14[14]), .B(n17227), .S0(n5809), .Y(n4765) );
  MXI2X1 U8826 ( .A(U1_pipe3[15]), .B(n19290), .S0(n19215), .Y(n5055) );
  MXI2X1 U8827 ( .A(U1_pipe5[10]), .B(n17124), .S0(n5804), .Y(n5106) );
  MXI2X1 U8828 ( .A(U0_pipe0[17]), .B(n24898), .S0(n24784), .Y(n4295) );
  MXI2X1 U8829 ( .A(U1_pipe6[15]), .B(n16691), .S0(n17187), .Y(n4940) );
  MXI2X1 U8830 ( .A(U0_pipe5[13]), .B(n22360), .S0(n6888), .Y(n4505) );
  NAND2X1 U8831 ( .A(n16802), .B(n16801), .Y(n17065) );
  MXI2X1 U8832 ( .A(U0_pipe8[14]), .B(n25590), .S0(n25611), .Y(n4420) );
  MXI2X1 U8833 ( .A(U0_pipe8[15]), .B(n25585), .S0(n25611), .Y(n4419) );
  MXI2X1 U8834 ( .A(U1_pipe13[10]), .B(n20126), .S0(n20025), .Y(n4733) );
  MXI2X1 U8835 ( .A(U0_pipe13[10]), .B(n25394), .S0(n6887), .Y(n4682) );
  MXI2X1 U8836 ( .A(U2_pipe2[23]), .B(n21621), .S0(n21700), .Y(n4193) );
  AND2X2 U8837 ( .A(n19563), .B(n7881), .Y(n7033) );
  MXI2X1 U8838 ( .A(U0_pipe0[16]), .B(n24907), .S0(n24784), .Y(n4296) );
  INVX1 U8839 ( .A(n25528), .Y(n7707) );
  MXI2X1 U8840 ( .A(U0_pipe4[15]), .B(n22229), .S0(n22543), .Y(n4332) );
  NOR2X1 U8841 ( .A(n17059), .B(n16796), .Y(n5968) );
  AOI21X1 U8842 ( .A0(n25722), .A1(n25702), .B0(n25701), .Y(n25712) );
  NAND3BX2 U8843 ( .AN(n14506), .B(n6040), .C(n14500), .Y(n6039) );
  NAND2X1 U8844 ( .A(n24706), .B(n24705), .Y(n24990) );
  MXI2X1 U8845 ( .A(U1_pipe0[14]), .B(n19447), .S0(n19405), .Y(n5117) );
  MXI2X1 U8846 ( .A(U0_pipe9[13]), .B(n25723), .S0(n6887), .Y(n4592) );
  INVXL U8847 ( .A(n20028), .Y(n20023) );
  MXI2X1 U8848 ( .A(U0_pipe4[14]), .B(n22234), .S0(n22543), .Y(n4333) );
  NAND2X1 U8849 ( .A(n25328), .B(n25327), .Y(n25685) );
  INVX1 U8850 ( .A(n19235), .Y(n5996) );
  AOI21X1 U8851 ( .A0(n24773), .A1(n24755), .B0(n24754), .Y(n24764) );
  OAI21X2 U8852 ( .A0(n21693), .A1(n21692), .B0(n7417), .Y(n6427) );
  MXI2X1 U8853 ( .A(U0_pipe13[12]), .B(n25380), .S0(n6887), .Y(n4680) );
  MXI2X1 U8854 ( .A(U1_pipe13[12]), .B(n20111), .S0(n20025), .Y(n4735) );
  NAND2BXL U8855 ( .AN(n19076), .B(n14895), .Y(n7746) );
  NAND2X1 U8856 ( .A(n25304), .B(n25303), .Y(n25666) );
  NAND2X1 U8857 ( .A(n20029), .B(n20028), .Y(n20331) );
  AOI21X1 U8858 ( .A0(n25370), .A1(n25350), .B0(n25349), .Y(n25360) );
  INVX1 U8859 ( .A(n16799), .Y(n7471) );
  MXI2X1 U8860 ( .A(U2_pipe0[24]), .B(n26996), .S0(n27040), .Y(n4091) );
  MXI2X1 U8861 ( .A(U0_pipe0[14]), .B(n24915), .S0(n5920), .Y(n4298) );
  MXI2X1 U8862 ( .A(U0_pipe10[15]), .B(n22796), .S0(n22853), .Y(n4562) );
  MXI2X1 U8863 ( .A(U0_pipe14[14]), .B(n22517), .S0(n22543), .Y(n4650) );
  AOI21XL U8864 ( .A0(n6954), .A1(n13704), .B0(n13703), .Y(n13705) );
  MXI2X1 U8865 ( .A(U0_pipe10[14]), .B(n22802), .S0(n22853), .Y(n4563) );
  NOR2X1 U8866 ( .A(n14968), .B(n20032), .Y(n16789) );
  NAND2X1 U8867 ( .A(n20041), .B(n5845), .Y(n20326) );
  NOR2X1 U8868 ( .A(n20046), .B(n20018), .Y(n20037) );
  MXI2X1 U8869 ( .A(U0_pipe0[15]), .B(n24910), .S0(n24784), .Y(n4297) );
  NAND2X1 U8870 ( .A(n14966), .B(n5845), .Y(n16797) );
  AOI21X1 U8871 ( .A0(n20386), .A1(n20366), .B0(n20365), .Y(n20375) );
  INVX1 U8872 ( .A(n19267), .Y(n19274) );
  MXI2X1 U8873 ( .A(U0_pipe8[13]), .B(n25593), .S0(n25611), .Y(n4421) );
  CLKINVX3 U8874 ( .A(n19567), .Y(n20333) );
  MXI2X1 U8875 ( .A(U0_pipe11[12]), .B(n23059), .S0(n22620), .Y(n4537) );
  MXI2X1 U8876 ( .A(U0_pipe15[12]), .B(n22664), .S0(n22620), .Y(n4624) );
  NOR2X1 U8877 ( .A(n5958), .B(n20355), .Y(n5957) );
  MXI2X1 U8878 ( .A(U1_pipe5[9]), .B(n17127), .S0(n5804), .Y(n5105) );
  NAND2X1 U8879 ( .A(n5847), .B(n24693), .Y(n22969) );
  MXI2X1 U8880 ( .A(U0_pipe5[10]), .B(n22379), .S0(n19405), .Y(n4309) );
  MXI2X1 U8881 ( .A(U1_pipe0[12]), .B(n19456), .S0(n19405), .Y(n5115) );
  MXI2X1 U8882 ( .A(U1_pipe0[13]), .B(n19449), .S0(n19405), .Y(n5116) );
  NAND2BX1 U8883 ( .AN(n24693), .B(n5846), .Y(n12342) );
  MXI2X1 U8884 ( .A(U1_pipe13[9]), .B(n20131), .S0(n20025), .Y(n4732) );
  AOI21X1 U8885 ( .A0(n13947), .A1(n6936), .B0(n13946), .Y(n6032) );
  MXI2X1 U8886 ( .A(U1_pipe13[11]), .B(n20116), .S0(n20025), .Y(n4734) );
  AOI21X1 U8887 ( .A0(n20101), .A1(n20082), .B0(n20081), .Y(n20092) );
  MXI2X1 U8888 ( .A(U0_pipe3[12]), .B(n24785), .S0(n24784), .Y(n4363) );
  OAI2BB2XL U8889 ( .B0(n5851), .B1(U1_A_r_d0[25]), .A0N(n7526), .A1N(n7525), 
        .Y(n6566) );
  NAND2X1 U8890 ( .A(n6954), .B(n19108), .Y(n19416) );
  MXI2X1 U8891 ( .A(U0_pipe13[11]), .B(n25384), .S0(n5920), .Y(n4681) );
  MXI2X1 U8892 ( .A(U1_pipe5[11]), .B(n17116), .S0(n5804), .Y(n4908) );
  MXI2X1 U8893 ( .A(U0_pipe5[12]), .B(n22368), .S0(n19215), .Y(n4506) );
  MXI2X1 U8894 ( .A(U0_pipe2[11]), .B(n24516), .S0(n24784), .Y(n4392) );
  MXI2X1 U8895 ( .A(U1_pipe9[10]), .B(n20410), .S0(n21972), .Y(n4820) );
  INVX1 U8896 ( .A(n19564), .Y(n7881) );
  AOI21X1 U8897 ( .A0(n16855), .A1(n16835), .B0(n7035), .Y(n16845) );
  MXI2X1 U8898 ( .A(U1_pipe15[11]), .B(n17384), .S0(n5812), .Y(n4790) );
  MXI2X1 U8899 ( .A(U1_pipe3[12]), .B(n19309), .S0(n19215), .Y(n5052) );
  MXI2X1 U8900 ( .A(U0_pipe1[12]), .B(n25054), .S0(n25091), .Y(n4272) );
  AOI21X1 U8901 ( .A0(n21879), .A1(n21863), .B0(n21862), .Y(n21871) );
  AOI21X1 U8902 ( .A0(n12270), .A1(n25311), .B0(n12269), .Y(n25664) );
  MXI2X1 U8903 ( .A(U1_pipe9[12]), .B(n20396), .S0(n21972), .Y(n4822) );
  NAND2X1 U8904 ( .A(n5846), .B(n24693), .Y(n24694) );
  CLKINVX2 U8905 ( .A(n14838), .Y(n7895) );
  INVXL U8906 ( .A(n20046), .Y(n6022) );
  MXI2X1 U8907 ( .A(U2_pipe2[18]), .B(n21368), .S0(n21700), .Y(n4183) );
  INVXL U8908 ( .A(n20045), .Y(n6021) );
  AOI21X1 U8909 ( .A0(n17664), .A1(n17646), .B0(n17645), .Y(n17655) );
  INVXL U8910 ( .A(n20346), .Y(n20049) );
  INVX1 U8911 ( .A(n19594), .Y(n6231) );
  MXI2X1 U8912 ( .A(U2_pipe2[20]), .B(n21485), .S0(n21700), .Y(n4187) );
  AOI21X1 U8913 ( .A0(n19637), .A1(n19619), .B0(n19618), .Y(n19627) );
  INVX1 U8914 ( .A(n19597), .Y(n19598) );
  AOI21X1 U8915 ( .A0(n17370), .A1(n17352), .B0(n17351), .Y(n17360) );
  MXI2X1 U8916 ( .A(U0_pipe7[8]), .B(n22057), .S0(n21972), .Y(n4454) );
  MXI2X1 U8917 ( .A(U1_pipe3[10]), .B(n19325), .S0(n19215), .Y(n5050) );
  NAND2X1 U8918 ( .A(n17309), .B(n17308), .Y(n17613) );
  MXI2X1 U8919 ( .A(U1_pipe2[12]), .B(n19161), .S0(n19215), .Y(n5024) );
  MXI2X1 U8920 ( .A(U0_pipe9[10]), .B(n25746), .S0(n6887), .Y(n4595) );
  NAND2X1 U8921 ( .A(n6936), .B(n14012), .Y(n16814) );
  NOR2BX1 U8922 ( .AN(n14575), .B(n5858), .Y(n6448) );
  NAND2BX1 U8923 ( .AN(n13966), .B(n16804), .Y(n17059) );
  MXI2X1 U8924 ( .A(U0_pipe14[15]), .B(n22512), .S0(n22543), .Y(n4649) );
  INVX1 U8925 ( .A(n21815), .Y(n21837) );
  AOI21X1 U8926 ( .A0(n22498), .A1(n14052), .B0(n14051), .Y(n22490) );
  MXI2X1 U8927 ( .A(U0_pipe9[12]), .B(n25731), .S0(n6887), .Y(n4593) );
  NAND2X1 U8928 ( .A(n5797), .B(n5845), .Y(n14967) );
  MXI2X1 U8929 ( .A(U2_pipe2[22]), .B(n21579), .S0(n21700), .Y(n4191) );
  MXI2X1 U8930 ( .A(U1_pipe10[12]), .B(n17534), .S0(n5809), .Y(n4850) );
  MXI2X1 U8931 ( .A(U1_pipe3[13]), .B(n19300), .S0(n19215), .Y(n5053) );
  MXI2X1 U8932 ( .A(U1_pipe15[9]), .B(n17398), .S0(n5812), .Y(n4788) );
  MXI2X1 U8933 ( .A(U0_pipe9[9]), .B(n25751), .S0(n6887), .Y(n4596) );
  AOI21X1 U8934 ( .A0(n19150), .A1(n19130), .B0(n19129), .Y(n19140) );
  MXI2X1 U8935 ( .A(U0_pipe3[10]), .B(n24801), .S0(n24784), .Y(n4365) );
  MXI2X1 U8936 ( .A(U0_pipe11[10]), .B(n23073), .S0(n24784), .Y(n4539) );
  MXI2X1 U8937 ( .A(U0_pipe2[10]), .B(n24528), .S0(n22853), .Y(n4393) );
  MXI2X1 U8938 ( .A(U2_pipe0[20]), .B(n26826), .S0(n27040), .Y(n4083) );
  MXI2X1 U8939 ( .A(U0_pipe0[12]), .B(n24925), .S0(n5920), .Y(n4300) );
  MXI2X1 U8940 ( .A(U1_pipe3[11]), .B(n19314), .S0(n19215), .Y(n5051) );
  MXI2X1 U8941 ( .A(U1_pipe2[10]), .B(n19177), .S0(n19215), .Y(n5022) );
  MXI2X1 U8942 ( .A(U2_pipe0[17]), .B(n26652), .S0(n27040), .Y(n4077) );
  MXI2X1 U8943 ( .A(U0_pipe11[11]), .B(n23063), .S0(n22620), .Y(n4538) );
  INVX1 U8944 ( .A(n7685), .Y(n19407) );
  MXI2X1 U8945 ( .A(U0_pipe10[13]), .B(n22806), .S0(n22853), .Y(n4564) );
  MXI2X1 U8946 ( .A(U0_pipe5[11]), .B(n22371), .S0(n22853), .Y(n4507) );
  MXI2X1 U8947 ( .A(U0_pipe10[12]), .B(n22815), .S0(n22853), .Y(n4565) );
  NAND2X1 U8948 ( .A(n14895), .B(n14893), .Y(n19069) );
  MXI2X1 U8949 ( .A(U2_pipe3[22]), .B(n18869), .S0(n18987), .Y(n4243) );
  MXI2X1 U8950 ( .A(U0_pipe10[10]), .B(n22829), .S0(n22853), .Y(n4567) );
  MXI2X1 U8951 ( .A(U0_pipe0[10]), .B(n24936), .S0(n5920), .Y(n4302) );
  NAND2X1 U8952 ( .A(n22456), .B(n29009), .Y(n22460) );
  NAND3X2 U8953 ( .A(n6030), .B(n12972), .C(n6029), .Y(n17664) );
  NAND2XL U8954 ( .A(n16958), .B(n8616), .Y(n8618) );
  MXI2X1 U8955 ( .A(U2_pipe0[18]), .B(n26708), .S0(n27040), .Y(n4079) );
  MXI2X1 U8956 ( .A(U1_pipe10[11]), .B(n17538), .S0(n5809), .Y(n4849) );
  MXI2X1 U8957 ( .A(U1_pipe2[11]), .B(n19165), .S0(n19215), .Y(n5023) );
  AOI21XL U8958 ( .A0(n8612), .A1(n6906), .B0(n7532), .Y(n8613) );
  XNOR2X1 U8959 ( .A(n25398), .B(n25397), .Y(n25399) );
  MXI2X1 U8960 ( .A(U1_pipe10[10]), .B(n17548), .S0(n5809), .Y(n4848) );
  NAND2X1 U8961 ( .A(n16826), .B(n16825), .Y(n17077) );
  AOI21X1 U8962 ( .A0(n25592), .A1(n25577), .B0(n25576), .Y(n25584) );
  MXI2X1 U8963 ( .A(U2_pipe0[23]), .B(n26953), .S0(n27040), .Y(n4089) );
  NAND2X1 U8964 ( .A(n17314), .B(n17313), .Y(n17617) );
  AND2X2 U8965 ( .A(n17174), .B(n17175), .Y(n7012) );
  MXI2X1 U8966 ( .A(U0_pipe14[10]), .B(n22539), .S0(n22543), .Y(n4654) );
  NOR2X1 U8967 ( .A(n22959), .B(n14570), .Y(n21961) );
  NOR2XL U8968 ( .A(n5851), .B(n29007), .Y(n6587) );
  NOR2X1 U8969 ( .A(n20010), .B(n20079), .Y(n20056) );
  MXI2X1 U8970 ( .A(U2_pipe0[19]), .B(n26766), .S0(n27040), .Y(n4081) );
  MXI2X1 U8971 ( .A(U0_pipe3[11]), .B(n24789), .S0(n24784), .Y(n4364) );
  AOI21X1 U8972 ( .A0(n19299), .A1(n19279), .B0(n19278), .Y(n19289) );
  MXI2X1 U8973 ( .A(U1_pipe3[9]), .B(n19329), .S0(n19215), .Y(n5049) );
  INVXL U8974 ( .A(n20308), .Y(n20065) );
  MXI2X1 U8975 ( .A(U0_pipe15[10]), .B(n22677), .S0(n22620), .Y(n4626) );
  INVX1 U8976 ( .A(n25125), .Y(n21805) );
  MXI2X1 U8977 ( .A(U0_pipe1[10]), .B(n25065), .S0(n25091), .Y(n4274) );
  MXI2X1 U8978 ( .A(U0_pipe12[12]), .B(n25215), .S0(n5810), .Y(n4509) );
  AOI21X1 U8979 ( .A0(n16993), .A1(n16978), .B0(n16977), .Y(n16985) );
  MXI2X1 U8980 ( .A(U0_pipe1[11]), .B(n25057), .S0(n25091), .Y(n4273) );
  MXI2X1 U8981 ( .A(U1_pipe9[11]), .B(n20400), .S0(n21972), .Y(n4821) );
  MXI2X1 U8982 ( .A(U0_pipe14[12]), .B(n22528), .S0(n22543), .Y(n4652) );
  MXI2X1 U8983 ( .A(U2_pipe2[21]), .B(n21535), .S0(n21700), .Y(n4189) );
  MXI2X1 U8984 ( .A(U2_pipe0[15]), .B(n26522), .S0(n27040), .Y(n4073) );
  MXI2X1 U8985 ( .A(U0_pipe15[11]), .B(n22668), .S0(n22620), .Y(n4625) );
  NAND2X1 U8986 ( .A(n12333), .B(n19791), .Y(n20189) );
  MXI2X1 U8987 ( .A(U1_pipe1[12]), .B(n19646), .S0(n20025), .Y(n5143) );
  MXI2X1 U8988 ( .A(U2_pipe2[16]), .B(n21272), .S0(n21700), .Y(n4179) );
  MXI2X1 U8989 ( .A(U1_pipe0[11]), .B(n19459), .S0(n19405), .Y(n5114) );
  NOR2XL U8990 ( .A(n5851), .B(U1_A_i_d0[25]), .Y(n7164) );
  NAND2X1 U8991 ( .A(n25311), .B(n25310), .Y(n25671) );
  INVX1 U8992 ( .A(n20072), .Y(n5958) );
  MXI2X1 U8993 ( .A(U2_pipe1[24]), .B(n24337), .S0(n27040), .Y(n4143) );
  INVX1 U8994 ( .A(n24687), .Y(n6239) );
  MXI2X1 U8995 ( .A(U1_pipe6[14]), .B(n16697), .S0(n5812), .Y(n4939) );
  MXI2X1 U8996 ( .A(U2_pipe2[17]), .B(n21314), .S0(n21700), .Y(n4181) );
  MXI2X1 U8997 ( .A(U2_pipe2[19]), .B(n21428), .S0(n21700), .Y(n4185) );
  MXI2X1 U8998 ( .A(U2_pipe2[14]), .B(n21128), .S0(n21700), .Y(n4175) );
  MXI2X1 U8999 ( .A(U0_pipe9[11]), .B(n25736), .S0(n6887), .Y(n4594) );
  AOI21X1 U9000 ( .A0(n22236), .A1(n22221), .B0(n22220), .Y(n22228) );
  MXI2X1 U9001 ( .A(U0_pipe6[12]), .B(n21889), .S0(n20438), .Y(n4478) );
  INVXL U9002 ( .A(n16819), .Y(n14011) );
  MXI2X1 U9003 ( .A(U0_pipe5[9]), .B(n22382), .S0(n22620), .Y(n4310) );
  MXI2X1 U9004 ( .A(U2_pipe0[22]), .B(n26913), .S0(n27040), .Y(n4087) );
  MXI2X1 U9005 ( .A(U1_pipe9[9]), .B(n20415), .S0(n21972), .Y(n4819) );
  MXI2X1 U9006 ( .A(U1_pipe14[12]), .B(n17238), .S0(n5809), .Y(n4763) );
  NAND2X1 U9007 ( .A(n17314), .B(n17318), .Y(n17306) );
  MXI2X1 U9008 ( .A(U2_pipe3[19]), .B(n18715), .S0(n18987), .Y(n4237) );
  INVX1 U9009 ( .A(n19595), .Y(n7804) );
  MXI2X1 U9010 ( .A(U1_pipe10[9]), .B(n17552), .S0(n5809), .Y(n4847) );
  AOI21X1 U9011 ( .A0(n5854), .A1(n22503), .B0(n22502), .Y(n22511) );
  NOR2X1 U9012 ( .A(n14963), .B(n20047), .Y(n13966) );
  OR2XL U9013 ( .A(n19790), .B(n29008), .Y(n7000) );
  MXI2X1 U9014 ( .A(U2_pipe3[21]), .B(n18823), .S0(n18987), .Y(n4241) );
  MXI2X1 U9015 ( .A(U2_pipe1[23]), .B(n24294), .S0(n21700), .Y(n4141) );
  MXI2X1 U9016 ( .A(U1_pipe2[9]), .B(n19181), .S0(n19215), .Y(n5021) );
  MXI2X1 U9017 ( .A(U0_pipe0[11]), .B(n24928), .S0(n5920), .Y(n4301) );
  MXI2X1 U9018 ( .A(U0_pipe4[12]), .B(n22245), .S0(n22543), .Y(n4335) );
  NAND2X1 U9019 ( .A(n7171), .B(n5861), .Y(n17314) );
  NAND2X1 U9020 ( .A(n24758), .B(n24757), .Y(n25032) );
  MXI2X1 U9021 ( .A(U2_pipe3[13]), .B(n18365), .S0(n18987), .Y(n4225) );
  NAND3BX1 U9022 ( .AN(n14944), .B(n7465), .C(n6160), .Y(n7454) );
  NAND2BX2 U9023 ( .AN(n9685), .B(n6507), .Y(n19150) );
  MXI2X1 U9024 ( .A(U1_pipe0[10]), .B(n19467), .S0(n19405), .Y(n5113) );
  MXI2X1 U9025 ( .A(U2_pipe0[21]), .B(n26871), .S0(n27040), .Y(n4085) );
  MXI2X1 U9026 ( .A(U2_pipe3[16]), .B(n18553), .S0(n18987), .Y(n4231) );
  MXI2X1 U9027 ( .A(U1_pipe14[10]), .B(n17250), .S0(n5809), .Y(n4761) );
  MXI2X1 U9028 ( .A(U0_pipe8[12]), .B(n25600), .S0(n25611), .Y(n4422) );
  MXI2X1 U9029 ( .A(U2_pipe3[17]), .B(n18601), .S0(n18987), .Y(n4233) );
  INVXL U9030 ( .A(n5975), .Y(n16858) );
  MXI2X1 U9031 ( .A(U2_pipe1[18]), .B(n24046), .S0(n27040), .Y(n4131) );
  NAND2X1 U9032 ( .A(n19560), .B(n19558), .Y(n19585) );
  MXI2X1 U9033 ( .A(U0_pipe1[9]), .B(n25068), .S0(n25091), .Y(n4275) );
  MXI2X1 U9034 ( .A(U1_pipe6[12]), .B(n16711), .S0(n5812), .Y(n4937) );
  NAND2X1 U9035 ( .A(n5855), .B(n7913), .Y(n20072) );
  MXI2X1 U9036 ( .A(U2_pipe1[17]), .B(n23988), .S0(n21700), .Y(n4129) );
  MXI2X1 U9037 ( .A(U1_pipe14[11]), .B(n17241), .S0(n5809), .Y(n4762) );
  MXI2X1 U9038 ( .A(U0_pipe6[11]), .B(n21893), .S0(n20438), .Y(n4479) );
  INVX1 U9039 ( .A(n17666), .Y(n17697) );
  MXI2X1 U9040 ( .A(U1_pipe4[10]), .B(n17011), .S0(n17187), .Y(n5078) );
  MXI2X1 U9041 ( .A(U1_pipe6[10]), .B(n16727), .S0(n5812), .Y(n4935) );
  XNOR2XL U9042 ( .A(n24917), .B(n24916), .Y(n24918) );
  NAND2X1 U9043 ( .A(n17191), .B(n17190), .Y(n17471) );
  INVXL U9044 ( .A(n19601), .Y(n19260) );
  MXI2X1 U9045 ( .A(U2_pipe1[22]), .B(n24253), .S0(n27040), .Y(n4139) );
  MXI2X1 U9046 ( .A(U0_pipe12[10]), .B(n25230), .S0(n5810), .Y(n4511) );
  MXI2X1 U9047 ( .A(U1_pipe11[6]), .B(n17713), .S0(n17187), .Y(n4872) );
  INVXL U9048 ( .A(n17627), .Y(n14502) );
  MXI2X1 U9049 ( .A(U2_pipe1[20]), .B(n24166), .S0(n27040), .Y(n4135) );
  MXI2X1 U9050 ( .A(U0_pipe12[11]), .B(n25219), .S0(n5810), .Y(n4510) );
  NAND2X1 U9051 ( .A(n17355), .B(n17354), .Y(n17649) );
  INVX1 U9052 ( .A(n22463), .Y(n22455) );
  MXI2X1 U9053 ( .A(U1_pipe3[8]), .B(n19333), .S0(n19215), .Y(n5048) );
  MXI2X1 U9054 ( .A(U2_pipe1[19]), .B(n24104), .S0(n21700), .Y(n4133) );
  MXI2X1 U9055 ( .A(U0_pipe0[9]), .B(n24939), .S0(n5920), .Y(n4303) );
  MXI2X1 U9056 ( .A(U0_pipe6[10]), .B(n21903), .S0(n20438), .Y(n4480) );
  NOR2X1 U9057 ( .A(n22959), .B(n24684), .Y(n22602) );
  MXI2X1 U9058 ( .A(U0_pipe3[9]), .B(n24805), .S0(n24784), .Y(n4366) );
  MXI2X1 U9059 ( .A(U2_pipe2[13]), .B(n21075), .S0(n21700), .Y(n4173) );
  INVXL U9060 ( .A(n20071), .Y(n7437) );
  MXI2X1 U9061 ( .A(U2_pipe0[14]), .B(n26465), .S0(n27040), .Y(n4071) );
  MXI2X1 U9062 ( .A(U2_pipe2[15]), .B(n21195), .S0(n21700), .Y(n4177) );
  MXI2X1 U9063 ( .A(U2_pipe0[16]), .B(n26611), .S0(n27040), .Y(n4075) );
  MXI2X1 U9064 ( .A(U0_pipe14[11]), .B(n22531), .S0(n22543), .Y(n4653) );
  AND2XL U9065 ( .A(n5797), .B(n19243), .Y(n7968) );
  INVX1 U9066 ( .A(n5851), .Y(n5816) );
  MXI2X1 U9067 ( .A(U0_pipe11[9]), .B(n23078), .S0(n24784), .Y(n4540) );
  AOI21X1 U9068 ( .A0(n25353), .A1(n12391), .B0(n12390), .Y(n12392) );
  NAND2X1 U9069 ( .A(n14124), .B(n22609), .Y(n22991) );
  MXI2X1 U9070 ( .A(U0_pipe14[9]), .B(n22544), .S0(n22543), .Y(n4655) );
  MXI2X1 U9071 ( .A(U1_pipe12[12]), .B(n19881), .S0(n20025), .Y(n4906) );
  MXI2X1 U9072 ( .A(U1_pipe12[10]), .B(n19897), .S0(n20025), .Y(n4904) );
  MXI2X1 U9073 ( .A(U0_pipe15[9]), .B(n22682), .S0(n22620), .Y(n4627) );
  NOR2XL U9074 ( .A(n13713), .B(n7074), .Y(n9715) );
  NAND2X1 U9075 ( .A(n5860), .B(n24435), .Y(n24876) );
  NAND2XL U9076 ( .A(n23006), .B(n23005), .Y(n23007) );
  MXI2X1 U9077 ( .A(U2_pipe1[21]), .B(n24211), .S0(n21700), .Y(n4137) );
  INVX1 U9078 ( .A(n24748), .Y(n24743) );
  INVX1 U9079 ( .A(n19998), .Y(n5855) );
  XNOR2X1 U9080 ( .A(n21120), .B(n21074), .Y(n21075) );
  INVX1 U9081 ( .A(n19262), .Y(n19258) );
  MXI2X1 U9082 ( .A(U0_pipe12[9]), .B(n25234), .S0(n5810), .Y(n4512) );
  MXI2X1 U9083 ( .A(U2_pipe1[16]), .B(n23941), .S0(n27040), .Y(n4127) );
  INVXL U9084 ( .A(n22617), .Y(n14111) );
  MXI2X1 U9085 ( .A(U0_pipe11[8]), .B(n23082), .S0(n24784), .Y(n4541) );
  NAND2X1 U9086 ( .A(n6580), .B(n8561), .Y(n7199) );
  MXI2X1 U9087 ( .A(U0_pipe6[9]), .B(n21906), .S0(n20438), .Y(n4481) );
  NAND2X1 U9088 ( .A(n7916), .B(n14960), .Y(n14503) );
  NAND2X1 U9089 ( .A(n19992), .B(n20103), .Y(n5944) );
  NAND2X1 U9090 ( .A(n6947), .B(n19554), .Y(n19601) );
  NAND2X1 U9091 ( .A(n17359), .B(n17358), .Y(n17653) );
  MXI2X1 U9092 ( .A(U2_pipe2[12]), .B(n21024), .S0(n21023), .Y(n4171) );
  OAI21XL U9093 ( .A0(n18986), .A1(n6254), .B0(n6252), .Y(n6251) );
  MXI2X1 U9094 ( .A(U2_pipe0[11]), .B(n26297), .S0(n8054), .Y(n4065) );
  NOR2X1 U9095 ( .A(n22933), .B(n13128), .Y(n22330) );
  MXI2X1 U9096 ( .A(U1_pipe0[9]), .B(n19470), .S0(n19405), .Y(n5112) );
  NAND2X1 U9097 ( .A(n22933), .B(n13128), .Y(n22329) );
  MXI2X1 U9098 ( .A(U2_pipe0[13]), .B(n26410), .S0(n27040), .Y(n4069) );
  NAND2X1 U9099 ( .A(n19553), .B(n5856), .Y(n17627) );
  NAND3X1 U9100 ( .A(n7467), .B(n16848), .C(n16842), .Y(n6160) );
  MXI2X1 U9101 ( .A(U2_pipe0[12]), .B(n26361), .S0(n8054), .Y(n4067) );
  XNOR2X1 U9102 ( .A(n26514), .B(n26464), .Y(n26465) );
  MXI2X1 U9103 ( .A(U0_pipe15[6]), .B(n22701), .S0(n22620), .Y(n4630) );
  AOI2BB2X1 U9104 ( .B0(n8003), .B1(n14834), .A0N(n20011), .A1N(n7914), .Y(
        n19256) );
  OR2X2 U9105 ( .A(n19999), .B(n7843), .Y(n20356) );
  NAND2X1 U9106 ( .A(n7612), .B(n22477), .Y(n22755) );
  MXI2X1 U9107 ( .A(U0_pipe15[7]), .B(n22693), .S0(n22620), .Y(n4629) );
  NOR2X1 U9108 ( .A(n25374), .B(n12382), .Y(n12384) );
  NAND3X1 U9109 ( .A(n5976), .B(n5978), .C(n14936), .Y(n5975) );
  MXI2X1 U9110 ( .A(U0_pipe15[8]), .B(n22686), .S0(n22620), .Y(n4628) );
  NOR2X1 U9111 ( .A(n19248), .B(n5861), .Y(n14509) );
  MXI2X1 U9112 ( .A(U2_pipe3[10]), .B(n18195), .S0(n8054), .Y(n4219) );
  INVX1 U9113 ( .A(n16836), .Y(n16843) );
  MXI2X1 U9114 ( .A(U2_pipe3[11]), .B(n18258), .S0(n8054), .Y(n4221) );
  MXI2X1 U9115 ( .A(U2_pipe3[12]), .B(n18309), .S0(n27040), .Y(n4223) );
  MXI2X1 U9116 ( .A(U0_pipe8[11]), .B(n25603), .S0(n25611), .Y(n4423) );
  NAND2X1 U9117 ( .A(n14955), .B(n19999), .Y(n17074) );
  NOR2X1 U9118 ( .A(n17109), .B(n13887), .Y(n13889) );
  NAND2BX1 U9119 ( .AN(n19999), .B(n5868), .Y(n16830) );
  OR2X2 U9120 ( .A(n12334), .B(U1_A_r_d0[25]), .Y(n12333) );
  MXI2X1 U9121 ( .A(U0_pipe8[10]), .B(n25612), .S0(n25611), .Y(n4424) );
  NAND2X1 U9122 ( .A(n19829), .B(n19828), .Y(n20217) );
  MXI2X1 U9123 ( .A(U2_pipe1[14]), .B(n23800), .S0(n27040), .Y(n4123) );
  MXI2X1 U9124 ( .A(U2_pipe2[11]), .B(n20964), .S0(n21023), .Y(n4169) );
  AOI21X1 U9125 ( .A0(n19870), .A1(n19850), .B0(n19849), .Y(n19860) );
  MXI2X1 U9126 ( .A(U2_pipe2[10]), .B(n20909), .S0(n21023), .Y(n4167) );
  NAND2X1 U9127 ( .A(n24641), .B(n14550), .Y(n25683) );
  INVXL U9128 ( .A(n17093), .Y(n17087) );
  MXI2X1 U9129 ( .A(U2_pipe1[11]), .B(n23640), .S0(n23695), .Y(n4117) );
  MXI2X1 U9130 ( .A(U0_pipe8[9]), .B(n25615), .S0(n6888), .Y(n4425) );
  MXI2X1 U9131 ( .A(U2_pipe1[13]), .B(n23749), .S0(n21700), .Y(n4121) );
  NAND2XL U9132 ( .A(n6253), .B(n18986), .Y(n6252) );
  INVXL U9133 ( .A(n24641), .Y(n6344) );
  MXI2X1 U9134 ( .A(U2_pipe1[12]), .B(n23696), .S0(n23695), .Y(n4119) );
  NAND2BX1 U9135 ( .AN(n16853), .B(n16849), .Y(n7467) );
  INVX1 U9136 ( .A(n24642), .Y(n6314) );
  NAND2X1 U9137 ( .A(n8675), .B(n7082), .Y(n19829) );
  INVXL U9138 ( .A(n25720), .Y(n25714) );
  INVX1 U9139 ( .A(n6762), .Y(n25753) );
  MXI2X1 U9140 ( .A(U2_pipe0[10]), .B(n26246), .S0(n8054), .Y(n4063) );
  OR2X2 U9141 ( .A(n24650), .B(n24649), .Y(n24648) );
  MXI2X1 U9142 ( .A(U2_pipe0[9]), .B(n26195), .S0(n8054), .Y(n4061) );
  INVX1 U9143 ( .A(n20388), .Y(n20417) );
  NAND2BX1 U9144 ( .AN(n14945), .B(n5862), .Y(n17093) );
  NAND2X1 U9145 ( .A(n6995), .B(n14003), .Y(n24456) );
  NAND2XL U9146 ( .A(n6441), .B(n6439), .Y(n6438) );
  NAND2X1 U9147 ( .A(n14957), .B(n7914), .Y(n13070) );
  NOR2X1 U9148 ( .A(n25140), .B(U2_A_r_d[23]), .Y(n25519) );
  NAND2X1 U9149 ( .A(n20379), .B(n20384), .Y(n20363) );
  MXI2X1 U9150 ( .A(U2_pipe2[9]), .B(n20859), .S0(n21023), .Y(n4165) );
  MXI2X1 U9151 ( .A(U2_pipe2[8]), .B(n20819), .S0(n21023), .Y(n4163) );
  NAND2X1 U9152 ( .A(n7543), .B(n7071), .Y(n19839) );
  AOI21X1 U9153 ( .A0(n14542), .A1(n22027), .B0(n7965), .Y(n14543) );
  MXI2X1 U9154 ( .A(U2_pipe3[9]), .B(n18147), .S0(n8054), .Y(n4217) );
  INVX1 U9155 ( .A(n20095), .Y(n20004) );
  NAND2X1 U9156 ( .A(n22447), .B(n22481), .Y(n22761) );
  NAND2X1 U9157 ( .A(n13527), .B(n24441), .Y(n24881) );
  INVX1 U9158 ( .A(n25048), .Y(n25070) );
  INVX1 U9159 ( .A(n14002), .Y(n24461) );
  NAND2BX2 U9160 ( .AN(n7158), .B(n6104), .Y(n20015) );
  INVXL U9161 ( .A(n17098), .Y(n7515) );
  CLKINVX3 U9162 ( .A(n24663), .Y(n24641) );
  NAND2X1 U9163 ( .A(n6452), .B(n12257), .Y(n6451) );
  NAND2X1 U9164 ( .A(n20002), .B(n6033), .Y(n17104) );
  AND2XL U9165 ( .A(n5867), .B(n19282), .Y(n8144) );
  AOI21X1 U9166 ( .A0(n12968), .A1(n12967), .B0(n12966), .Y(n17667) );
  NAND2XL U9167 ( .A(n19750), .B(n19872), .Y(n6688) );
  OR2X2 U9168 ( .A(n24661), .B(n24643), .Y(n25018) );
  NAND2XL U9169 ( .A(n24646), .B(n14553), .Y(n25363) );
  INVX1 U9170 ( .A(n17638), .Y(n17633) );
  NAND2X1 U9171 ( .A(n19987), .B(n12970), .Y(n7018) );
  MXI2X1 U9172 ( .A(U2_pipe2[7]), .B(n20757), .S0(n21023), .Y(n4161) );
  MXI2X1 U9173 ( .A(U2_pipe2[6]), .B(n20702), .S0(n21023), .Y(n4159) );
  INVX1 U9174 ( .A(n17526), .Y(n17555) );
  MXI2X1 U9175 ( .A(U2_pipe3[6]), .B(n17984), .S0(n8054), .Y(n4211) );
  INVX1 U9176 ( .A(n24919), .Y(n24941) );
  INVX1 U9177 ( .A(n19152), .Y(n19184) );
  INVXL U9178 ( .A(n6258), .Y(n6254) );
  MXI2X1 U9179 ( .A(U2_pipe1[10]), .B(n23581), .S0(n23695), .Y(n4115) );
  MXI2X1 U9180 ( .A(U2_pipe1[9]), .B(n23531), .S0(n23695), .Y(n4113) );
  MXI2X1 U9181 ( .A(U2_pipe1[7]), .B(n23435), .S0(n23695), .Y(n4109) );
  INVXL U9182 ( .A(n24786), .Y(n25051) );
  NAND2XL U9183 ( .A(n14482), .B(U2_A_r_d[22]), .Y(n7041) );
  INVX1 U9184 ( .A(n24503), .Y(n24535) );
  INVX2 U9185 ( .A(n14548), .Y(n12388) );
  OR2X2 U9186 ( .A(n24620), .B(n24631), .Y(n9004) );
  OAI21XL U9187 ( .A0(n19873), .A1(n19748), .B0(n19747), .Y(n19749) );
  MXI2X1 U9188 ( .A(U2_pipe2[5]), .B(n20656), .S0(n21023), .Y(n4157) );
  INVX1 U9189 ( .A(n22492), .Y(n5818) );
  INVX1 U9190 ( .A(n21886), .Y(n22116) );
  MXI2X1 U9191 ( .A(U2_pipe1[5]), .B(n23328), .S0(n23695), .Y(n4105) );
  INVX1 U9192 ( .A(n17232), .Y(n17257) );
  INVX1 U9193 ( .A(n6580), .Y(n17016) );
  NAND2X1 U9194 ( .A(n18980), .B(n18979), .Y(n6258) );
  INVX1 U9195 ( .A(n23741), .Y(n23794) );
  CLKINVX3 U9196 ( .A(n14929), .Y(n19987) );
  MXI2X1 U9197 ( .A(U2_pipe1[6]), .B(n23371), .S0(n23695), .Y(n4107) );
  AOI21XL U9198 ( .A0(n18812), .A1(n18811), .B0(n18810), .Y(n18813) );
  MXI2X1 U9199 ( .A(U2_pipe1[8]), .B(n23487), .S0(n23695), .Y(n4111) );
  MXI2X1 U9200 ( .A(U2_pipe0[7]), .B(n26087), .S0(n8054), .Y(n4057) );
  INVXL U9201 ( .A(n14547), .Y(n5864) );
  NAND2BX1 U9202 ( .AN(n14955), .B(n19272), .Y(n17638) );
  OR2X2 U9203 ( .A(n14950), .B(n19541), .Y(n13554) );
  INVX2 U9204 ( .A(n24646), .Y(n5820) );
  NAND2BXL U9205 ( .AN(n5880), .B(n7885), .Y(n19304) );
  AOI21X1 U9206 ( .A0(n6633), .A1(n5792), .B0(n6669), .Y(n6668) );
  NAND2X1 U9207 ( .A(n7727), .B(n5894), .Y(n6309) );
  NAND2XL U9208 ( .A(n12963), .B(n19330), .Y(n17680) );
  AOI21X1 U9209 ( .A0(n22707), .A1(n12528), .B0(n12527), .Y(n22687) );
  NAND2X1 U9210 ( .A(n13082), .B(n5892), .Y(n6152) );
  NAND2X2 U9211 ( .A(n5991), .B(n5936), .Y(n5935) );
  INVX1 U9212 ( .A(n21189), .Y(n20958) );
  INVX1 U9213 ( .A(n25189), .Y(n14445) );
  CLKINVX3 U9214 ( .A(n19980), .Y(n14926) );
  INVX1 U9215 ( .A(n13506), .Y(n24509) );
  NAND2XL U9216 ( .A(n7907), .B(n7911), .Y(n7910) );
  INVX1 U9217 ( .A(n14530), .Y(n14535) );
  NOR2X1 U9218 ( .A(n20005), .B(n19544), .Y(n19620) );
  AND2X1 U9219 ( .A(n19758), .B(U1_A_r_d0[14]), .Y(n19759) );
  MXI2X1 U9220 ( .A(U2_pipe0[6]), .B(n26041), .S0(n8054), .Y(n4055) );
  INVX1 U9221 ( .A(n16889), .Y(n16907) );
  NAND2X1 U9222 ( .A(n14930), .B(n5880), .Y(n20113) );
  NAND2X1 U9223 ( .A(n19977), .B(n19976), .Y(n20117) );
  OR2X2 U9224 ( .A(n14940), .B(n14930), .Y(n13881) );
  INVX1 U9225 ( .A(n25193), .Y(n14444) );
  XOR2X1 U9226 ( .A(n27035), .B(n21698), .Y(n21699) );
  NAND2X1 U9227 ( .A(n7441), .B(n7442), .Y(n7440) );
  OR2X2 U9228 ( .A(n14923), .B(n14902), .Y(n13801) );
  NAND2X1 U9229 ( .A(n21311), .B(n21310), .Y(n21416) );
  AND2XL U9230 ( .A(n5880), .B(n19311), .Y(n8146) );
  NOR2X1 U9231 ( .A(n21175), .B(n21180), .Y(n21183) );
  AND2X2 U9232 ( .A(n13973), .B(n13975), .Y(n7011) );
  INVX1 U9233 ( .A(n24327), .Y(n24328) );
  INVX1 U9234 ( .A(n14073), .Y(n13398) );
  CLKINVX3 U9235 ( .A(n6048), .Y(n5990) );
  XOR2X1 U9236 ( .A(n24375), .B(n18985), .Y(n18986) );
  NAND2X1 U9237 ( .A(n5985), .B(n13032), .Y(n13024) );
  AND2XL U9238 ( .A(n5876), .B(U2_A_r_d[11]), .Y(n24506) );
  OR2XL U9239 ( .A(n27035), .B(n27034), .Y(n27037) );
  INVX1 U9240 ( .A(n26986), .Y(n26987) );
  CLKINVX3 U9241 ( .A(n7786), .Y(n6044) );
  INVX1 U9242 ( .A(n18770), .Y(n6417) );
  INVX1 U9243 ( .A(n26904), .Y(n26905) );
  NAND2X1 U9244 ( .A(n6226), .B(n14821), .Y(n7224) );
  NAND2X1 U9245 ( .A(n12189), .B(n12208), .Y(n12190) );
  XNOR2X2 U9246 ( .A(n13869), .B(n13868), .Y(n14927) );
  NOR2X1 U9247 ( .A(n21073), .B(n21072), .Y(n21175) );
  MXI2X1 U9248 ( .A(Q7[25]), .B(n18994), .S0(U1_valid[1]), .Y(n3934) );
  INVX1 U9249 ( .A(n13963), .Y(n13969) );
  NOR2X1 U9250 ( .A(n20962), .B(n20961), .Y(n21063) );
  NAND2X1 U9251 ( .A(n13019), .B(n5896), .Y(n5985) );
  NAND2BX1 U9252 ( .AN(n6000), .B(n5879), .Y(n6702) );
  INVX1 U9253 ( .A(n8575), .Y(n8584) );
  MXI2X1 U9254 ( .A(Q2[25]), .B(n24394), .S0(n23239), .Y(n3597) );
  NAND2X1 U9255 ( .A(n14816), .B(n5897), .Y(n6226) );
  MXI2X1 U9256 ( .A(Q5[53]), .B(n21729), .S0(n23239), .Y(n3987) );
  INVXL U9257 ( .A(n14840), .Y(n7890) );
  MXI2X1 U9258 ( .A(Q2[53]), .B(n27056), .S0(n24128), .Y(n3623) );
  INVX1 U9259 ( .A(n23480), .Y(n23364) );
  NAND2X1 U9260 ( .A(n26993), .B(n26992), .Y(n27029) );
  NAND2X1 U9261 ( .A(n18713), .B(n18712), .Y(n18808) );
  INVX1 U9262 ( .A(n18769), .Y(n6416) );
  NAND2X1 U9263 ( .A(n5878), .B(n13057), .Y(n6075) );
  INVX1 U9264 ( .A(n7641), .Y(n7639) );
  NAND2X1 U9265 ( .A(n24334), .B(n24333), .Y(n24370) );
  MXI2X1 U9266 ( .A(Q7[53]), .B(n21708), .S0(n23239), .Y(n3908) );
  INVX1 U9267 ( .A(n13905), .Y(n7837) );
  NAND2X2 U9268 ( .A(n7840), .B(n7841), .Y(n5959) );
  OR2X2 U9269 ( .A(n24163), .B(n24162), .Y(n24161) );
  NOR2XL U9270 ( .A(n13583), .B(n7834), .Y(n7833) );
  AOI21X1 U9271 ( .A0(n9062), .A1(n8961), .B0(n8941), .Y(n8946) );
  INVX1 U9272 ( .A(n7667), .Y(n7665) );
  INVX1 U9273 ( .A(n13967), .Y(n13968) );
  MXI2X1 U9274 ( .A(Q6[53]), .B(n21715), .S0(n23239), .Y(n3856) );
  INVX1 U9275 ( .A(n25231), .Y(n14380) );
  MXI2X1 U9276 ( .A(Q3[25]), .B(n24387), .S0(n24128), .Y(n3545) );
  AND2X2 U9277 ( .A(n12259), .B(n12262), .Y(n6926) );
  MXI2X1 U9278 ( .A(Q4[53]), .B(n21722), .S0(n24128), .Y(n4050) );
  NAND2X1 U9279 ( .A(n7278), .B(n13600), .Y(n13576) );
  MXI2X1 U9280 ( .A(Q1[25]), .B(n24408), .S0(n23239), .Y(n3466) );
  NAND2X1 U9281 ( .A(n7176), .B(n13566), .Y(n7175) );
  NAND2X1 U9282 ( .A(n12267), .B(n12271), .Y(n12268) );
  NAND2X1 U9283 ( .A(n12283), .B(n12355), .Y(n12284) );
  MXI2X1 U9284 ( .A(Q0[25]), .B(n24401), .S0(n24128), .Y(n3518) );
  MXI2X1 U9285 ( .A(Q1[53]), .B(n27070), .S0(n23239), .Y(n3492) );
  MXI2X1 U9286 ( .A(Q0[53]), .B(n27063), .S0(n23239), .Y(n3429) );
  INVXL U9287 ( .A(n14839), .Y(n7889) );
  MXI2X1 U9288 ( .A(Q3[53]), .B(n27049), .S0(n23239), .Y(n3571) );
  ADDFHX1 U9289 ( .A(n21362), .B(n21361), .CI(U2_A_r_d[17]), .CO(n21363), .S(
        n21311) );
  NAND2XL U9290 ( .A(n6442), .B(n5893), .Y(n6437) );
  NAND2X1 U9291 ( .A(n12274), .B(n12278), .Y(n12277) );
  AND2X2 U9292 ( .A(n14681), .B(n14849), .Y(n6966) );
  AND2X2 U9293 ( .A(n13634), .B(n13644), .Y(n7003) );
  INVXL U9294 ( .A(n26909), .Y(n21574) );
  INVX1 U9295 ( .A(n21694), .Y(n21695) );
  AND2X2 U9296 ( .A(n6849), .B(n9219), .Y(n6848) );
  NOR2XL U9297 ( .A(n14797), .B(n7891), .Y(n7160) );
  NAND2X1 U9298 ( .A(n18496), .B(n18497), .Y(n18593) );
  NAND2X1 U9299 ( .A(n13054), .B(n13072), .Y(n13055) );
  ADDFHX2 U9300 ( .A(n21122), .B(n21121), .CI(U2_A_r_d[13]), .CO(n21123), .S(
        n21073) );
  NAND2X1 U9301 ( .A(n13606), .B(n13605), .Y(n13614) );
  INVX1 U9302 ( .A(n19732), .Y(n8657) );
  OR2X2 U9303 ( .A(n19520), .B(n19969), .Y(n19505) );
  NAND2X1 U9304 ( .A(n14860), .B(n14859), .Y(n14861) );
  AND2X2 U9305 ( .A(n13986), .B(n13989), .Y(n6957) );
  INVX1 U9306 ( .A(n12278), .Y(n12279) );
  NOR2X1 U9307 ( .A(n18497), .B(n18496), .Y(n18591) );
  NAND2X1 U9308 ( .A(n9484), .B(n9483), .Y(n9485) );
  INVX1 U9309 ( .A(n9034), .Y(n9150) );
  INVX4 U9310 ( .A(n9189), .Y(n5821) );
  NOR2X1 U9311 ( .A(n26191), .B(n26190), .Y(n26238) );
  NAND2X1 U9312 ( .A(n26463), .B(n26462), .Y(n26595) );
  INVX1 U9313 ( .A(n13950), .Y(n5937) );
  CLKINVX3 U9314 ( .A(n7888), .Y(n5882) );
  INVXL U9315 ( .A(n13954), .Y(n6481) );
  AND2X2 U9316 ( .A(n13932), .B(n13951), .Y(n6978) );
  NAND2XL U9317 ( .A(n6931), .B(n7922), .Y(n7921) );
  INVX1 U9318 ( .A(n18981), .Y(n18982) );
  AND2XL U9319 ( .A(n9072), .B(n9165), .Y(n7228) );
  NAND2X1 U9320 ( .A(n13965), .B(n13964), .Y(n13967) );
  NAND2XL U9321 ( .A(n6931), .B(n13580), .Y(n7834) );
  INVX1 U9322 ( .A(n8619), .Y(n6669) );
  NAND2X1 U9323 ( .A(n13940), .B(n13939), .Y(n13941) );
  NAND2X2 U9324 ( .A(n6133), .B(n6008), .Y(n7802) );
  NAND3X1 U9325 ( .A(n7831), .B(n7832), .C(n5949), .Y(n5948) );
  NAND2X1 U9326 ( .A(n9190), .B(n9201), .Y(n9193) );
  INVXL U9327 ( .A(n14463), .Y(n6521) );
  AND2X2 U9328 ( .A(n5892), .B(n13080), .Y(n7004) );
  INVX1 U9329 ( .A(n25235), .Y(n21758) );
  NOR2X1 U9330 ( .A(n20698), .B(n20697), .Y(n20744) );
  OAI21X1 U9331 ( .A0(n7827), .A1(n12891), .B0(n6007), .Y(n12781) );
  INVX1 U9332 ( .A(n13938), .Y(n13940) );
  INVX1 U9333 ( .A(n13796), .Y(n13791) );
  NAND2X1 U9334 ( .A(n8565), .B(n8567), .Y(n8566) );
  INVX1 U9335 ( .A(n13073), .Y(n13051) );
  NAND2X1 U9336 ( .A(n5889), .B(n9185), .Y(n9160) );
  AND2X2 U9337 ( .A(n5890), .B(n8622), .Y(n8623) );
  NAND2BXL U9338 ( .AN(n9220), .B(n9202), .Y(n6849) );
  INVX1 U9339 ( .A(n26356), .Y(n21017) );
  CLKINVX3 U9340 ( .A(n26290), .Y(n20959) );
  INVX1 U9341 ( .A(n13591), .Y(n5884) );
  INVXL U9342 ( .A(n13578), .Y(n7506) );
  OR2X2 U9343 ( .A(n12261), .B(n12260), .Y(n12259) );
  INVX1 U9344 ( .A(n9154), .Y(n9033) );
  NAND2X1 U9345 ( .A(n12261), .B(n12260), .Y(n12262) );
  INVX1 U9346 ( .A(n13164), .Y(n13173) );
  OAI2BB1X2 U9347 ( .A0N(n14774), .A1N(n14657), .B0(n6131), .Y(n7886) );
  NAND2X1 U9348 ( .A(n13164), .B(n13172), .Y(n13165) );
  AND2X2 U9349 ( .A(n13628), .B(n13637), .Y(n6967) );
  INVX1 U9350 ( .A(n14845), .Y(n6125) );
  NAND2X1 U9351 ( .A(n12276), .B(n12275), .Y(n12278) );
  NOR2X1 U9352 ( .A(n14794), .B(n14798), .Y(n14674) );
  AND2X2 U9353 ( .A(n9475), .B(n9474), .Y(n6919) );
  NAND2X1 U9354 ( .A(n9428), .B(n9427), .Y(n9429) );
  AND2X2 U9355 ( .A(n9527), .B(n9526), .Y(n6961) );
  XOR2X1 U9356 ( .A(n14768), .B(n14705), .Y(n19969) );
  NAND2X1 U9357 ( .A(n13636), .B(n13635), .Y(n13644) );
  INVXL U9358 ( .A(n13041), .Y(n7172) );
  INVX1 U9359 ( .A(n12082), .Y(n12077) );
  NOR2X1 U9360 ( .A(n20653), .B(n20652), .Y(n20740) );
  NOR2X1 U9361 ( .A(n17941), .B(n17940), .Y(n18040) );
  AOI21X1 U9362 ( .A0(n5988), .A1(n14764), .B0(n14759), .Y(n7812) );
  OR2X2 U9363 ( .A(n14683), .B(n14682), .Y(n14681) );
  AND2X2 U9364 ( .A(n14811), .B(n14810), .Y(n6968) );
  XOR2X1 U9365 ( .A(n14688), .B(n14687), .Y(n14689) );
  AND2X2 U9366 ( .A(n5896), .B(n13032), .Y(n13033) );
  NAND2X1 U9367 ( .A(n14686), .B(n14685), .Y(n14859) );
  NAND2X1 U9368 ( .A(n7898), .B(n14805), .Y(n14806) );
  NAND2X1 U9369 ( .A(n13867), .B(n13866), .Y(n13868) );
  INVX1 U9370 ( .A(n7522), .Y(n6007) );
  INVX1 U9371 ( .A(n26189), .Y(n20855) );
  NOR2X1 U9372 ( .A(n9422), .B(n9420), .Y(n9438) );
  AND2X2 U9373 ( .A(n8633), .B(n8632), .Y(n6964) );
  NAND2X1 U9374 ( .A(n5897), .B(n14821), .Y(n14822) );
  INVX1 U9375 ( .A(n9468), .Y(n9470) );
  NAND2X1 U9376 ( .A(n8149), .B(n8624), .Y(n8625) );
  NAND2X1 U9377 ( .A(n7884), .B(n14777), .Y(n14778) );
  INVX1 U9378 ( .A(n9420), .Y(n9428) );
  INVX1 U9379 ( .A(n9427), .Y(n9421) );
  AND2X1 U9380 ( .A(n9126), .B(n9125), .Y(n6940) );
  NAND2X1 U9381 ( .A(n13641), .B(n13640), .Y(n13652) );
  NAND2X1 U9382 ( .A(n12569), .B(n12584), .Y(n12570) );
  AND2X2 U9383 ( .A(n13018), .B(n13017), .Y(n6896) );
  INVXL U9384 ( .A(n7726), .Y(n6376) );
  NAND2X1 U9385 ( .A(n12072), .B(n12079), .Y(n12073) );
  INVXL U9386 ( .A(n13914), .Y(n7432) );
  NAND2X1 U9387 ( .A(n5893), .B(n12343), .Y(n9230) );
  NAND2X1 U9388 ( .A(n12164), .B(n12178), .Y(n12165) );
  NAND2X1 U9389 ( .A(n13174), .B(n13179), .Y(n13177) );
  NAND2X1 U9390 ( .A(n5894), .B(n9091), .Y(n9092) );
  NAND2X1 U9391 ( .A(n5898), .B(n12157), .Y(n12145) );
  NAND2BX1 U9392 ( .AN(n13163), .B(n6449), .Y(n13164) );
  NAND2XL U9393 ( .A(n13930), .B(n13931), .Y(n13951) );
  AND2X2 U9394 ( .A(n9073), .B(n9152), .Y(n6973) );
  INVX1 U9395 ( .A(n13949), .Y(n5822) );
  NAND2X2 U9396 ( .A(n13924), .B(n13925), .Y(n13939) );
  INVX1 U9397 ( .A(n13179), .Y(n13180) );
  NOR2X1 U9398 ( .A(n13586), .B(n13587), .Y(n13591) );
  INVX1 U9399 ( .A(n14479), .Y(n14269) );
  INVX1 U9400 ( .A(n13474), .Y(n13288) );
  NAND2X1 U9401 ( .A(n5895), .B(n9128), .Y(n9129) );
  OR2X2 U9402 ( .A(n24588), .B(n13099), .Y(n12118) );
  NAND2X1 U9403 ( .A(n13903), .B(n13902), .Y(n13921) );
  OR2X2 U9404 ( .A(n13597), .B(n13596), .Y(n13595) );
  NAND2X1 U9405 ( .A(n13597), .B(n13596), .Y(n13607) );
  INVX1 U9406 ( .A(n11462), .Y(n11476) );
  NOR2X1 U9407 ( .A(n11483), .B(n11490), .Y(n11455) );
  AND2XL U9408 ( .A(n19709), .B(U1_A_r_d0[0]), .Y(n20304) );
  INVX1 U9409 ( .A(n9152), .Y(n9037) );
  NAND2X1 U9410 ( .A(n13157), .B(n13156), .Y(n13159) );
  NAND2X1 U9411 ( .A(n13183), .B(n13182), .Y(n13186) );
  NAND2X1 U9412 ( .A(n13287), .B(n13286), .Y(n13474) );
  NAND2X1 U9413 ( .A(n13176), .B(n13175), .Y(n13179) );
  OR2X2 U9414 ( .A(n14907), .B(n19952), .Y(n13833) );
  NAND2X1 U9415 ( .A(n13293), .B(n13292), .Y(n13483) );
  NAND2X1 U9416 ( .A(n9192), .B(n9191), .Y(n9201) );
  OR2X2 U9417 ( .A(n9223), .B(n9222), .Y(n9221) );
  NAND2X1 U9418 ( .A(n9223), .B(n9222), .Y(n9231) );
  NAND2X1 U9419 ( .A(n9235), .B(n9234), .Y(n12348) );
  OR2X2 U9420 ( .A(n9182), .B(n9181), .Y(n9180) );
  NAND2X1 U9421 ( .A(n8454), .B(n8453), .Y(n8627) );
  NAND2BX1 U9422 ( .AN(n8456), .B(n6522), .Y(n8633) );
  NAND2X1 U9423 ( .A(n8750), .B(n8822), .Y(n8751) );
  INVX1 U9424 ( .A(n8990), .Y(n8963) );
  NAND2X1 U9425 ( .A(n13028), .B(n13027), .Y(n13029) );
  NAND2X1 U9426 ( .A(n12645), .B(n12644), .Y(n13136) );
  NOR2X1 U9427 ( .A(n9159), .B(n9158), .Y(n9186) );
  AND2X2 U9428 ( .A(n5901), .B(n8823), .Y(n8817) );
  NAND2X1 U9429 ( .A(n12628), .B(n12629), .Y(n12639) );
  AOI21X1 U9430 ( .A0(n19064), .A1(n19063), .B0(n19062), .Y(n25845) );
  INVX1 U9431 ( .A(n12156), .Y(n12146) );
  INVX1 U9432 ( .A(n14429), .Y(n14431) );
  AND2X2 U9433 ( .A(n8529), .B(n8528), .Y(n6925) );
  INVX1 U9434 ( .A(n14438), .Y(n14433) );
  INVX1 U9435 ( .A(n12158), .Y(n12142) );
  NOR2X1 U9436 ( .A(n14271), .B(n14270), .Y(n14491) );
  NAND2X1 U9437 ( .A(n14271), .B(n14270), .Y(n14492) );
  INVXL U9438 ( .A(n23429), .Y(n18052) );
  NAND2X1 U9439 ( .A(n14268), .B(n14267), .Y(n14479) );
  INVX1 U9440 ( .A(n23481), .Y(n18092) );
  NAND2X1 U9441 ( .A(n12768), .B(n12787), .Y(n12769) );
  AOI21X1 U9442 ( .A0(n16623), .A1(n16622), .B0(n16621), .Y(n23174) );
  AND2XL U9443 ( .A(n19709), .B(U1_A_i_d0[0]), .Y(n17046) );
  NAND2BXL U9444 ( .AN(n9352), .B(n9350), .Y(n7659) );
  NOR2X1 U9445 ( .A(n14265), .B(n14264), .Y(n14473) );
  INVX1 U9446 ( .A(n23576), .Y(n18188) );
  OR2X2 U9447 ( .A(n14262), .B(n14261), .Y(n14260) );
  NAND2X1 U9448 ( .A(n14262), .B(n14261), .Y(n14470) );
  INVX1 U9449 ( .A(n14020), .Y(n14061) );
  NAND2X1 U9450 ( .A(n7933), .B(n12937), .Y(n12899) );
  INVX1 U9451 ( .A(n13871), .Y(n13855) );
  NAND2X1 U9452 ( .A(n12924), .B(n12923), .Y(n12925) );
  NOR2X1 U9453 ( .A(n11456), .B(U2_B_r[24]), .Y(n11462) );
  NAND2X1 U9454 ( .A(n14258), .B(n14257), .Y(n14466) );
  NAND2X1 U9455 ( .A(n11456), .B(U2_B_r[24]), .Y(n11475) );
  NAND2X1 U9456 ( .A(n14244), .B(n14243), .Y(n14398) );
  NAND2X1 U9457 ( .A(n12953), .B(n12952), .Y(n12994) );
  BUFX4 U9458 ( .A(B2_addr[3]), .Y(n7135) );
  XOR2X1 U9459 ( .A(n9393), .B(n9392), .Y(n13665) );
  NAND2X1 U9460 ( .A(n7044), .B(n14656), .Y(n14777) );
  NOR2X1 U9461 ( .A(n9063), .B(n9064), .Y(n9090) );
  XOR2X1 U9462 ( .A(n13830), .B(n13829), .Y(n14905) );
  XOR2X1 U9463 ( .A(U0_U1_y0[40]), .B(U0_U1_y2[40]), .Y(n13190) );
  XNOR2X1 U9464 ( .A(n13841), .B(n13840), .Y(n14911) );
  NAND2X1 U9465 ( .A(n9036), .B(n9035), .Y(n9152) );
  AOI211XL U9466 ( .A0(n5918), .A1(n28544), .B0(n28543), .C0(n28542), .Y(
        n28545) );
  NAND2X1 U9467 ( .A(n12985), .B(n12984), .Y(n13017) );
  NOR2X1 U9468 ( .A(n13783), .B(n13784), .Y(n13792) );
  AND2X2 U9469 ( .A(n5902), .B(n12474), .Y(n12471) );
  INVX1 U9470 ( .A(n13364), .Y(n13371) );
  INVX1 U9471 ( .A(n8581), .Y(n5900) );
  NAND2X1 U9472 ( .A(n13280), .B(n13279), .Y(n13433) );
  NAND2X1 U9473 ( .A(n13284), .B(n13283), .Y(n13471) );
  XOR2X1 U9474 ( .A(U0_U0_y0[40]), .B(U0_U0_y1[40]), .Y(n13298) );
  XOR2X1 U9475 ( .A(n8873), .B(n8872), .Y(n24851) );
  CLKINVX3 U9476 ( .A(n8953), .Y(n8897) );
  NOR2X1 U9477 ( .A(n12544), .B(n12543), .Y(n12559) );
  XOR2X1 U9478 ( .A(n14730), .B(n14729), .Y(n20179) );
  XOR2X1 U9479 ( .A(n12855), .B(n12854), .Y(n19507) );
  XOR2X1 U9480 ( .A(n12115), .B(n12114), .Y(n13098) );
  INVX1 U9481 ( .A(n8475), .Y(n8472) );
  AOI211XL U9482 ( .A0(n5918), .A1(n27744), .B0(n28557), .C0(n27743), .Y(
        n27745) );
  XOR2X1 U9483 ( .A(n8507), .B(n8506), .Y(n19709) );
  OR2X2 U9484 ( .A(n19954), .B(n19952), .Y(n14866) );
  NAND2X1 U9485 ( .A(n14771), .B(n14770), .Y(n14772) );
  INVXL U9486 ( .A(n23322), .Y(n17939) );
  XOR2X1 U9487 ( .A(U0_U0_y0[40]), .B(U0_U0_y2[40]), .Y(n14273) );
  AND2X2 U9488 ( .A(n14762), .B(n14761), .Y(n6921) );
  INVXL U9489 ( .A(n11540), .Y(n6177) );
  NOR2X1 U9490 ( .A(n12141), .B(n12140), .Y(n12156) );
  OAI21X1 U9491 ( .A0(n14760), .A1(n14763), .B0(n14761), .Y(n14774) );
  INVX1 U9492 ( .A(n10519), .Y(n8236) );
  NAND2X1 U9493 ( .A(n28630), .B(n11975), .Y(n28635) );
  XOR2X1 U9494 ( .A(U1_U2_y2[26]), .B(U1_U2_y0[26]), .Y(n7839) );
  CLKINVX3 U9495 ( .A(U2_B_i[18]), .Y(n11445) );
  AND2X2 U9496 ( .A(U1_U2_y2[26]), .B(U1_U2_y0[26]), .Y(n5934) );
  INVX1 U9497 ( .A(n14349), .Y(n14356) );
  INVX1 U9498 ( .A(U2_B_i[24]), .Y(n11456) );
  NAND2X1 U9499 ( .A(U2_B_r[19]), .B(n11446), .Y(n11508) );
  NAND2X1 U9500 ( .A(n12898), .B(n12897), .Y(n12937) );
  NOR2X1 U9501 ( .A(n11995), .B(n29241), .Y(A0_CEN) );
  NAND2X1 U9502 ( .A(n14240), .B(n14239), .Y(n14411) );
  NAND2X1 U9503 ( .A(n13780), .B(n13779), .Y(n13813) );
  NOR2X1 U9504 ( .A(n11995), .B(n11994), .Y(A4_CEN) );
  XOR2X1 U9505 ( .A(n8514), .B(n8509), .Y(n12288) );
  NAND2X1 U9506 ( .A(n12943), .B(n12942), .Y(n12976) );
  NAND2X1 U9507 ( .A(n12467), .B(n12466), .Y(n12473) );
  NAND2X1 U9508 ( .A(n8749), .B(n8748), .Y(n8822) );
  NAND2X1 U9509 ( .A(n8466), .B(n8465), .Y(n8467) );
  XOR2X1 U9510 ( .A(U1_U0_y0[40]), .B(U1_U0_y2[40]), .Y(n8460) );
  XOR2X1 U9511 ( .A(U0_U1_y0[40]), .B(U0_U1_y1[40]), .Y(n12346) );
  NAND2X1 U9512 ( .A(n8813), .B(n8812), .Y(n8831) );
  XOR2X1 U9513 ( .A(n14740), .B(n14732), .Y(n19954) );
  NAND2X1 U9514 ( .A(n13306), .B(n13305), .Y(n7009) );
  NOR2X1 U9515 ( .A(n14760), .B(n14758), .Y(n14775) );
  NAND2X1 U9516 ( .A(n13325), .B(n13324), .Y(n13326) );
  NAND2X1 U9517 ( .A(n8427), .B(n8428), .Y(n8544) );
  NAND2X1 U9518 ( .A(n8836), .B(n8835), .Y(n8971) );
  INVX1 U9519 ( .A(U2_B_i[19]), .Y(n11446) );
  INVXL U9520 ( .A(U2_B_i[15]), .Y(n11439) );
  INVX1 U9521 ( .A(U2_B_i[21]), .Y(n11451) );
  INVX1 U9522 ( .A(n7107), .Y(n7108) );
  INVX1 U9523 ( .A(n7097), .Y(n7098) );
  NOR2X2 U9524 ( .A(n12062), .B(n12063), .Y(n12092) );
  INVX1 U9525 ( .A(n7105), .Y(n7106) );
  INVXL U9526 ( .A(U0_U2_y2[23]), .Y(n6430) );
  NOR2X2 U9527 ( .A(n12761), .B(n12762), .Y(n12813) );
  INVX1 U9528 ( .A(U0_U2_y0[23]), .Y(n6431) );
  INVX4 U9529 ( .A(n5799), .Y(n16559) );
  NOR2X1 U9530 ( .A(n11993), .B(n11992), .Y(n11995) );
  NAND2X1 U9531 ( .A(n6513), .B(n6512), .Y(n9350) );
  CMPR22X1 U9532 ( .A(U1_U1_y2[22]), .B(U1_U1_y0[22]), .CO(n12895), .S(n12892)
         );
  CLKINVX3 U9533 ( .A(n27088), .Y(n28055) );
  INVX1 U9534 ( .A(n7091), .Y(n7092) );
  INVX1 U9535 ( .A(n7093), .Y(n7094) );
  NOR2X1 U9536 ( .A(n14651), .B(n14650), .Y(n14758) );
  OAI21X2 U9537 ( .A0(n6330), .A1(n29106), .B0(n11423), .Y(U2_B_i[24]) );
  INVX8 U9538 ( .A(n11900), .Y(B1_addr[6]) );
  INVX1 U9539 ( .A(n18747), .Y(n18682) );
  NAND2X1 U9540 ( .A(n11650), .B(n11649), .Y(T1_rom_addr[6]) );
  INVX1 U9541 ( .A(n21459), .Y(n21395) );
  INVX1 U9542 ( .A(n26797), .Y(n26735) );
  INVX1 U9543 ( .A(n11880), .Y(n11881) );
  INVX1 U9544 ( .A(n18734), .Y(n18671) );
  XOR2X2 U9545 ( .A(n6405), .B(n10055), .Y(U2_U0_z2[9]) );
  NAND3X1 U9546 ( .A(n7744), .B(n7262), .C(n7743), .Y(n6171) );
  NAND2X1 U9547 ( .A(n9623), .B(n7088), .Y(n11587) );
  INVX8 U9548 ( .A(n27205), .Y(n5823) );
  INVX1 U9549 ( .A(n24148), .Y(n24062) );
  INVX1 U9550 ( .A(n24136), .Y(n24073) );
  CMPR22X1 U9551 ( .A(U1_U0_y1[18]), .B(U1_U0_y0[18]), .CO(n9301), .S(n9296)
         );
  NOR2X2 U9552 ( .A(n14644), .B(n14645), .Y(n14692) );
  INVX1 U9553 ( .A(n18759), .Y(n18693) );
  INVX1 U9554 ( .A(n24123), .Y(n24084) );
  AOI21X1 U9555 ( .A0(n11214), .A1(n11213), .B0(n11212), .Y(n11215) );
  CMPR22X1 U9556 ( .A(U1_U1_y1[22]), .B(U1_U1_y0[22]), .CO(n14651), .S(n14648)
         );
  NAND2X1 U9557 ( .A(n8313), .B(U2_B_r[4]), .Y(n11583) );
  INVX1 U9558 ( .A(n7085), .Y(n7086) );
  CLKINVX3 U9559 ( .A(n5924), .Y(n6880) );
  CMPR22X1 U9560 ( .A(U1_U1_y1[19]), .B(U1_U1_y0[19]), .CO(n14645), .S(n14642)
         );
  NAND2X1 U9561 ( .A(n8412), .B(n8411), .Y(n8485) );
  INVX4 U9562 ( .A(n5924), .Y(n5909) );
  CLKBUFX8 U9563 ( .A(n28050), .Y(n7140) );
  NOR2X1 U9564 ( .A(n8803), .B(n8802), .Y(n8845) );
  INVX1 U9565 ( .A(n7109), .Y(n7110) );
  AOI21XL U9566 ( .A0(n8797), .A1(n8875), .B0(n8796), .Y(n8798) );
  INVX4 U9567 ( .A(n5924), .Y(n5915) );
  NOR2X1 U9568 ( .A(n8738), .B(n8739), .Y(n8851) );
  INVX1 U9569 ( .A(U2_U0_y2[13]), .Y(n17752) );
  NOR2X1 U9570 ( .A(n11952), .B(n11874), .Y(n28661) );
  INVX1 U9571 ( .A(n7103), .Y(n7104) );
  INVX1 U9572 ( .A(n7101), .Y(n7102) );
  NOR2X1 U9573 ( .A(n14219), .B(n14218), .Y(n14282) );
  NAND2X1 U9574 ( .A(n12698), .B(n12699), .Y(n12818) );
  NAND2X1 U9575 ( .A(n14216), .B(n14215), .Y(n14299) );
  NAND2BX2 U9576 ( .AN(n11421), .B(n6331), .Y(n11425) );
  INVX1 U9577 ( .A(n7099), .Y(n7100) );
  INVX2 U9578 ( .A(U2_B_i[17]), .Y(n5824) );
  XOR2X1 U9579 ( .A(n6404), .B(BOPA[45]), .Y(n6403) );
  INVX1 U9580 ( .A(n7115), .Y(n7116) );
  INVX1 U9581 ( .A(n7111), .Y(n7112) );
  INVX1 U9582 ( .A(n7089), .Y(n7090) );
  INVX1 U9583 ( .A(n7113), .Y(n7114) );
  INVX1 U9584 ( .A(n11908), .Y(n28641) );
  NAND2X1 U9585 ( .A(n13245), .B(n13244), .Y(n13352) );
  NAND2X1 U9586 ( .A(n8801), .B(n8800), .Y(n8856) );
  NOR2X1 U9587 ( .A(n8801), .B(n8800), .Y(n8855) );
  OR2XL U9588 ( .A(n25101), .B(U0_pipe1[25]), .Y(n9238) );
  AOI21X1 U9589 ( .A0(n27976), .A1(Q1[37]), .B0(n27972), .Y(n28525) );
  NOR2X1 U9590 ( .A(n12455), .B(n12454), .Y(n12488) );
  NAND2X1 U9591 ( .A(n12455), .B(n12454), .Y(n12489) );
  NAND2X1 U9592 ( .A(n5921), .B(B_sel_reg[0]), .Y(n28050) );
  NOR2X1 U9593 ( .A(n12756), .B(n12755), .Y(n12872) );
  INVX4 U9594 ( .A(n11891), .Y(n5825) );
  AOI21X1 U9595 ( .A0(n27976), .A1(Q1[32]), .B0(n27951), .Y(n28490) );
  INVX1 U9596 ( .A(U0_U2_y0[16]), .Y(n6355) );
  NOR2X1 U9597 ( .A(n5922), .B(n28704), .Y(n27078) );
  NAND2X1 U9598 ( .A(n28964), .B(n7123), .Y(n27159) );
  NOR2X1 U9599 ( .A(n5922), .B(n28674), .Y(n27081) );
  NAND2X1 U9600 ( .A(n28983), .B(n7123), .Y(n27274) );
  NOR2X1 U9601 ( .A(n11984), .B(n28666), .Y(n11897) );
  OAI21X1 U9602 ( .A0(Q5[43]), .A1(n7123), .B0(n27237), .Y(n27752) );
  NAND2X1 U9603 ( .A(n28955), .B(n7123), .Y(n27123) );
  INVXL U9604 ( .A(n13827), .Y(n6068) );
  INVX1 U9605 ( .A(n10397), .Y(n10398) );
  NAND2X4 U9606 ( .A(n11929), .B(n28675), .Y(n27772) );
  NOR2X1 U9607 ( .A(n5922), .B(n28680), .Y(n27084) );
  NAND2X1 U9608 ( .A(n14210), .B(n14209), .Y(n14328) );
  NAND2X1 U9609 ( .A(n28967), .B(n7123), .Y(n27172) );
  NAND2X1 U9610 ( .A(n28969), .B(n7123), .Y(n27180) );
  NAND2X1 U9611 ( .A(n28968), .B(n7123), .Y(n27176) );
  NOR2X1 U9612 ( .A(n5922), .B(n28703), .Y(n15028) );
  NAND2X1 U9613 ( .A(n14214), .B(n14213), .Y(n14303) );
  NOR2X1 U9614 ( .A(n5922), .B(n28673), .Y(n14988) );
  NAND2X1 U9615 ( .A(n28957), .B(n7123), .Y(n27131) );
  NAND2X1 U9616 ( .A(n28956), .B(n7123), .Y(n27127) );
  NAND2X1 U9617 ( .A(n28984), .B(n7123), .Y(n27278) );
  NAND2X1 U9618 ( .A(n8406), .B(n8405), .Y(n8512) );
  NOR2X1 U9619 ( .A(n5922), .B(n28679), .Y(n27073) );
  CLKINVX3 U9620 ( .A(n11940), .Y(n5827) );
  NOR2X1 U9621 ( .A(n13775), .B(n13776), .Y(n13836) );
  NOR2X1 U9622 ( .A(n12694), .B(n12695), .Y(n12865) );
  NAND2X1 U9623 ( .A(n28976), .B(n7123), .Y(n27245) );
  NOR2X1 U9624 ( .A(n13774), .B(U1_U2_y2[13]), .Y(n13826) );
  CLKINVX3 U9625 ( .A(n7095), .Y(n7096) );
  INVX1 U9626 ( .A(n27950), .Y(n27951) );
  INVX1 U9627 ( .A(n27967), .Y(n27968) );
  INVX1 U9628 ( .A(n27855), .Y(n27856) );
  INVX1 U9629 ( .A(n9746), .Y(n9809) );
  NAND2X1 U9630 ( .A(n11427), .B(BOPA[15]), .Y(n8241) );
  INVX1 U9631 ( .A(n27815), .Y(n27816) );
  INVX1 U9632 ( .A(n7008), .Y(n6824) );
  INVX1 U9633 ( .A(n27958), .Y(n27960) );
  BUFX2 U9634 ( .A(n28284), .Y(n7120) );
  NAND2X1 U9635 ( .A(n11427), .B(BOPA[18]), .Y(n11402) );
  INVX1 U9636 ( .A(n27975), .Y(n27977) );
  NAND2X1 U9637 ( .A(n11427), .B(BOPA[24]), .Y(n11423) );
  OAI21X2 U9638 ( .A0(n28687), .A1(n11428), .B0(n11424), .Y(U2_B_r[24]) );
  NAND2X1 U9639 ( .A(n11427), .B(BOPA[19]), .Y(n11404) );
  INVX1 U9640 ( .A(n27954), .Y(n27955) );
  INVX1 U9641 ( .A(n27971), .Y(n27972) );
  NAND2X1 U9642 ( .A(n11427), .B(BOPA[17]), .Y(n8248) );
  NAND2X1 U9643 ( .A(n11427), .B(BOPA[25]), .Y(n11426) );
  XOR2X1 U9644 ( .A(n10690), .B(n10689), .Y(U1_U0_z0[2]) );
  NAND2X1 U9645 ( .A(n11427), .B(BOPA[16]), .Y(n11405) );
  NOR3X2 U9646 ( .A(n27236), .B(C_sel_reg[0]), .C(A_sel_reg[0]), .Y(n28322) );
  CLKINVX8 U9647 ( .A(n11709), .Y(n5828) );
  INVX8 U9648 ( .A(n5806), .Y(n16165) );
  INVX1 U9649 ( .A(n27835), .Y(n27836) );
  INVX4 U9650 ( .A(n11997), .Y(n5829) );
  INVX2 U9651 ( .A(n11956), .Y(n5830) );
  INVX1 U9652 ( .A(n27819), .Y(n27820) );
  INVX1 U9653 ( .A(n27851), .Y(n27852) );
  NAND2BX1 U9654 ( .AN(n8257), .B(n6159), .Y(n6158) );
  INVX1 U9655 ( .A(n27938), .Y(n27939) );
  INVX1 U9656 ( .A(n27823), .Y(n27824) );
  NOR2X1 U9657 ( .A(n8795), .B(U0_U1_y1[13]), .Y(n8884) );
  INVX1 U9658 ( .A(n10180), .Y(n7580) );
  CLKINVX8 U9659 ( .A(n11678), .Y(n5831) );
  CLKINVX8 U9660 ( .A(n11710), .Y(n5832) );
  INVX1 U9661 ( .A(n27839), .Y(n27840) );
  INVX1 U9662 ( .A(n27843), .Y(n27844) );
  INVX1 U9663 ( .A(n27827), .Y(n27828) );
  OR2XL U9664 ( .A(n6888), .B(U1_pipe6[26]), .Y(n7347) );
  INVX1 U9665 ( .A(n27946), .Y(n27947) );
  CLKINVX8 U9666 ( .A(n11684), .Y(n5833) );
  INVX1 U9667 ( .A(n27831), .Y(n27832) );
  AOI21X1 U9668 ( .A0(n27976), .A1(Q1[30]), .B0(n27943), .Y(n28476) );
  NAND2X1 U9669 ( .A(n10091), .B(n10093), .Y(n10096) );
  INVX1 U9670 ( .A(n11373), .Y(n11395) );
  OR2XL U9671 ( .A(U0_U2_y1[12]), .B(U0_U2_y0[12]), .Y(n8719) );
  NAND2X1 U9672 ( .A(n28973), .B(n5927), .Y(n27232) );
  AND2X2 U9673 ( .A(n10787), .B(n10786), .Y(n6918) );
  NAND2X1 U9674 ( .A(n10968), .B(n10967), .Y(n10969) );
  NAND2X1 U9675 ( .A(n10827), .B(n10826), .Y(n10828) );
  NAND2X1 U9676 ( .A(n10476), .B(n10475), .Y(n6916) );
  AND2XL U9677 ( .A(n11102), .B(n11101), .Y(n7010) );
  INVX1 U9678 ( .A(n10921), .Y(n10922) );
  AND2X2 U9679 ( .A(n11248), .B(n11247), .Y(n6960) );
  NAND2X1 U9680 ( .A(n10758), .B(n10757), .Y(n10759) );
  AND2X2 U9681 ( .A(n10552), .B(n10551), .Y(n6924) );
  NAND2X1 U9682 ( .A(n10984), .B(n10983), .Y(n10985) );
  AOI21XL U9683 ( .A0(n14592), .A1(n14591), .B0(n14590), .Y(n14593) );
  NAND2X1 U9684 ( .A(n8290), .B(n11092), .Y(n11080) );
  INVX4 U9685 ( .A(n17249), .Y(n17641) );
  NAND2X1 U9686 ( .A(n10717), .B(n10716), .Y(n10718) );
  NAND2X1 U9687 ( .A(n11057), .B(n11056), .Y(n11058) );
  NAND2X1 U9688 ( .A(n11120), .B(n8286), .Y(n8288) );
  AND2X2 U9689 ( .A(n9981), .B(n9980), .Y(n7008) );
  AND2X2 U9690 ( .A(n10928), .B(n10927), .Y(n6895) );
  NAND2X1 U9691 ( .A(n10533), .B(n10672), .Y(n10534) );
  NAND2X1 U9692 ( .A(n11089), .B(n11088), .Y(n11090) );
  NAND2BX1 U9693 ( .AN(n9793), .B(n9763), .Y(n6402) );
  NAND2X1 U9694 ( .A(n11232), .B(n11381), .Y(n11233) );
  NAND2X1 U9695 ( .A(n10631), .B(n10630), .Y(n10632) );
  NOR2BX1 U9696 ( .AN(n11088), .B(n6222), .Y(n6221) );
  NAND2X1 U9697 ( .A(n9866), .B(n9865), .Y(n10126) );
  NAND2X1 U9698 ( .A(n28963), .B(n5927), .Y(n27155) );
  NAND2X1 U9699 ( .A(n10179), .B(n10181), .Y(n10184) );
  NAND2X1 U9700 ( .A(n11193), .B(n11192), .Y(n11194) );
  AND2X2 U9701 ( .A(n9950), .B(n9949), .Y(n10215) );
  NAND2X1 U9702 ( .A(n10652), .B(n10651), .Y(n10653) );
  CLKINVX8 U9703 ( .A(n5808), .Y(n5834) );
  NAND2X1 U9704 ( .A(n9835), .B(n9834), .Y(n10168) );
  NAND2X1 U9705 ( .A(n10728), .B(n10727), .Y(n10729) );
  NAND2X1 U9706 ( .A(n9954), .B(n9953), .Y(n10244) );
  OR2XL U9707 ( .A(n20438), .B(U0_pipe6[26]), .Y(n6727) );
  NAND2X1 U9708 ( .A(n10487), .B(n10486), .Y(n10488) );
  NAND2X1 U9709 ( .A(n11152), .B(n11151), .Y(n11153) );
  NAND2X1 U9710 ( .A(n10818), .B(n8251), .Y(n6422) );
  NAND2X1 U9711 ( .A(n9843), .B(n9842), .Y(n10188) );
  INVX1 U9712 ( .A(n5812), .Y(n5835) );
  NAND2XL U9713 ( .A(n13746), .B(n13752), .Y(n13754) );
  NAND2X1 U9714 ( .A(n11341), .B(n11340), .Y(n11342) );
  NAND2X1 U9715 ( .A(n11143), .B(n11142), .Y(n11144) );
  NAND2X1 U9716 ( .A(BOPA[7]), .B(n11430), .Y(n9611) );
  NAND2X1 U9717 ( .A(n10367), .B(n10366), .Y(n10368) );
  NAND2X1 U9718 ( .A(n11046), .B(n11209), .Y(n11047) );
  NAND2X1 U9719 ( .A(n10942), .B(n10941), .Y(n10943) );
  NAND2X1 U9720 ( .A(n10822), .B(n10821), .Y(n10823) );
  NAND2X1 U9721 ( .A(n11336), .B(n8336), .Y(n11322) );
  NAND2X1 U9722 ( .A(n10876), .B(n11022), .Y(n10877) );
  NAND2X1 U9723 ( .A(n10902), .B(n10901), .Y(n10903) );
  AOI22X1 U9724 ( .A0(n7305), .A1(n14996), .B0(C_sel_reg[8]), .B1(n14995), .Y(
        n14997) );
  NAND2X1 U9725 ( .A(n9805), .B(n9804), .Y(n10081) );
  INVXL U9726 ( .A(n25330), .Y(n5971) );
  INVXL U9727 ( .A(n25330), .Y(n5940) );
  AOI21XL U9728 ( .A0(n13739), .A1(n8143), .B0(n13738), .Y(n13740) );
  CLKBUFX8 U9729 ( .A(n25330), .Y(n6888) );
  NAND2X1 U9730 ( .A(BOPA[10]), .B(n11430), .Y(n9618) );
  AND2XL U9731 ( .A(n12689), .B(U1_U1_y0[13]), .Y(n6998) );
  INVX8 U9732 ( .A(n27976), .Y(n27814) );
  INVX1 U9733 ( .A(n11146), .Y(n11160) );
  INVX1 U9734 ( .A(n9748), .Y(n9750) );
  INVX1 U9735 ( .A(n11128), .Y(n11143) );
  NOR2X1 U9736 ( .A(n11288), .B(n11284), .Y(n11276) );
  AOI21XL U9737 ( .A0(n13743), .A1(n13749), .B0(n13748), .Y(n13755) );
  CLKBUFX8 U9738 ( .A(n25330), .Y(n21972) );
  INVX8 U9739 ( .A(n27213), .Y(n5927) );
  INVX1 U9740 ( .A(n9859), .Y(n9861) );
  NAND2X1 U9741 ( .A(n11976), .B(cnt[10]), .Y(n11632) );
  INVX1 U9742 ( .A(n9793), .Y(n9795) );
  OAI21X1 U9743 ( .A0(n11100), .A1(n11105), .B0(n11101), .Y(n11093) );
  NOR2X1 U9744 ( .A(n10866), .B(n10868), .Y(n10896) );
  NOR2X1 U9745 ( .A(n10930), .B(n10926), .Y(n10920) );
  INVX1 U9746 ( .A(n11310), .Y(n11324) );
  INVX1 U9747 ( .A(n9938), .Y(n9940) );
  INVX1 U9748 ( .A(n9982), .Y(n9984) );
  NOR2XL U9749 ( .A(n14170), .B(U0_U0_y0[13]), .Y(n14160) );
  INVX1 U9750 ( .A(n10223), .Y(n10226) );
  INVX1 U9751 ( .A(n10435), .Y(n10449) );
  INVX1 U9752 ( .A(n9907), .Y(n9909) );
  INVX1 U9753 ( .A(n10315), .Y(n10318) );
  INVX1 U9754 ( .A(n10515), .Y(n10348) );
  CLKBUFX8 U9755 ( .A(n25330), .Y(n20438) );
  INVX4 U9756 ( .A(n20240), .Y(n5837) );
  NOR2X1 U9757 ( .A(n10272), .B(n10301), .Y(n10274) );
  INVXL U9758 ( .A(U0_U2_y0[13]), .Y(n6364) );
  NOR2X1 U9759 ( .A(n10755), .B(n10756), .Y(n10746) );
  CLKBUFX8 U9760 ( .A(n25330), .Y(n22620) );
  INVX1 U9761 ( .A(n10954), .Y(n10968) );
  INVX1 U9762 ( .A(n10846), .Y(n10706) );
  CLKBUFX8 U9763 ( .A(n25330), .Y(n19215) );
  INVX1 U9764 ( .A(n10147), .Y(n10148) );
  INVX1 U9765 ( .A(n9812), .Y(n8353) );
  INVX1 U9766 ( .A(n9826), .Y(n9828) );
  INVX1 U9767 ( .A(n10090), .Y(n10093) );
  INVX1 U9768 ( .A(n9986), .Y(n9988) );
  CLKBUFX8 U9769 ( .A(n25330), .Y(n22853) );
  NAND2X1 U9770 ( .A(n11418), .B(BOPA[2]), .Y(n8304) );
  CLKBUFX8 U9771 ( .A(n25330), .Y(n19405) );
  NAND2X1 U9772 ( .A(n11418), .B(BOPA[4]), .Y(n8307) );
  INVX1 U9773 ( .A(n9818), .Y(n9866) );
  INVX1 U9774 ( .A(n18987), .Y(n5929) );
  INVX2 U9775 ( .A(n25330), .Y(n17249) );
  INVX1 U9776 ( .A(B1_q[8]), .Y(n16323) );
  NAND2X1 U9777 ( .A(W1[15]), .B(n7976), .Y(n10255) );
  NOR2X1 U9778 ( .A(n8159), .B(BOPD[48]), .Y(n10726) );
  NOR2X1 U9779 ( .A(n8162), .B(BOPD[47]), .Y(n10693) );
  NOR2X1 U9780 ( .A(n8152), .B(BOPD[50]), .Y(n10846) );
  NAND2X1 U9781 ( .A(n8152), .B(BOPD[50]), .Y(n10849) );
  INVX1 U9782 ( .A(B1_q[49]), .Y(n16369) );
  NOR2X1 U9783 ( .A(n6950), .B(AOPD[44]), .Y(n10911) );
  NOR2X2 U9784 ( .A(n8112), .B(AOPD[43]), .Y(n10926) );
  NAND2X1 U9785 ( .A(n8112), .B(AOPD[43]), .Y(n10927) );
  INVX1 U9786 ( .A(B1_q[48]), .Y(n16373) );
  INVX1 U9787 ( .A(B1_q[47]), .Y(n16378) );
  NOR2X1 U9788 ( .A(n8088), .B(AOPD[50]), .Y(n11020) );
  NOR2X1 U9789 ( .A(AOPD[25]), .B(n8056), .Y(n11024) );
  NAND2X1 U9790 ( .A(n8088), .B(AOPD[50]), .Y(n11023) );
  INVX1 U9791 ( .A(B1_q[46]), .Y(n16382) );
  INVX2 U9792 ( .A(n9831), .Y(n5839) );
  NAND2X1 U9793 ( .A(n8065), .B(AOPD[33]), .Y(n8317) );
  INVX1 U9794 ( .A(B0_q[51]), .Y(n16361) );
  INVX1 U9795 ( .A(B1_q[50]), .Y(n16365) );
  INVX8 U9796 ( .A(n28697), .Y(n24380) );
  NAND2X1 U9797 ( .A(n8066), .B(AOPB[33]), .Y(n10482) );
  NAND2X1 U9798 ( .A(n8021), .B(W3[19]), .Y(n10012) );
  NOR2X1 U9799 ( .A(n8110), .B(AOPB[44]), .Y(n10387) );
  NOR2X1 U9800 ( .A(n8092), .B(AOPB[49]), .Y(n10365) );
  NOR2X1 U9801 ( .A(n8089), .B(AOPB[50]), .Y(n10512) );
  NOR2X1 U9802 ( .A(AOPB[25]), .B(n8073), .Y(n10516) );
  NAND2X1 U9803 ( .A(n8089), .B(AOPB[50]), .Y(n10515) );
  NAND2X1 U9804 ( .A(W2[13]), .B(W2[29]), .Y(n9882) );
  AND2XL U9805 ( .A(U1_U0_y2[12]), .B(U1_U0_y0[12]), .Y(n8398) );
  OR2XL U9806 ( .A(U1_U0_y2[8]), .B(U1_U0_y0[8]), .Y(n8386) );
  NAND2X1 U9807 ( .A(n8175), .B(BOPB[43]), .Y(n10588) );
  NOR2X1 U9808 ( .A(n8163), .B(BOPB[46]), .Y(n10553) );
  NOR2X1 U9809 ( .A(n8160), .B(BOPB[47]), .Y(n10559) );
  NOR2X1 U9810 ( .A(BOPB[25]), .B(n8129), .Y(n10674) );
  INVXL U9811 ( .A(U1_A_r_d0[20]), .Y(n6189) );
  INVX1 U9812 ( .A(B1_q[19]), .Y(n16494) );
  NAND2X1 U9813 ( .A(W3[9]), .B(W3[25]), .Y(n9787) );
  INVX1 U9814 ( .A(B1_q[12]), .Y(n16523) );
  INVX1 U9815 ( .A(B1_q[13]), .Y(n16519) );
  INVX1 U9816 ( .A(B1_q[14]), .Y(n16303) );
  NOR2X1 U9817 ( .A(W3[20]), .B(W3[4]), .Y(n9778) );
  INVX1 U9818 ( .A(B1_q[17]), .Y(n16504) );
  INVX1 U9819 ( .A(B1_q[23]), .Y(n16477) );
  BUFX8 U9820 ( .A(U1_valid[0]), .Y(n25330) );
  INVX1 U9821 ( .A(B1_q[24]), .Y(n16473) );
  OR2XL U9822 ( .A(U1_U0_y1[8]), .B(U1_U0_y0[8]), .Y(n9271) );
  INVX1 U9823 ( .A(B1_q[21]), .Y(n16485) );
  INVX1 U9824 ( .A(B5_q[43]), .Y(n15807) );
  INVX1 U9825 ( .A(B5_q[25]), .Y(n15879) );
  INVX1 U9826 ( .A(B5_q[48]), .Y(n15787) );
  INVX1 U9827 ( .A(B5_q[36]), .Y(n15835) );
  INVX1 U9828 ( .A(B5_q[49]), .Y(n15783) );
  INVX1 U9829 ( .A(B7_q[45]), .Y(n15799) );
  INVX1 U9830 ( .A(B5_q[32]), .Y(n15650) );
  INVX1 U9831 ( .A(B5_q[26]), .Y(n15875) );
  INVX1 U9832 ( .A(B5_q[1]), .Y(n15980) );
  INVX1 U9833 ( .A(B5_q[18]), .Y(n15701) );
  INVX1 U9834 ( .A(B1_q[10]), .Y(n16531) );
  INVX1 U9835 ( .A(B2_q[18]), .Y(n16287) );
  INVX4 U9836 ( .A(n16136), .Y(n5841) );
  INVX1 U9837 ( .A(B1_q[33]), .Y(n16435) );
  NAND2X1 U9838 ( .A(n8087), .B(AOPC[50]), .Y(n11382) );
  NOR2X1 U9839 ( .A(AOPC[25]), .B(n8055), .Y(n11383) );
  NOR2X1 U9840 ( .A(n8087), .B(AOPC[50]), .Y(n11379) );
  INVX1 U9841 ( .A(B0_q[29]), .Y(n16451) );
  INVX1 U9842 ( .A(B3_q[41]), .Y(n16205) );
  INVX1 U9843 ( .A(B1_q[44]), .Y(n16390) );
  INVX1 U9844 ( .A(B0_q[37]), .Y(n16419) );
  NAND2X1 U9845 ( .A(n8151), .B(BOPC[50]), .Y(n11210) );
  INVX1 U9846 ( .A(B0_q[38]), .Y(n16414) );
  NOR2X1 U9847 ( .A(n8161), .B(BOPC[47]), .Y(n11075) );
  NOR2X1 U9848 ( .A(n8158), .B(BOPC[48]), .Y(n11064) );
  INVX1 U9849 ( .A(B1_q[39]), .Y(n16410) );
  INVX1 U9850 ( .A(B1_q[3]), .Y(n16342) );
  OR2X2 U9851 ( .A(W3[14]), .B(W3[30]), .Y(n9740) );
  OR2XL U9852 ( .A(U1_U2_y2[10]), .B(U1_U2_y0[10]), .Y(n13763) );
  OR2X2 U9853 ( .A(U1_U2_y2[9]), .B(U1_U2_y0[9]), .Y(n13760) );
  OR2XL U9854 ( .A(U1_U2_y2[8]), .B(U1_U2_y0[8]), .Y(n13761) );
  NOR2X1 U9855 ( .A(W3[13]), .B(W3[29]), .Y(n9742) );
  NAND2X1 U9856 ( .A(W3[13]), .B(W3[29]), .Y(n9743) );
  INVX1 U9857 ( .A(B3_q[28]), .Y(n16251) );
  OR2X2 U9858 ( .A(BOPA[49]), .B(BOPA[48]), .Y(n6407) );
  NAND2X1 U9859 ( .A(W3[12]), .B(W3[28]), .Y(n9804) );
  NAND2X1 U9860 ( .A(n8037), .B(W3[22]), .Y(n10044) );
  AOI22X1 U9861 ( .A0(cnt[7]), .A1(n28673), .B0(cnt[5]), .B1(n28703), .Y(
        n11610) );
  OR2XL U9862 ( .A(U0_U1_y2[8]), .B(U0_U1_y0[8]), .Y(n12434) );
  OR2XL U9863 ( .A(U0_U0_y2[8]), .B(U0_U0_y0[8]), .Y(n14176) );
  OR2XL U9864 ( .A(U0_U0_y2[12]), .B(U0_U0_y0[12]), .Y(n14161) );
  OR2XL U9865 ( .A(U0_U2_y1[8]), .B(U0_U2_y0[8]), .Y(n8720) );
  INVXL U9866 ( .A(U1_A_r_d0[12]), .Y(n6182) );
  INVX1 U9867 ( .A(n6832), .Y(n22297) );
  NAND3XL U9868 ( .A(n7030), .B(n7483), .C(n7481), .Y(n4979) );
  NAND2XL U9869 ( .A(n6529), .B(n6525), .Y(n4405) );
  OAI21XL U9870 ( .A0(U1_pipe7[23]), .A1(n5812), .B0(n6077), .Y(n4976) );
  INVXL U9871 ( .A(n19388), .Y(n19389) );
  INVX1 U9872 ( .A(n14582), .Y(n14583) );
  NAND3BX1 U9873 ( .AN(n6096), .B(n7488), .C(n6095), .Y(n4836) );
  MXI2XL U9874 ( .A(n6019), .B(U1_pipe13[22]), .S0(n5811), .Y(n4745) );
  XOR2X1 U9875 ( .A(n7813), .B(n6099), .Y(n20027) );
  MXI2X1 U9876 ( .A(n6081), .B(U1_pipe13[25]), .S0(n5811), .Y(n4748) );
  XOR2X1 U9877 ( .A(n6020), .B(n20049), .Y(n6019) );
  XOR2X1 U9878 ( .A(n13995), .B(n6045), .Y(n7511) );
  OAI21XL U9879 ( .A0(n6341), .A1(n8053), .B0(n9238), .Y(n4406) );
  OAI21XL U9880 ( .A0(n19387), .A1(n19386), .B0(n19385), .Y(n19388) );
  NAND2X1 U9881 ( .A(n6126), .B(n6128), .Y(n6099) );
  INVX1 U9882 ( .A(n19569), .Y(n19570) );
  AOI2BB1X2 U9883 ( .A0N(n6045), .A1N(n17050), .B0(n6004), .Y(n6003) );
  MXI2XL U9884 ( .A(n6599), .B(U1_pipe6[23]), .S0(n6598), .Y(n4948) );
  MXI2XL U9885 ( .A(n7661), .B(U1_pipe10[25]), .S0(n8053), .Y(n4863) );
  NAND3BX1 U9886 ( .AN(n6634), .B(n6577), .C(n6573), .Y(n6572) );
  NAND2XL U9887 ( .A(n7651), .B(n7631), .Y(n7625) );
  XOR2X1 U9888 ( .A(n25658), .B(n6456), .Y(n25659) );
  INVX1 U9889 ( .A(n7866), .Y(n20053) );
  INVXL U9890 ( .A(n22457), .Y(n22458) );
  MXI2XL U9891 ( .A(n6199), .B(U0_pipe7[24]), .S0(n5838), .Y(n4438) );
  NOR2X1 U9892 ( .A(n6115), .B(n6112), .Y(n19232) );
  MXI2XL U9893 ( .A(n7163), .B(U1_pipe6[27]), .S0(n8053), .Y(n4952) );
  MXI2XL U9894 ( .A(n7783), .B(U1_pipe11[27]), .S0(n8053), .Y(n4893) );
  NOR2X1 U9895 ( .A(n7475), .B(n6135), .Y(n20334) );
  XOR2X1 U9896 ( .A(n25653), .B(n7006), .Y(n12285) );
  XNOR2X1 U9897 ( .A(n17473), .B(n17472), .Y(n17474) );
  XOR2X1 U9898 ( .A(n6201), .B(n6200), .Y(n6199) );
  NOR2XL U9899 ( .A(n7486), .B(n7938), .Y(n7484) );
  MXI2XL U9900 ( .A(n6362), .B(U0_pipe1[16]), .S0(n6361), .Y(n4268) );
  XOR2X1 U9901 ( .A(n6600), .B(n16947), .Y(n6599) );
  XOR2X1 U9902 ( .A(n6388), .B(n25329), .Y(n25331) );
  NAND2XL U9903 ( .A(n14108), .B(n7213), .Y(n7212) );
  INVX1 U9904 ( .A(n7208), .Y(n6798) );
  NAND3BX2 U9905 ( .AN(n12406), .B(n25289), .C(n12403), .Y(n6302) );
  MXI2XL U9906 ( .A(n6672), .B(U1_pipe6[22]), .S0(n6671), .Y(n4947) );
  AOI21X2 U9907 ( .A0(n25663), .A1(n6990), .B0(n7557), .Y(n25661) );
  CLKINVX3 U9908 ( .A(n7157), .Y(n20350) );
  NAND2XL U9909 ( .A(n7551), .B(n17305), .Y(n17310) );
  NAND2XL U9910 ( .A(n6585), .B(n16961), .Y(n16963) );
  NAND2XL U9911 ( .A(n6677), .B(n19804), .Y(n19809) );
  XOR2X1 U9912 ( .A(n7348), .B(n23007), .Y(n23008) );
  XOR2X1 U9913 ( .A(n6775), .B(n24722), .Y(n24723) );
  XOR2X1 U9914 ( .A(n6363), .B(n25032), .Y(n6362) );
  NAND2X1 U9915 ( .A(n7470), .B(n16793), .Y(n6080) );
  NAND2XL U9916 ( .A(n7939), .B(n25330), .Y(n7486) );
  INVXL U9917 ( .A(n22592), .Y(n6797) );
  NAND2BXL U9918 ( .AN(n7939), .B(n25330), .Y(n7479) );
  NAND3X1 U9919 ( .A(n6517), .B(n8688), .C(n6516), .Y(n7166) );
  XOR2X1 U9920 ( .A(n6842), .B(n22324), .Y(n22325) );
  NOR2XL U9921 ( .A(n7938), .B(n17249), .Y(n7482) );
  INVXL U9922 ( .A(n17081), .Y(n17076) );
  INVX1 U9923 ( .A(n24988), .Y(n5842) );
  NOR2XL U9924 ( .A(n14107), .B(n7504), .Y(n7503) );
  NAND3X1 U9925 ( .A(n16633), .B(n6518), .C(n8689), .Y(n6517) );
  NAND2X1 U9926 ( .A(n17304), .B(n7860), .Y(n6150) );
  INVXL U9927 ( .A(n16633), .Y(n16652) );
  INVX2 U9928 ( .A(n17602), .Y(n17625) );
  NAND2XL U9929 ( .A(n7444), .B(n20355), .Y(n20358) );
  INVXL U9930 ( .A(n7938), .Y(n7480) );
  AND2X2 U9931 ( .A(n6298), .B(n12341), .Y(n6530) );
  NAND2BX1 U9932 ( .AN(n25651), .B(n6474), .Y(n6473) );
  MXI2XL U9933 ( .A(n6503), .B(U0_pipe4[20]), .S0(n5838), .Y(n4327) );
  INVXL U9934 ( .A(n22979), .Y(n22980) );
  INVXL U9935 ( .A(n17456), .Y(n7617) );
  NAND2BXL U9936 ( .AN(n14128), .B(n7210), .Y(n7209) );
  NAND2XL U9937 ( .A(n25654), .B(n24696), .Y(n6317) );
  NAND2XL U9938 ( .A(n9603), .B(n7312), .Y(n7311) );
  INVXL U9939 ( .A(n17347), .Y(n17339) );
  ADDFHX2 U9940 ( .A(n25123), .B(n29009), .CI(n21810), .CO(n21808), .S(n21811)
         );
  NAND2BX1 U9941 ( .AN(n14894), .B(n7746), .Y(n7745) );
  OAI2BB1X2 U9942 ( .A0N(n17323), .A1N(n17370), .B0(n7782), .Y(n17347) );
  OAI21X1 U9943 ( .A0(n16969), .A1(n16959), .B0(n16960), .Y(n6586) );
  AND2X2 U9944 ( .A(n12342), .B(n12341), .Y(n24698) );
  INVXL U9945 ( .A(n19575), .Y(n7810) );
  NAND2XL U9946 ( .A(n7643), .B(n7646), .Y(n7630) );
  NOR2BX2 U9947 ( .AN(n14567), .B(n6538), .Y(n6537) );
  NAND2X1 U9948 ( .A(n22594), .B(n7735), .Y(n6238) );
  NAND2X1 U9949 ( .A(n14006), .B(n5965), .Y(n5961) );
  INVXL U9950 ( .A(n17457), .Y(n7618) );
  NAND3X1 U9951 ( .A(n5966), .B(n5965), .C(n14007), .Y(n5964) );
  OR2XL U9952 ( .A(n14976), .B(n7814), .Y(n7047) );
  INVX1 U9953 ( .A(n7735), .Y(n22595) );
  AND2X2 U9954 ( .A(n22594), .B(n22593), .Y(n22974) );
  NAND2BXL U9955 ( .AN(n25292), .B(n25652), .Y(n6475) );
  OAI21X2 U9956 ( .A0(n7415), .A1(n7414), .B0(n6427), .Y(n6426) );
  INVXL U9957 ( .A(n9604), .Y(n7315) );
  INVXL U9958 ( .A(n17605), .Y(n17606) );
  AOI21X1 U9959 ( .A0(n13623), .A1(n17301), .B0(n7494), .Y(n6149) );
  NAND2X2 U9960 ( .A(n25321), .B(n12397), .Y(n6379) );
  XOR2X1 U9961 ( .A(n17636), .B(n17635), .Y(n17637) );
  INVX1 U9962 ( .A(n20194), .Y(n20206) );
  XNOR2XL U9963 ( .A(n25046), .B(n25045), .Y(n25047) );
  NAND3X1 U9964 ( .A(n16809), .B(n7455), .C(n16855), .Y(n6167) );
  XOR2X1 U9965 ( .A(n6005), .B(n19260), .Y(n19261) );
  AND2X1 U9966 ( .A(n20023), .B(n20029), .Y(n20024) );
  NAND3X2 U9967 ( .A(n6039), .B(n6036), .C(n6035), .Y(n17602) );
  AND2X2 U9968 ( .A(n20019), .B(n20038), .Y(n6093) );
  INVXL U9969 ( .A(n17465), .Y(n17466) );
  INVXL U9970 ( .A(n19566), .Y(n7877) );
  XOR2X1 U9971 ( .A(n6857), .B(n14105), .Y(n14106) );
  NAND2X1 U9972 ( .A(n20037), .B(n20019), .Y(n20031) );
  INVXL U9973 ( .A(n20341), .Y(n7864) );
  NAND2BXL U9974 ( .AN(n19835), .B(n7530), .Y(n7529) );
  INVXL U9975 ( .A(n17297), .Y(n7504) );
  NOR2X1 U9976 ( .A(n7437), .B(n5957), .Y(n20316) );
  NAND2BXL U9977 ( .AN(n12338), .B(n12337), .Y(n7715) );
  NAND2BXL U9978 ( .AN(n17177), .B(n17175), .Y(n7750) );
  INVX1 U9979 ( .A(n22185), .Y(n22197) );
  NAND2BXL U9980 ( .AN(n14976), .B(n7861), .Y(n7784) );
  NAND2X1 U9981 ( .A(n20029), .B(n7255), .Y(n7254) );
  INVX1 U9982 ( .A(n17296), .Y(n13651) );
  AND2X2 U9983 ( .A(n7177), .B(n6231), .Y(n6232) );
  AND2X2 U9984 ( .A(n6934), .B(n21984), .Y(n22324) );
  NAND2X1 U9985 ( .A(n6240), .B(n6239), .Y(n7735) );
  NAND3X1 U9986 ( .A(n17524), .B(n9517), .C(n17478), .Y(n7626) );
  NAND2XL U9987 ( .A(n7650), .B(n7649), .Y(n7648) );
  INVX1 U9988 ( .A(n13948), .Y(n6046) );
  OAI21XL U9989 ( .A0(U1_pipe12[26]), .A1(n5810), .B0(n6620), .Y(n6619) );
  INVXL U9990 ( .A(n22972), .Y(n6815) );
  INVXL U9991 ( .A(n6626), .Y(n6623) );
  NAND2XL U9992 ( .A(n7527), .B(n6621), .Y(n6620) );
  NAND2BX2 U9993 ( .AN(n19415), .B(n6954), .Y(n13706) );
  AOI2BB1X2 U9994 ( .A0N(n14504), .A1N(n6041), .B0(n6037), .Y(n6036) );
  INVXL U9995 ( .A(n20345), .Y(n20321) );
  AND2XL U9996 ( .A(n14575), .B(n24676), .Y(n8082) );
  XNOR2XL U9997 ( .A(n20101), .B(n20100), .Y(n20102) );
  XNOR2XL U9998 ( .A(n21879), .B(n21878), .Y(n21880) );
  NOR2XL U9999 ( .A(n5816), .B(U1_A_i_d0[25]), .Y(n6609) );
  XNOR2XL U10000 ( .A(n25722), .B(n25721), .Y(n25723) );
  XOR2XL U10001 ( .A(n22212), .B(n22216), .Y(n22217) );
  NAND3X2 U10002 ( .A(n6175), .B(n21656), .C(n6174), .Y(n7417) );
  NAND2XL U10003 ( .A(n22498), .B(n5818), .Y(n7574) );
  INVXL U10004 ( .A(n17178), .Y(n17176) );
  INVX1 U10005 ( .A(n20333), .Y(n5843) );
  NAND2XL U10006 ( .A(n7671), .B(n7670), .Y(n7669) );
  NAND2X1 U10007 ( .A(n20033), .B(n20032), .Y(n20329) );
  NAND2BXL U10008 ( .AN(n7654), .B(n9547), .Y(n7650) );
  OAI2BB1XL U10009 ( .A0N(n9548), .A1N(n9547), .B0(n7654), .Y(n7649) );
  INVXL U10010 ( .A(n24897), .Y(n24892) );
  NAND2X1 U10011 ( .A(n14505), .B(n6040), .Y(n6035) );
  NAND3X1 U10012 ( .A(n17370), .B(n17323), .C(n13563), .Y(n7497) );
  NOR2BX1 U10013 ( .AN(n14972), .B(n19233), .Y(n17596) );
  INVX1 U10014 ( .A(n24873), .Y(n24885) );
  NAND2X1 U10015 ( .A(n20061), .B(n20059), .Y(n6016) );
  NOR2X1 U10016 ( .A(n17306), .B(n17307), .Y(n13624) );
  NAND2BX1 U10017 ( .AN(n25010), .B(n25008), .Y(n6366) );
  XNOR2XL U10018 ( .A(n25205), .B(n25204), .Y(n25206) );
  INVXL U10019 ( .A(n25694), .Y(n25340) );
  INVXL U10020 ( .A(n25309), .Y(n6469) );
  INVX1 U10021 ( .A(n20032), .Y(n20020) );
  INVXL U10022 ( .A(n9722), .Y(n7351) );
  NAND3X2 U10023 ( .A(n6839), .B(n6837), .C(n22928), .Y(n23049) );
  AOI21X1 U10024 ( .A0(n20325), .A1(n20324), .B0(n20323), .Y(n7478) );
  OR2X2 U10025 ( .A(n24685), .B(n24684), .Y(n24686) );
  AOI21X1 U10026 ( .A0(n20009), .A1(n20085), .B0(n20008), .Y(n6017) );
  XNOR2XL U10027 ( .A(n19150), .B(n19149), .Y(n19151) );
  NAND3BX2 U10028 ( .AN(n13525), .B(n6545), .C(n6546), .Y(n24873) );
  INVXL U10029 ( .A(n6508), .Y(n25138) );
  INVXL U10030 ( .A(n19585), .Y(n19249) );
  NAND2BX1 U10031 ( .AN(n13996), .B(n6551), .Y(n24897) );
  NAND3X2 U10032 ( .A(n5980), .B(n5979), .C(n5977), .Y(n16855) );
  NAND2BX1 U10033 ( .AN(n23052), .B(n6838), .Y(n6837) );
  AND2X2 U10034 ( .A(n14966), .B(n14961), .Y(n6086) );
  NAND2X1 U10035 ( .A(n6314), .B(n6313), .Y(n12394) );
  INVXL U10036 ( .A(n24501), .Y(n24449) );
  INVXL U10037 ( .A(n19787), .Y(n7525) );
  OR2X2 U10038 ( .A(n6047), .B(n5969), .Y(n14009) );
  INVX1 U10039 ( .A(n17064), .Y(n16804) );
  INVXL U10040 ( .A(n19788), .Y(n6650) );
  NOR2X1 U10041 ( .A(n13556), .B(n7517), .Y(n7516) );
  NOR2X1 U10042 ( .A(n13945), .B(n17083), .Y(n14007) );
  AND2X2 U10043 ( .A(n13622), .B(n17314), .Y(n7495) );
  NAND2X1 U10044 ( .A(n14546), .B(n22024), .Y(n7152) );
  INVXL U10045 ( .A(n19825), .Y(n7530) );
  INVXL U10046 ( .A(n9536), .Y(n7670) );
  NOR2X2 U10047 ( .A(n6073), .B(n17643), .Y(n14500) );
  NAND2BX1 U10048 ( .AN(n19423), .B(n19118), .Y(n19410) );
  XNOR2XL U10049 ( .A(n19299), .B(n19298), .Y(n19300) );
  AND2XL U10050 ( .A(n5817), .B(n14960), .Y(n7956) );
  NAND2X2 U10051 ( .A(n6190), .B(n6189), .Y(n6954) );
  INVXL U10052 ( .A(n17471), .Y(n17472) );
  NAND2X1 U10053 ( .A(n16826), .B(n16830), .Y(n14008) );
  INVXL U10054 ( .A(n17194), .Y(n9602) );
  NAND2BXL U10055 ( .AN(n18904), .B(n7376), .Y(n7380) );
  INVXL U10056 ( .A(n14564), .Y(n13131) );
  NAND2X1 U10057 ( .A(n14966), .B(n19243), .Y(n17308) );
  NAND2X1 U10058 ( .A(n20085), .B(n20090), .Y(n20010) );
  NOR2X1 U10059 ( .A(n19556), .B(n19596), .Y(n6102) );
  INVXL U10060 ( .A(n16628), .Y(n6576) );
  INVX1 U10061 ( .A(n22960), .Y(n6240) );
  INVXL U10062 ( .A(n7696), .Y(n9703) );
  CLKINVX3 U10063 ( .A(n14961), .Y(n5845) );
  INVX1 U10064 ( .A(n13717), .Y(n9720) );
  OR2X2 U10065 ( .A(n22958), .B(n24680), .Y(n14124) );
  AOI21X1 U10066 ( .A0(n13038), .A1(n13009), .B0(n8145), .Y(n6072) );
  INVXL U10067 ( .A(n17330), .Y(n7502) );
  NOR2X1 U10068 ( .A(n8614), .B(n16959), .Y(n8616) );
  INVXL U10069 ( .A(n16661), .Y(n7532) );
  INVXL U10070 ( .A(n24725), .Y(n6776) );
  OR2X2 U10071 ( .A(n19790), .B(n29007), .Y(n7526) );
  NAND2X1 U10072 ( .A(n20373), .B(n7005), .Y(n14887) );
  NAND3X2 U10073 ( .A(n6185), .B(n6183), .C(n13689), .Y(n7685) );
  INVXL U10074 ( .A(n25343), .Y(n25692) );
  NAND2XL U10075 ( .A(n13713), .B(U1_A_i_d0[23]), .Y(n17184) );
  NAND2X1 U10076 ( .A(n13889), .B(n17107), .Y(n5960) );
  INVXL U10077 ( .A(n19423), .Y(n19123) );
  NAND2BX2 U10078 ( .AN(n8560), .B(n7199), .Y(n16993) );
  INVXL U10079 ( .A(n19415), .Y(n19112) );
  NAND2X1 U10080 ( .A(n13009), .B(n13015), .Y(n6073) );
  INVXL U10081 ( .A(n16830), .Y(n17075) );
  OR2X2 U10082 ( .A(n14560), .B(n22933), .Y(n14552) );
  AND2X2 U10083 ( .A(n14560), .B(n22933), .Y(n14561) );
  OR2X2 U10084 ( .A(n19786), .B(U1_A_i_d0[25]), .Y(n8689) );
  AND2X2 U10085 ( .A(n6123), .B(n19243), .Y(n5994) );
  INVX1 U10086 ( .A(n16857), .Y(n16887) );
  AOI21X1 U10087 ( .A0(n19803), .A1(n19781), .B0(n19780), .Y(n19795) );
  INVXL U10088 ( .A(n22322), .Y(n13133) );
  NAND2X1 U10089 ( .A(n16857), .B(n5981), .Y(n5980) );
  NOR2X1 U10090 ( .A(n13713), .B(U1_A_r_d0[23]), .Y(n19085) );
  AOI21X1 U10091 ( .A0(n20377), .A1(n20379), .B0(n14883), .Y(n20364) );
  INVXL U10092 ( .A(n7467), .Y(n7466) );
  INVX1 U10093 ( .A(n6477), .Y(n25716) );
  INVXL U10094 ( .A(n14968), .Y(n14510) );
  INVXL U10095 ( .A(n19605), .Y(n19600) );
  INVX1 U10096 ( .A(n6743), .Y(n22353) );
  INVX2 U10097 ( .A(n22968), .Y(n5847) );
  NAND2X1 U10098 ( .A(n17639), .B(n13070), .Y(n14499) );
  OAI21X1 U10099 ( .A0(n16889), .A1(n14925), .B0(n5982), .Y(n16857) );
  AOI21XL U10100 ( .A0(n25377), .A1(n25375), .B0(n12380), .Y(n12381) );
  INVXL U10101 ( .A(n19752), .Y(n19763) );
  INVX1 U10102 ( .A(n13709), .Y(n5848) );
  NAND2BXL U10103 ( .AN(n8684), .B(n16646), .Y(n6657) );
  NAND2X1 U10104 ( .A(n22010), .B(n7016), .Y(n14559) );
  NOR2X1 U10105 ( .A(n25132), .B(U2_A_i_d[24]), .Y(n22175) );
  NAND2X1 U10106 ( .A(n25132), .B(U2_A_i_d[24]), .Y(n22174) );
  INVXL U10107 ( .A(n17221), .Y(n17215) );
  INVX1 U10108 ( .A(n22454), .Y(n14158) );
  NAND2X1 U10109 ( .A(n25132), .B(U2_A_r_d[24]), .Y(n25522) );
  NOR2X1 U10110 ( .A(n19616), .B(n19549), .Y(n19595) );
  NAND2X1 U10111 ( .A(n25353), .B(n25358), .Y(n12393) );
  NOR2X1 U10112 ( .A(n7913), .B(n19998), .Y(n6014) );
  NAND2X1 U10113 ( .A(n6334), .B(n6333), .Y(n22024) );
  AND2X2 U10114 ( .A(n16665), .B(n16961), .Y(n16965) );
  INVXL U10115 ( .A(n7602), .Y(n24504) );
  OR2X2 U10116 ( .A(n6440), .B(n6442), .Y(n6359) );
  INVX1 U10117 ( .A(n12334), .Y(n19786) );
  INVXL U10118 ( .A(n19552), .Y(n7792) );
  NAND2X1 U10119 ( .A(n19605), .B(n6947), .Y(n19556) );
  NAND3X2 U10120 ( .A(n6553), .B(n13512), .C(n6552), .Y(n24917) );
  AOI21XL U10121 ( .A0(n7018), .A1(n17110), .B0(n13885), .Y(n13886) );
  INVXL U10122 ( .A(n25703), .Y(n25710) );
  INVX1 U10123 ( .A(n14550), .Y(n5852) );
  CLKINVX3 U10124 ( .A(n14852), .Y(n20048) );
  NAND2X1 U10125 ( .A(n22453), .B(U2_A_r_d[24]), .Y(n24425) );
  NAND2BX1 U10126 ( .AN(n13395), .B(n7586), .Y(n7602) );
  INVXL U10127 ( .A(n19604), .Y(n7879) );
  CLKINVX3 U10128 ( .A(n14960), .Y(n5853) );
  CLKINVX3 U10129 ( .A(n22446), .Y(n5854) );
  NAND3X2 U10130 ( .A(n5938), .B(n5935), .C(n13952), .Y(n7836) );
  OR2X2 U10131 ( .A(n14529), .B(n22058), .Y(n6334) );
  NAND2X1 U10132 ( .A(n7672), .B(n9518), .Y(n9525) );
  INVXL U10133 ( .A(n24445), .Y(n24880) );
  INVXL U10134 ( .A(n17345), .Y(n17338) );
  NAND2X1 U10135 ( .A(n7409), .B(n5820), .Y(n25040) );
  OR2X2 U10136 ( .A(n9700), .B(U1_A_r_d0[17]), .Y(n9689) );
  INVXL U10137 ( .A(n17639), .Y(n7215) );
  NOR2X1 U10138 ( .A(n6188), .B(n13684), .Y(n19451) );
  INVX1 U10139 ( .A(n13690), .Y(n6186) );
  INVXL U10140 ( .A(n25358), .Y(n25351) );
  NAND2X1 U10141 ( .A(n6995), .B(n24461), .Y(n13524) );
  OR2X2 U10142 ( .A(n22926), .B(n24633), .Y(n23056) );
  NAND4X2 U10143 ( .A(n6453), .B(n6451), .C(n6450), .D(n12254), .Y(n12264) );
  INVXL U10144 ( .A(n23009), .Y(n23004) );
  NOR2XL U10145 ( .A(n13690), .B(n19452), .Y(n6184) );
  NOR2X1 U10146 ( .A(n17668), .B(n12973), .Y(n6031) );
  INVXL U10147 ( .A(n16848), .Y(n14952) );
  NAND2X1 U10148 ( .A(n19287), .B(n14830), .Y(n14832) );
  INVX1 U10149 ( .A(n12600), .Y(n22638) );
  INVXL U10150 ( .A(n16647), .Y(n6674) );
  AND2XL U10151 ( .A(n9694), .B(U1_A_i_d0[16]), .Y(n9505) );
  AND2X2 U10152 ( .A(n6938), .B(n20094), .Y(n6018) );
  CLKINVX3 U10153 ( .A(n13037), .Y(n14954) );
  NAND3X2 U10154 ( .A(n6702), .B(n13961), .C(n5992), .Y(n13970) );
  AND2XL U10155 ( .A(n7543), .B(U1_A_r_d0[18]), .Y(n7039) );
  AND2XL U10156 ( .A(n8675), .B(U1_A_r_d0[20]), .Y(n19768) );
  INVXL U10157 ( .A(n19259), .Y(n7916) );
  NAND2X1 U10158 ( .A(n17099), .B(n17104), .Y(n17083) );
  NAND2X1 U10159 ( .A(n22453), .B(U2_A_i_d[24]), .Y(n22469) );
  AND2XL U10160 ( .A(n21784), .B(U2_A_i_d[20]), .Y(n21785) );
  CLKINVX3 U10161 ( .A(n14959), .Y(n5856) );
  CLKINVX2 U10162 ( .A(n14851), .Y(n20051) );
  AOI21X2 U10163 ( .A0(n5991), .A1(n13950), .B0(n6480), .Y(n5939) );
  NAND2X1 U10164 ( .A(n6480), .B(n5822), .Y(n5938) );
  AND2X2 U10165 ( .A(n16890), .B(n14903), .Y(n5974) );
  AND2X2 U10166 ( .A(n19776), .B(U1_A_i_d0[21]), .Y(n16646) );
  OR2X2 U10167 ( .A(n24647), .B(n14548), .Y(n12204) );
  INVX1 U10168 ( .A(n22959), .Y(n5858) );
  INVXL U10169 ( .A(n16853), .Y(n16847) );
  AND2XL U10170 ( .A(n21784), .B(U2_A_r_d[20]), .Y(n14454) );
  AND2X2 U10171 ( .A(n6951), .B(n22156), .Y(n22206) );
  INVXL U10172 ( .A(n22932), .Y(n7229) );
  OR2X2 U10173 ( .A(n12388), .B(n24647), .Y(n12385) );
  INVXL U10174 ( .A(n7603), .Y(n7601) );
  CLKINVX3 U10175 ( .A(n14555), .Y(n13125) );
  INVX4 U10176 ( .A(n12224), .Y(n12247) );
  INVX1 U10177 ( .A(n23051), .Y(n23081) );
  NAND2X1 U10178 ( .A(n8523), .B(n6579), .Y(n6580) );
  INVXL U10179 ( .A(n24890), .Y(n13520) );
  NAND2X1 U10180 ( .A(n24645), .B(n24652), .Y(n25033) );
  NOR2XL U10181 ( .A(n23066), .B(n23068), .Y(n6802) );
  OR2X2 U10182 ( .A(n13513), .B(n24920), .Y(n6552) );
  INVX1 U10183 ( .A(n24434), .Y(n5860) );
  INVXL U10184 ( .A(n16674), .Y(n16968) );
  NAND2X2 U10185 ( .A(n6452), .B(n7243), .Y(n6450) );
  INVXL U10186 ( .A(n17117), .Y(n13883) );
  INVXL U10187 ( .A(n13912), .Y(n17099) );
  AND2XL U10188 ( .A(n19767), .B(U1_A_i_d0[19]), .Y(n16659) );
  AND2XL U10189 ( .A(n12379), .B(n22917), .Y(n7965) );
  AND2X2 U10190 ( .A(n13686), .B(n13685), .Y(n6188) );
  AND2XL U10191 ( .A(n19758), .B(U1_A_i_d0[14]), .Y(n8669) );
  INVX1 U10192 ( .A(n19751), .Y(n19761) );
  INVXL U10193 ( .A(n22010), .Y(n22004) );
  OR2X2 U10194 ( .A(n24647), .B(n24649), .Y(n9136) );
  OR2X2 U10195 ( .A(n12388), .B(n22936), .Y(n14549) );
  INVXL U10196 ( .A(n20117), .Y(n19982) );
  CLKINVX3 U10197 ( .A(n14963), .Y(n5861) );
  NOR2BX1 U10198 ( .AN(n13114), .B(n24615), .Y(n25389) );
  OR2X2 U10199 ( .A(n22938), .B(n24649), .Y(n22937) );
  NAND2XL U10200 ( .A(n24631), .B(n24620), .Y(n24786) );
  OR2X2 U10201 ( .A(n20002), .B(n20001), .Y(n19995) );
  INVXL U10202 ( .A(n24619), .Y(n24634) );
  INVXL U10203 ( .A(n21575), .Y(n6173) );
  NAND2X2 U10204 ( .A(n5990), .B(n7200), .Y(n5993) );
  OR2X2 U10205 ( .A(n22449), .B(U2_A_i_d[22]), .Y(n22447) );
  NAND2X1 U10206 ( .A(n6309), .B(n9091), .Y(n6533) );
  MXI2X2 U10207 ( .A(n7776), .B(n7228), .S0(n9077), .Y(n7227) );
  OR2X2 U10208 ( .A(n22449), .B(U2_A_r_d[22]), .Y(n13527) );
  NOR2XL U10209 ( .A(n6228), .B(n6227), .Y(n13450) );
  NAND2X1 U10210 ( .A(n9681), .B(n6182), .Y(n19158) );
  OR2X2 U10211 ( .A(n19754), .B(U1_A_i_d0[14]), .Y(n8580) );
  NAND2BXL U10212 ( .AN(n9681), .B(U1_A_r_d0[12]), .Y(n19157) );
  INVXL U10213 ( .A(n14532), .Y(n12379) );
  AND2XL U10214 ( .A(n9681), .B(U1_A_r_d0[12]), .Y(n9682) );
  INVXL U10215 ( .A(n19542), .Y(n7520) );
  INVXL U10216 ( .A(n22774), .Y(n7292) );
  NAND2XL U10217 ( .A(n13399), .B(n24506), .Y(n7600) );
  OR2X2 U10218 ( .A(n22925), .B(n24631), .Y(n22919) );
  INVXL U10219 ( .A(n22935), .Y(n22939) );
  AND2XL U10220 ( .A(n14445), .B(U2_A_i_d[16]), .Y(n21776) );
  NAND2X1 U10221 ( .A(n9681), .B(n5787), .Y(n6991) );
  NAND2BXL U10222 ( .AN(n9681), .B(U1_A_i_d0[12]), .Y(n17236) );
  AND2X2 U10223 ( .A(n24286), .B(n7382), .Y(n6263) );
  OR2X2 U10224 ( .A(n22936), .B(n24649), .Y(n12612) );
  INVXL U10225 ( .A(n17662), .Y(n17657) );
  AND2XL U10226 ( .A(n14445), .B(U2_A_r_d[16]), .Y(n14446) );
  AND2XL U10227 ( .A(n9681), .B(U1_A_i_d0[12]), .Y(n9456) );
  OAI21XL U10228 ( .A0(n9419), .A1(n17557), .B0(n9418), .Y(n17526) );
  OR2X2 U10229 ( .A(n14825), .B(n19541), .Y(n14824) );
  AND2XL U10230 ( .A(n21764), .B(U2_A_i_d[12]), .Y(n21765) );
  OR2X2 U10231 ( .A(n19754), .B(U1_A_r_d0[14]), .Y(n12310) );
  AND2XL U10232 ( .A(n9680), .B(U1_A_i_d0[11]), .Y(n17529) );
  NOR2X1 U10233 ( .A(n19986), .B(n14929), .Y(n14873) );
  OR2X2 U10234 ( .A(n22918), .B(n24631), .Y(n12572) );
  INVXL U10235 ( .A(n19287), .Y(n19280) );
  AOI21X1 U10236 ( .A0(n13573), .A1(n13572), .B0(n13571), .Y(n7190) );
  NAND3BX2 U10237 ( .AN(n13583), .B(n6043), .C(n6042), .Y(n7919) );
  NAND3X2 U10238 ( .A(n7370), .B(n14844), .C(n7371), .Y(n5987) );
  NAND2X2 U10239 ( .A(n6152), .B(n13080), .Y(n7381) );
  OR2X2 U10240 ( .A(n22936), .B(n14548), .Y(n13122) );
  NAND2X1 U10241 ( .A(n7200), .B(n13939), .Y(n6063) );
  NOR2X1 U10242 ( .A(n20007), .B(n19282), .Y(n19281) );
  XOR2XL U10243 ( .A(n23689), .B(n23486), .Y(n23487) );
  INVX2 U10244 ( .A(n25178), .Y(n5863) );
  NAND2X1 U10245 ( .A(n9184), .B(n5821), .Y(n6357) );
  AND2XL U10246 ( .A(n13398), .B(U2_A_i_d[12]), .Y(n14082) );
  INVX1 U10247 ( .A(n26605), .Y(n26354) );
  OR2X2 U10248 ( .A(n14099), .B(U2_A_i_d[17]), .Y(n14098) );
  CLKINVX3 U10249 ( .A(n14099), .Y(n14047) );
  NAND2BXL U10250 ( .AN(n24537), .B(n6981), .Y(n7589) );
  OR2X2 U10251 ( .A(n19984), .B(n14930), .Y(n14874) );
  AOI21X1 U10252 ( .A0(n7890), .A1(n6010), .B0(n7889), .Y(n7191) );
  NAND2X1 U10253 ( .A(n6417), .B(n6416), .Y(n18812) );
  INVXL U10254 ( .A(n18945), .Y(n7378) );
  INVX1 U10255 ( .A(n18495), .Y(n18252) );
  NOR2X1 U10256 ( .A(n13598), .B(n13601), .Y(n6141) );
  OR2X2 U10257 ( .A(n13687), .B(U1_A_i_d0[11]), .Y(n9577) );
  OR2X2 U10258 ( .A(n20001), .B(n19541), .Y(n19540) );
  AND2X2 U10259 ( .A(n24377), .B(n24376), .Y(n24378) );
  NAND2BXL U10260 ( .AN(n24287), .B(n24245), .Y(n7382) );
  AND2X2 U10261 ( .A(n7383), .B(n24246), .Y(n6264) );
  INVX1 U10262 ( .A(n19272), .Y(n5865) );
  OR2X2 U10263 ( .A(n19758), .B(U1_A_r_d0[14]), .Y(n19755) );
  INVX1 U10264 ( .A(n19282), .Y(n5866) );
  OR2X2 U10265 ( .A(n14940), .B(n19311), .Y(n13545) );
  NAND2BX2 U10266 ( .AN(n7506), .B(n6044), .Y(n6043) );
  INVX1 U10267 ( .A(n14955), .Y(n5868) );
  INVXL U10268 ( .A(n20005), .Y(n14828) );
  OR2X2 U10269 ( .A(n13035), .B(n19541), .Y(n13034) );
  INVX1 U10270 ( .A(n14930), .Y(n19985) );
  OR2X2 U10271 ( .A(n8524), .B(n17018), .Y(n6579) );
  OR2X2 U10272 ( .A(n13687), .B(U1_A_r_d0[11]), .Y(n13680) );
  INVXL U10273 ( .A(n9519), .Y(n7673) );
  NAND2X2 U10274 ( .A(n9480), .B(n7628), .Y(n7680) );
  NAND2XL U10275 ( .A(n8663), .B(n16706), .Y(n8665) );
  AND2X2 U10276 ( .A(n18654), .B(n18702), .Y(n18655) );
  OR2X2 U10277 ( .A(n14527), .B(n22887), .Y(n14514) );
  INVXL U10278 ( .A(n19311), .Y(n7885) );
  OR2X2 U10279 ( .A(n19736), .B(U1_A_r_d0[11]), .Y(n12300) );
  OR2X2 U10280 ( .A(n18867), .B(n18866), .Y(n18865) );
  OR2X2 U10281 ( .A(n18820), .B(n18819), .Y(n6935) );
  OR2X2 U10282 ( .A(n19520), .B(n14923), .Y(n13534) );
  NOR2X1 U10283 ( .A(n7175), .B(n7174), .Y(n13602) );
  AND2X2 U10284 ( .A(n6644), .B(n8633), .Y(n6641) );
  INVX4 U10285 ( .A(n5959), .Y(n7146) );
  NAND2XL U10286 ( .A(n18909), .B(n18908), .Y(n18945) );
  NAND3X1 U10287 ( .A(n6051), .B(n7721), .C(n6076), .Y(n6053) );
  XOR2X1 U10288 ( .A(n8584), .B(n8583), .Y(n12311) );
  OR2X2 U10289 ( .A(n19736), .B(U1_A_i_d0[11]), .Y(n8553) );
  INVX2 U10290 ( .A(n9123), .Y(n9135) );
  AND2XL U10291 ( .A(n19745), .B(U1_A_r_d0[12]), .Y(n19746) );
  INVXL U10292 ( .A(n22918), .Y(n22925) );
  INVXL U10293 ( .A(n26816), .Y(n7546) );
  OR2X2 U10294 ( .A(n19745), .B(U1_A_r_d0[12]), .Y(n19735) );
  INVX1 U10295 ( .A(n23935), .Y(n23689) );
  NAND3X1 U10296 ( .A(n12959), .B(n12945), .C(n12977), .Y(n5946) );
  AND2XL U10297 ( .A(n19745), .B(U1_A_i_d0[12]), .Y(n8662) );
  OR2X2 U10298 ( .A(n19970), .B(n14923), .Y(n14903) );
  INVX1 U10299 ( .A(n14935), .Y(n12965) );
  NAND2XL U10300 ( .A(n7748), .B(n7718), .Y(n7717) );
  OR2X2 U10301 ( .A(n14527), .B(n24584), .Y(n12362) );
  NAND2X1 U10302 ( .A(n13619), .B(n13631), .Y(n13620) );
  INVX1 U10303 ( .A(n13614), .Y(n13615) );
  OR2X2 U10304 ( .A(n22887), .B(n13108), .Y(n13097) );
  AND2XL U10305 ( .A(U1_A_i_d0[11]), .B(n19744), .Y(n16705) );
  AND2XL U10306 ( .A(n9668), .B(U1_A_r_d0[7]), .Y(n9669) );
  NAND2XL U10307 ( .A(n18041), .B(n18047), .Y(n18049) );
  NAND2X1 U10308 ( .A(n7247), .B(n12244), .Y(n12223) );
  NAND2X1 U10309 ( .A(n7244), .B(n12254), .Y(n12250) );
  NOR2X1 U10310 ( .A(n26993), .B(n26992), .Y(n27030) );
  ADDFHX2 U10311 ( .A(n21309), .B(n21308), .CI(U2_A_r_d[16]), .CO(n21310), .S(
        n21268) );
  ADDFHX2 U10312 ( .A(n21480), .B(n21479), .CI(U2_A_r_d[19]), .CO(n21481), .S(
        n21426) );
  NAND2XL U10313 ( .A(n9176), .B(n9062), .Y(n6435) );
  ADDFHX1 U10314 ( .A(n21574), .B(n21573), .CI(U2_A_r_d[21]), .CO(n21576), .S(
        n21532) );
  OR2X2 U10315 ( .A(n26823), .B(n26822), .Y(n26821) );
  INVX1 U10316 ( .A(n25226), .Y(n5871) );
  INVX1 U10317 ( .A(n18980), .Y(n5872) );
  INVX1 U10318 ( .A(n18979), .Y(n5873) );
  OR2X2 U10319 ( .A(n9668), .B(U1_A_i_d0[7]), .Y(n9365) );
  ADDFHX2 U10320 ( .A(n18818), .B(n18817), .CI(U2_A_i_d[20]), .CO(n18819), .S(
        n18770) );
  INVXL U10321 ( .A(n12242), .Y(n7250) );
  NOR2X1 U10322 ( .A(n24251), .B(n24250), .Y(n24287) );
  NOR2X1 U10323 ( .A(n24334), .B(n24333), .Y(n24371) );
  OR2X2 U10324 ( .A(n19969), .B(n14902), .Y(n14865) );
  NAND2X1 U10325 ( .A(n20962), .B(n20961), .Y(n21065) );
  NAND2X1 U10326 ( .A(n21019), .B(n21018), .Y(n21064) );
  NOR2XL U10327 ( .A(n7641), .B(n9486), .Y(n7640) );
  NOR2X1 U10328 ( .A(n21124), .B(n21123), .Y(n21180) );
  AOI21XL U10329 ( .A0(n25620), .A1(n25242), .B0(n25470), .Y(n25471) );
  OR2X2 U10330 ( .A(n14074), .B(U2_A_r_d[11]), .Y(n13507) );
  OAI21XL U10331 ( .A0(n19210), .A1(n19490), .B0(n19211), .Y(n13672) );
  NAND2X2 U10332 ( .A(n5948), .B(n7823), .Y(n12959) );
  AND2X2 U10333 ( .A(n13599), .B(n13048), .Y(n6142) );
  OR2X2 U10334 ( .A(n14074), .B(U2_A_i_d[11]), .Y(n14029) );
  OR2X2 U10335 ( .A(n24584), .B(n13108), .Y(n12087) );
  INVXL U10336 ( .A(n13975), .Y(n6723) );
  NAND2X1 U10337 ( .A(n24621), .B(n24617), .Y(n25058) );
  INVXL U10338 ( .A(n13959), .Y(n7493) );
  NAND2X1 U10339 ( .A(n12191), .B(n12209), .Y(n12192) );
  INVX4 U10340 ( .A(n12258), .Y(n5875) );
  NAND2X1 U10341 ( .A(n7894), .B(n14674), .Y(n14840) );
  INVX1 U10342 ( .A(n7830), .Y(n13594) );
  ADDFHX1 U10343 ( .A(n20903), .B(n20902), .CI(U2_A_r_d[9]), .CO(n20904), .S(
        n20857) );
  INVX1 U10344 ( .A(n12262), .Y(n12263) );
  ADDFHX1 U10345 ( .A(n21071), .B(n21070), .CI(U2_A_r_d[12]), .CO(n21072), .S(
        n21019) );
  ADDFHX2 U10346 ( .A(n21191), .B(n21190), .CI(U2_A_r_d[14]), .CO(n21192), .S(
        n21124) );
  ADDFHX2 U10347 ( .A(n26820), .B(n26819), .CI(U2_A_r_d[19]), .CO(n26822), .S(
        n26762) );
  INVXL U10348 ( .A(n12244), .Y(n7246) );
  NAND2X1 U10349 ( .A(n7699), .B(n9477), .Y(n9478) );
  XOR2X1 U10350 ( .A(n13791), .B(n13790), .Y(n14901) );
  NAND2BXL U10351 ( .AN(n9072), .B(n9165), .Y(n7775) );
  OR2X2 U10352 ( .A(n13676), .B(U1_A_r_d0[7]), .Y(n13664) );
  NOR2X2 U10353 ( .A(n26293), .B(n26292), .Y(n26350) );
  NAND2X1 U10354 ( .A(n26357), .B(n26358), .Y(n26455) );
  NAND2X2 U10355 ( .A(n7242), .B(n7241), .Y(n7247) );
  OR2X2 U10356 ( .A(n24610), .B(n24584), .Y(n8839) );
  OR2X2 U10357 ( .A(n14025), .B(U2_A_i_d[7]), .Y(n14015) );
  NAND2XL U10358 ( .A(n14065), .B(U2_A_r_d[5]), .Y(n24553) );
  INVX1 U10359 ( .A(n13644), .Y(n13645) );
  INVX1 U10360 ( .A(n14074), .Y(n5876) );
  NAND2XL U10361 ( .A(n6582), .B(U1_A_i_d0[6]), .Y(n16748) );
  OR2X2 U10362 ( .A(n24611), .B(n24610), .Y(n24585) );
  NAND2X1 U10363 ( .A(n13087), .B(n13567), .Y(n13077) );
  NAND2X1 U10364 ( .A(n14799), .B(n7159), .Y(n6917) );
  OR2X2 U10365 ( .A(n19727), .B(U1_A_i_d0[7]), .Y(n8641) );
  AND2X2 U10366 ( .A(n5822), .B(n13952), .Y(n13933) );
  NAND2X1 U10367 ( .A(n13936), .B(n13935), .Y(n13937) );
  NOR2BX1 U10368 ( .AN(n7886), .B(n7888), .Y(n7220) );
  NOR2X1 U10369 ( .A(n18410), .B(n18409), .Y(n18486) );
  NOR2X1 U10370 ( .A(n6794), .B(n13134), .Y(n6793) );
  INVXL U10371 ( .A(n6791), .Y(n6767) );
  XOR2X2 U10372 ( .A(n11572), .B(n11571), .Y(U2_U0_z0[8]) );
  NOR2X1 U10373 ( .A(n6025), .B(n7432), .Y(n6024) );
  NAND2BX1 U10374 ( .AN(n7259), .B(n6125), .Y(n6124) );
  AOI21X1 U10375 ( .A0(n9155), .A1(n9154), .B0(n6847), .Y(n9187) );
  NAND2X1 U10376 ( .A(n13642), .B(n13652), .Y(n13643) );
  INVXL U10377 ( .A(n9481), .Y(n7642) );
  INVXL U10378 ( .A(n13659), .Y(n13649) );
  AOI21X1 U10379 ( .A0(n17163), .A1(n13833), .B0(n13834), .Y(n17160) );
  OR2X2 U10380 ( .A(n24596), .B(n24595), .Y(n8850) );
  OR2X2 U10381 ( .A(n9093), .B(n9061), .Y(n6316) );
  NAND2X1 U10382 ( .A(n9446), .B(n9445), .Y(n9447) );
  NAND2BXL U10383 ( .AN(n9226), .B(n6443), .Y(n6442) );
  NAND2X1 U10384 ( .A(n12266), .B(n12265), .Y(n12271) );
  INVX1 U10385 ( .A(n14071), .Y(n5877) );
  OR2X2 U10386 ( .A(n13636), .B(n13635), .Y(n13634) );
  NAND2X2 U10387 ( .A(n7867), .B(n7868), .Y(n6084) );
  OR2X2 U10388 ( .A(n12276), .B(n12275), .Y(n12274) );
  INVX1 U10389 ( .A(n14849), .Y(n14684) );
  INVX1 U10390 ( .A(n9526), .Y(n9338) );
  NAND2X1 U10391 ( .A(n6640), .B(n8632), .Y(n6562) );
  NAND2X1 U10392 ( .A(n13957), .B(n13956), .Y(n13961) );
  AND2X2 U10393 ( .A(n19724), .B(n7068), .Y(n6583) );
  ADDFHX2 U10394 ( .A(n18596), .B(n18595), .CI(U2_A_i_d[16]), .CO(n18597), .S(
        n18549) );
  ADDFHX2 U10395 ( .A(n18651), .B(n18650), .CI(U2_A_i_d[17]), .CO(n18652), .S(
        n18598) );
  INVXL U10396 ( .A(n19724), .Y(n6582) );
  AND2X2 U10397 ( .A(n8572), .B(n8571), .Y(n8573) );
  NAND2X1 U10398 ( .A(n8603), .B(n8602), .Y(n8604) );
  INVXL U10399 ( .A(n14844), .Y(n7259) );
  AND2X2 U10400 ( .A(n6665), .B(n8593), .Y(n8594) );
  NAND2BX1 U10401 ( .AN(n14846), .B(n14847), .Y(n6094) );
  AND2X2 U10402 ( .A(n8578), .B(n8577), .Y(n8579) );
  INVX1 U10403 ( .A(n13962), .Y(n5879) );
  NAND2X1 U10404 ( .A(n13144), .B(n13149), .Y(n13145) );
  NAND2XL U10405 ( .A(n9486), .B(n9487), .Y(n7718) );
  NAND2X1 U10406 ( .A(n14266), .B(n14479), .Y(n14480) );
  AND2XL U10407 ( .A(n21751), .B(U2_A_r_d[7]), .Y(n14345) );
  OR2X2 U10408 ( .A(n12296), .B(U1_A_r_d0[7]), .Y(n12286) );
  INVXL U10409 ( .A(n9487), .Y(n7719) );
  AND2X2 U10410 ( .A(n13915), .B(n13914), .Y(n13916) );
  INVX1 U10411 ( .A(n13607), .Y(n13608) );
  NAND2X1 U10412 ( .A(n9236), .B(n12348), .Y(n9237) );
  NAND2X1 U10413 ( .A(n9221), .B(n9231), .Y(n9224) );
  INVXL U10414 ( .A(n9190), .Y(n6852) );
  INVXL U10415 ( .A(n19984), .Y(n5880) );
  NAND2XL U10416 ( .A(n7703), .B(n14430), .Y(n7702) );
  INVXL U10417 ( .A(n12195), .Y(n12197) );
  NAND2X2 U10418 ( .A(n12625), .B(n12619), .Y(n12626) );
  AND2X2 U10419 ( .A(n9470), .B(n9469), .Y(n6958) );
  INVX2 U10420 ( .A(n9188), .Y(n5881) );
  XOR2X1 U10421 ( .A(n12776), .B(n12775), .Y(n19518) );
  NAND2X1 U10422 ( .A(n14475), .B(n14474), .Y(n14476) );
  XOR2X1 U10423 ( .A(n14700), .B(n14699), .Y(n19965) );
  NAND2X1 U10424 ( .A(n13479), .B(n13478), .Y(n13480) );
  NOR2X1 U10425 ( .A(n13618), .B(n13617), .Y(n13632) );
  NAND2X1 U10426 ( .A(n13618), .B(n13617), .Y(n13631) );
  AND2XL U10427 ( .A(n7159), .B(n14798), .Y(n7049) );
  INVXL U10428 ( .A(n14793), .Y(n7442) );
  ADDFHX1 U10429 ( .A(n26291), .B(n26290), .CI(U2_A_r_d[10]), .CO(n26292), .S(
        n26244) );
  XOR2X1 U10430 ( .A(n9359), .B(n9358), .Y(n13674) );
  INVXL U10431 ( .A(n16777), .Y(n8644) );
  INVX1 U10432 ( .A(n13637), .Y(n13638) );
  NAND2X1 U10433 ( .A(n13979), .B(n13978), .Y(n13980) );
  INVXL U10434 ( .A(n7159), .Y(n7891) );
  NAND2X1 U10435 ( .A(n13013), .B(n13043), .Y(n13014) );
  INVXL U10436 ( .A(n9438), .Y(n7615) );
  NAND2X1 U10437 ( .A(n13439), .B(n13438), .Y(n13440) );
  OR2X2 U10438 ( .A(n25243), .B(U2_A_r_d[7]), .Y(n25242) );
  XNOR2X1 U10439 ( .A(n8920), .B(n8919), .Y(n24600) );
  NOR2BX1 U10440 ( .AN(U2_U0_y0[36]), .B(n6411), .Y(n24331) );
  NAND2X1 U10441 ( .A(n13010), .B(n13060), .Y(n13011) );
  NAND2BXL U10442 ( .AN(n9212), .B(n9215), .Y(n6443) );
  INVX1 U10443 ( .A(n9231), .Y(n9232) );
  ADDFHX1 U10444 ( .A(n18189), .B(n18188), .CI(U2_A_i_d[9]), .CO(n18190), .S(
        n18145) );
  NAND2X1 U10445 ( .A(n9215), .B(n9225), .Y(n9218) );
  NAND2BXL U10446 ( .AN(n9213), .B(n9215), .Y(n6444) );
  OR2X2 U10447 ( .A(n9343), .B(n9342), .Y(n9341) );
  INVXL U10448 ( .A(n9177), .Y(n6433) );
  AND2X2 U10449 ( .A(n13444), .B(n13443), .Y(n6922) );
  XNOR2X1 U10450 ( .A(n12127), .B(n12126), .Y(n13101) );
  INVXL U10451 ( .A(n13575), .Y(n7279) );
  NAND2X1 U10452 ( .A(n5764), .B(n9314), .Y(n9440) );
  NAND2X1 U10453 ( .A(n11516), .B(n11515), .Y(n11517) );
  NAND2XL U10454 ( .A(n13387), .B(n7607), .Y(n7606) );
  INVXL U10455 ( .A(n9362), .Y(n9359) );
  INVXL U10456 ( .A(n14842), .Y(n7805) );
  AND2XL U10457 ( .A(n9397), .B(U1_A_r_d0[1]), .Y(n9652) );
  NAND2X1 U10458 ( .A(n13648), .B(n13647), .Y(n13658) );
  OR2X2 U10459 ( .A(n19369), .B(n14912), .Y(n13535) );
  NAND2XL U10460 ( .A(n13577), .B(n13580), .Y(n7922) );
  INVXL U10461 ( .A(n8596), .Y(n8598) );
  INVXL U10462 ( .A(n7184), .Y(n7464) );
  NOR2X1 U10463 ( .A(n13985), .B(n13984), .Y(n13990) );
  INVXL U10464 ( .A(n13978), .Y(n6721) );
  INVX1 U10465 ( .A(n14021), .Y(n14062) );
  INVXL U10466 ( .A(n13580), .Y(n7923) );
  NAND2X1 U10467 ( .A(n14680), .B(n14679), .Y(n14847) );
  NOR2X1 U10468 ( .A(n23527), .B(n23526), .Y(n23573) );
  AOI21X1 U10469 ( .A0(n7883), .A1(n7884), .B0(n6132), .Y(n6131) );
  NAND2X1 U10470 ( .A(n12138), .B(n6781), .Y(n6786) );
  NAND2X1 U10471 ( .A(n9097), .B(n9105), .Y(n9098) );
  INVXL U10472 ( .A(n9433), .Y(n9435) );
  INVXL U10473 ( .A(n13137), .Y(n6792) );
  INVX1 U10474 ( .A(n19951), .Y(n5883) );
  XNOR3X2 U10475 ( .A(n5781), .B(n23871), .C(n23870), .Y(n23798) );
  INVXL U10476 ( .A(n9473), .Y(n9475) );
  AND2X2 U10477 ( .A(n8969), .B(n8968), .Y(n8970) );
  AOI211XL U10478 ( .A0(n5826), .A1(n27787), .B0(n28625), .C0(n27262), .Y(
        n27263) );
  NAND2X1 U10479 ( .A(n13611), .B(n13610), .Y(n13625) );
  AOI211XL U10480 ( .A0(n5826), .A1(n27775), .B0(n28625), .C0(n27254), .Y(
        n27255) );
  AND2X2 U10481 ( .A(n12547), .B(n12560), .Y(n12548) );
  OAI21XL U10482 ( .A0(n9080), .A1(n9088), .B0(n9081), .Y(n9154) );
  INVXL U10483 ( .A(n14424), .Y(n7705) );
  AND2XL U10484 ( .A(n9397), .B(U1_A_i_d0[1]), .Y(n9398) );
  INVXL U10485 ( .A(n9469), .Y(n7690) );
  NAND2X1 U10486 ( .A(n13878), .B(n13893), .Y(n13879) );
  NAND2XL U10487 ( .A(n14423), .B(n14431), .Y(n7703) );
  AND2X2 U10488 ( .A(n9075), .B(n9165), .Y(n9076) );
  OR2X2 U10489 ( .A(n13630), .B(n13629), .Y(n13628) );
  AOI211XL U10490 ( .A0(n5826), .A1(n27635), .B0(n28452), .C0(n27169), .Y(
        n27170) );
  AND2X2 U10491 ( .A(n9086), .B(n9085), .Y(n9087) );
  NAND2X1 U10492 ( .A(n14467), .B(n14466), .Y(n14468) );
  NAND2X1 U10493 ( .A(n9346), .B(n9345), .Y(n9543) );
  NAND2X1 U10494 ( .A(n9334), .B(n9333), .Y(n9522) );
  AND2X2 U10495 ( .A(n13860), .B(n13871), .Y(n13861) );
  INVX1 U10496 ( .A(n9185), .Y(n6358) );
  NAND2X1 U10497 ( .A(n14433), .B(n14439), .Y(n14440) );
  NAND2X2 U10498 ( .A(n14246), .B(n14396), .Y(n7595) );
  NAND2X1 U10499 ( .A(n8637), .B(n8636), .Y(n8638) );
  INVX1 U10500 ( .A(n9201), .Y(n9202) );
  NAND2BXL U10501 ( .AN(n8627), .B(n8633), .Y(n6640) );
  AND2X2 U10502 ( .A(n14436), .B(n14435), .Y(n14437) );
  INVX1 U10503 ( .A(n13159), .Y(n13160) );
  ADDHXL U10504 ( .A(U0_U2_y2[39]), .B(U0_U2_y0[39]), .CO(n12358), .S(n12281)
         );
  XNOR2X1 U10505 ( .A(n13816), .B(n13815), .Y(n14904) );
  AND2X2 U10506 ( .A(n8997), .B(n9014), .Y(n8998) );
  XNOR2X1 U10507 ( .A(n14365), .B(n14364), .Y(n25235) );
  AOI211XL U10508 ( .A0(n5826), .A1(n28613), .B0(n28625), .C0(n28043), .Y(
        n28044) );
  NAND2X2 U10509 ( .A(n9308), .B(n9309), .Y(n9427) );
  AND2XL U10510 ( .A(n22727), .B(n13098), .Y(n22421) );
  NAND2X1 U10511 ( .A(n12631), .B(n12630), .Y(n12638) );
  AOI211XL U10512 ( .A0(n5827), .A1(n27732), .B0(n28543), .C0(n27731), .Y(
        n27733) );
  XNOR2X1 U10513 ( .A(n9379), .B(n9378), .Y(n13670) );
  AOI211XL U10514 ( .A0(n27631), .A1(n27708), .B0(n28515), .C0(n27707), .Y(
        n27709) );
  INVX1 U10515 ( .A(n19709), .Y(n16780) );
  INVX1 U10516 ( .A(n13134), .Y(n5885) );
  NAND2X2 U10517 ( .A(n6345), .B(n6346), .Y(n9073) );
  AND2XL U10518 ( .A(n21735), .B(U2_A_i_d[1]), .Y(n21736) );
  XNOR2X1 U10519 ( .A(n9408), .B(n9407), .Y(n13669) );
  OR2X2 U10520 ( .A(n13667), .B(U1_A_r_d0[1]), .Y(n13666) );
  AOI211XL U10521 ( .A0(n27631), .A1(n28329), .B0(n28328), .C0(n28327), .Y(
        n28330) );
  AOI211XL U10522 ( .A0(n27631), .A1(n28343), .B0(n28342), .C0(n28341), .Y(
        n28344) );
  AOI211XL U10523 ( .A0(n27631), .A1(n28350), .B0(n28349), .C0(n28348), .Y(
        n28351) );
  AOI211XL U10524 ( .A0(n27631), .A1(n27501), .B0(n7120), .C0(n27500), .Y(
        n27502) );
  XOR2XL U10525 ( .A(U1_U2_y0[40]), .B(U1_U2_y1[40]), .Y(n13662) );
  OR2X2 U10526 ( .A(n13157), .B(n13156), .Y(n13155) );
  NOR2X1 U10527 ( .A(n9309), .B(n9308), .Y(n9420) );
  NAND2X1 U10528 ( .A(n11499), .B(n11498), .Y(n11500) );
  OR2X2 U10529 ( .A(n13176), .B(n13175), .Y(n13174) );
  AOI211XL U10530 ( .A0(n27631), .A1(n28558), .B0(n28557), .C0(n28556), .Y(
        n28559) );
  OR2XL U10531 ( .A(n14057), .B(U2_A_i_d[1]), .Y(n14059) );
  NAND2X1 U10532 ( .A(n13163), .B(n13162), .Y(n13172) );
  INVXL U10533 ( .A(n13162), .Y(n6449) );
  AOI211XL U10534 ( .A0(n5798), .A1(n28365), .B0(n28364), .C0(n28363), .Y(
        n28366) );
  CLKINVX3 U10535 ( .A(n23870), .Y(n5888) );
  XOR2X1 U10536 ( .A(n13190), .B(n13189), .Y(n13191) );
  NAND2X1 U10537 ( .A(n8451), .B(n8450), .Y(n8624) );
  NAND2X1 U10538 ( .A(n8538), .B(n8537), .Y(n8539) );
  AND2X2 U10539 ( .A(n8550), .B(n8549), .Y(n8551) );
  INVX1 U10540 ( .A(n23742), .Y(n18360) );
  INVX1 U10541 ( .A(n25458), .Y(n25285) );
  AND2XL U10542 ( .A(n20179), .B(n14905), .Y(n20455) );
  AND2XL U10543 ( .A(n21735), .B(U2_A_r_d[1]), .Y(n14325) );
  NOR2X1 U10544 ( .A(n13143), .B(n13142), .Y(n13150) );
  NAND2X1 U10545 ( .A(n9159), .B(n9158), .Y(n9185) );
  INVX1 U10546 ( .A(n9186), .Y(n5889) );
  OR2X2 U10547 ( .A(n13667), .B(U1_A_i_d0[1]), .Y(n9570) );
  AND2X1 U10548 ( .A(n12706), .B(n12778), .Y(n6939) );
  OR2XL U10549 ( .A(n14057), .B(U2_A_r_d[1]), .Y(n13350) );
  AND2XL U10550 ( .A(n16932), .B(n14905), .Y(n17163) );
  XNOR2X1 U10551 ( .A(n12825), .B(n12824), .Y(n19363) );
  INVX1 U10552 ( .A(n14905), .Y(n20180) );
  NOR2X1 U10553 ( .A(n13795), .B(n13792), .Y(n13847) );
  NAND2X1 U10554 ( .A(n8448), .B(n8447), .Y(n8622) );
  INVX1 U10555 ( .A(n8621), .Y(n5890) );
  NOR2X1 U10556 ( .A(n9039), .B(n9038), .Y(n9153) );
  INVX1 U10557 ( .A(n13665), .Y(n19231) );
  INVXL U10558 ( .A(n9013), .Y(n9002) );
  CLKINVX3 U10559 ( .A(n9017), .Y(n5891) );
  NAND2X1 U10560 ( .A(n14660), .B(n14661), .Y(n14818) );
  AOI211XL U10561 ( .A0(n5798), .A1(n28481), .B0(n28480), .C0(n28479), .Y(
        n28482) );
  NAND2X1 U10562 ( .A(n12944), .B(n12976), .Y(n12945) );
  AND2X2 U10563 ( .A(n9182), .B(n9181), .Y(n9195) );
  AND2X2 U10564 ( .A(n13418), .B(n13417), .Y(n13419) );
  INVX1 U10565 ( .A(n13098), .Y(n25449) );
  XOR2X1 U10566 ( .A(n14273), .B(n14272), .Y(n14274) );
  INVX1 U10567 ( .A(n13078), .Y(n5892) );
  INVXL U10568 ( .A(n8951), .Y(n7222) );
  NAND3X2 U10569 ( .A(n6413), .B(n7231), .C(n13314), .Y(n6412) );
  OR2X2 U10570 ( .A(n13287), .B(n13286), .Y(n13285) );
  INVXL U10571 ( .A(n8966), .Y(n8828) );
  NAND2X1 U10572 ( .A(n12957), .B(n12977), .Y(n12958) );
  INVXL U10573 ( .A(n9108), .Y(n9110) );
  NAND2X1 U10574 ( .A(n14265), .B(n14264), .Y(n14474) );
  OR2X2 U10575 ( .A(n13293), .B(n13292), .Y(n13291) );
  INVXL U10576 ( .A(n9165), .Y(n7774) );
  NAND2X1 U10577 ( .A(n13290), .B(n13289), .Y(n13478) );
  NAND2X1 U10578 ( .A(n9198), .B(n9197), .Y(n9212) );
  NAND2X1 U10579 ( .A(n13411), .B(n13410), .Y(n13412) );
  NAND2X1 U10580 ( .A(n13390), .B(n13389), .Y(n13391) );
  OAI21X1 U10581 ( .A0(n8897), .A1(n8948), .B0(n8952), .Y(n8825) );
  OR2X2 U10582 ( .A(n14268), .B(n14267), .Y(n14266) );
  INVXL U10583 ( .A(n14809), .Y(n14811) );
  NAND2X2 U10584 ( .A(n12067), .B(n12088), .Y(n12134) );
  NOR2X1 U10585 ( .A(n12078), .B(n12081), .Y(n12133) );
  INVXL U10586 ( .A(n13016), .Y(n13018) );
  INVXL U10587 ( .A(n13371), .Y(n7084) );
  OR2XL U10588 ( .A(n14018), .B(U2_A_i_d[1]), .Y(n14017) );
  NOR2X1 U10589 ( .A(n8458), .B(n8457), .Y(n8635) );
  NAND2X1 U10590 ( .A(n13785), .B(n13786), .Y(n13793) );
  INVX1 U10591 ( .A(n11535), .Y(n11440) );
  NAND2X1 U10592 ( .A(n13874), .B(n13875), .Y(n13893) );
  NAND2X1 U10593 ( .A(n8458), .B(n8457), .Y(n8636) );
  INVXL U10594 ( .A(n13388), .Y(n13390) );
  OR2X2 U10595 ( .A(n9217), .B(n9216), .Y(n9215) );
  NAND2X1 U10596 ( .A(n11445), .B(U2_B_r[18]), .Y(n11515) );
  AND2X2 U10597 ( .A(n9374), .B(n9373), .Y(n9375) );
  INVXL U10598 ( .A(n8455), .Y(n6522) );
  XNOR2X1 U10599 ( .A(n8519), .B(n8518), .Y(n12290) );
  NAND2X1 U10600 ( .A(n8940), .B(n8939), .Y(n8981) );
  INVXL U10601 ( .A(n8582), .Y(n6656) );
  NAND2X1 U10602 ( .A(n13784), .B(n13783), .Y(n13794) );
  NAND2BXL U10603 ( .AN(n8931), .B(n8938), .Y(n7290) );
  NOR2X1 U10604 ( .A(n11453), .B(U2_B_r[23]), .Y(n11483) );
  INVX1 U10605 ( .A(n13370), .Y(n13365) );
  INVXL U10606 ( .A(n13389), .Y(n7609) );
  OR2X2 U10607 ( .A(n12288), .B(U1_A_i_d0[1]), .Y(n8510) );
  INVX1 U10608 ( .A(n12974), .Y(n12957) );
  AND2X2 U10609 ( .A(n14372), .B(n14371), .Y(n14373) );
  OAI211XL U10610 ( .A0(n7125), .A1(n16464), .B0(n16463), .C0(n16462), .Y(
        n16465) );
  INVX1 U10611 ( .A(n14289), .Y(n14286) );
  OAI211XL U10612 ( .A0(n7125), .A1(n16402), .B0(n16401), .C0(n16400), .Y(
        n16403) );
  XNOR2X1 U10613 ( .A(n14715), .B(n14714), .Y(n19960) );
  OAI211XL U10614 ( .A0(n7125), .A1(n16394), .B0(n16393), .C0(n16392), .Y(
        n16395) );
  NAND2X1 U10615 ( .A(n8827), .B(n8826), .Y(n8965) );
  OAI211XL U10616 ( .A0(n7125), .A1(n16414), .B0(n16413), .C0(n16412), .Y(
        n16415) );
  OR2X2 U10617 ( .A(n25281), .B(U2_A_r_d[1]), .Y(n25280) );
  INVX1 U10618 ( .A(n9090), .Y(n5894) );
  XNOR2X1 U10619 ( .A(n12526), .B(n12525), .Y(n22890) );
  CLKINVX4 U10620 ( .A(n9931), .Y(U1_U2_z2[16]) );
  NOR2X2 U10621 ( .A(n14656), .B(n7044), .Y(n14776) );
  INVX1 U10622 ( .A(n9127), .Y(n5895) );
  INVXL U10623 ( .A(n12977), .Y(n7820) );
  NAND2XL U10624 ( .A(n12974), .B(n12977), .Y(n7819) );
  INVX1 U10625 ( .A(n7798), .Y(n7449) );
  NAND2X2 U10626 ( .A(n14249), .B(n14248), .Y(n14439) );
  NOR2X2 U10627 ( .A(n6467), .B(n7632), .Y(n9319) );
  XNOR2X1 U10628 ( .A(n14335), .B(n14334), .Y(n25275) );
  OR2X2 U10629 ( .A(n12288), .B(U1_A_r_d0[1]), .Y(n12287) );
  OAI211XL U10630 ( .A0(n7125), .A1(n16386), .B0(n16385), .C0(n16384), .Y(
        n16387) );
  OAI211XL U10631 ( .A0(n7125), .A1(n16361), .B0(n16360), .C0(n16359), .Y(
        n16362) );
  INVX1 U10632 ( .A(n9036), .Y(n6345) );
  INVX1 U10633 ( .A(n9035), .Y(n6346) );
  INVXL U10634 ( .A(U1_U2_y0[33]), .Y(n7905) );
  OR2X2 U10635 ( .A(n25281), .B(U2_A_i_d[1]), .Y(n21942) );
  XOR2X1 U10636 ( .A(n8460), .B(n8459), .Y(n8461) );
  NOR2X2 U10637 ( .A(n13280), .B(n13279), .Y(n13432) );
  INVXL U10638 ( .A(n11539), .Y(n11534) );
  ADDHXL U10639 ( .A(U0_U0_y1[39]), .B(U0_U0_y0[39]), .CO(n13297), .S(n13295)
         );
  NAND2X2 U10640 ( .A(n13273), .B(n13274), .Y(n13447) );
  CLKBUFX8 U10641 ( .A(B0_addr[3]), .Y(n7124) );
  NAND2X1 U10642 ( .A(n8984), .B(n8983), .Y(n9045) );
  INVX1 U10643 ( .A(n14820), .Y(n5897) );
  INVX2 U10644 ( .A(n12159), .Y(n5898) );
  ADDHX2 U10645 ( .A(U0_U0_y2[32]), .B(U0_U0_y0[32]), .CO(n14253), .S(n14250)
         );
  CMPR22X1 U10646 ( .A(U0_U0_y2[34]), .B(U0_U0_y0[34]), .CO(n14258), .S(n14254) );
  INVXL U10647 ( .A(n14766), .Y(n7859) );
  INVXL U10648 ( .A(n7681), .Y(n7714) );
  NOR2X2 U10649 ( .A(n12898), .B(n12897), .Y(n12939) );
  CLKINVX8 U10650 ( .A(n11877), .Y(B0_addr[5]) );
  NAND2X1 U10651 ( .A(n10972), .B(n6378), .Y(n10978) );
  CLKINVX8 U10652 ( .A(n11882), .Y(B0_addr[1]) );
  CMPR22X1 U10653 ( .A(U0_U0_y1[33]), .B(U0_U0_y0[33]), .CO(n13280), .S(n13277) );
  XOR2X1 U10654 ( .A(U0_U1_y1[24]), .B(U0_U1_y0[24]), .Y(n8942) );
  INVXL U10655 ( .A(n9357), .Y(n7431) );
  CLKINVX8 U10656 ( .A(n11888), .Y(B1_addr[0]) );
  BUFX12 U10657 ( .A(n28055), .Y(n27959) );
  INVXL U10658 ( .A(n11443), .Y(n11523) );
  NAND2X2 U10659 ( .A(U2_B_i[13]), .B(n6170), .Y(n6989) );
  CLKINVX8 U10660 ( .A(n11884), .Y(B2_addr[1]) );
  AOI21X1 U10661 ( .A0(n8809), .A1(n8906), .B0(n8808), .Y(n8937) );
  INVX1 U10662 ( .A(n14691), .Y(n7451) );
  INVXL U10663 ( .A(n13314), .Y(n6549) );
  INVX1 U10664 ( .A(n8525), .Y(n5899) );
  INVX1 U10665 ( .A(n12803), .Y(n6027) );
  NOR2X2 U10666 ( .A(n12704), .B(n12705), .Y(n12780) );
  NOR2X2 U10667 ( .A(n12813), .B(n12811), .Y(n12763) );
  AND2X2 U10668 ( .A(U0_U2_y0[24]), .B(U0_U2_y2[24]), .Y(n6752) );
  NAND2X1 U10669 ( .A(n9303), .B(n9302), .Y(n9354) );
  NAND2X1 U10670 ( .A(n8747), .B(n8746), .Y(n8823) );
  INVX1 U10671 ( .A(n14690), .Y(n14740) );
  AND4XL U10672 ( .A(n11692), .B(n11691), .C(n11690), .D(n11689), .Y(n5273) );
  AND4XL U10673 ( .A(n11659), .B(n11658), .C(n11657), .D(n11656), .Y(n5271) );
  AND4XL U10674 ( .A(n11704), .B(n11703), .C(n11702), .D(n11701), .Y(n5267) );
  AND4XL U10675 ( .A(n11787), .B(n11786), .C(n11785), .D(n11784), .Y(n5257) );
  AND4XL U10676 ( .A(n11827), .B(n11826), .C(n11825), .D(n11824), .Y(n5255) );
  NOR2X1 U10677 ( .A(n14228), .B(n14227), .Y(n14349) );
  AND4XL U10678 ( .A(n11767), .B(n11766), .C(n11765), .D(n11764), .Y(n5249) );
  NAND2X1 U10679 ( .A(n14230), .B(n14229), .Y(n14352) );
  AND4XL U10680 ( .A(n11847), .B(n11846), .C(n11845), .D(n11844), .Y(n5245) );
  AND4XL U10681 ( .A(n11731), .B(n11730), .C(n11729), .D(n11728), .Y(n5243) );
  AND4XL U10682 ( .A(n11683), .B(n11682), .C(n11681), .D(n11680), .Y(n5241) );
  AND4XL U10683 ( .A(n11747), .B(n11746), .C(n11745), .D(n11744), .Y(n5239) );
  AND4XL U10684 ( .A(n11775), .B(n11774), .C(n11773), .D(n11772), .Y(n5289) );
  AND4XL U10685 ( .A(n11667), .B(n11666), .C(n11665), .D(n11664), .Y(n5287) );
  AND4XL U10686 ( .A(n11851), .B(n11850), .C(n11849), .D(n11848), .Y(n5285) );
  NAND2X1 U10687 ( .A(n14651), .B(n14650), .Y(n14763) );
  AND4XL U10688 ( .A(n11799), .B(n11798), .C(n11797), .D(n11796), .Y(n5283) );
  AND4XL U10689 ( .A(n11771), .B(n11770), .C(n11769), .D(n11768), .Y(n5281) );
  AND4XL U10690 ( .A(n11700), .B(n11699), .C(n11698), .D(n11697), .Y(n5279) );
  AND4XL U10691 ( .A(n11755), .B(n11754), .C(n11753), .D(n11752), .Y(n5275) );
  NOR2X1 U10692 ( .A(n13836), .B(n13837), .Y(n13802) );
  ADDHXL U10693 ( .A(U2_U0_y2[13]), .B(n23132), .CO(n23175), .S(n21730) );
  NOR2X1 U10694 ( .A(n8811), .B(n8810), .Y(n8830) );
  NAND2X1 U10695 ( .A(n12062), .B(n12063), .Y(n12098) );
  AND2X2 U10696 ( .A(U0_U0_y1[23]), .B(U0_U0_y0[23]), .Y(n7569) );
  NOR2X2 U10697 ( .A(n14647), .B(n14646), .Y(n14767) );
  OAI21X1 U10698 ( .A0(n14692), .A1(n14697), .B0(n14693), .Y(n14701) );
  CLKINVX8 U10699 ( .A(n11890), .Y(B1_addr[2]) );
  AND4XL U10700 ( .A(n11872), .B(n11871), .C(n11870), .D(n11869), .Y(n5201) );
  AND4XL U10701 ( .A(n11803), .B(n11802), .C(n11801), .D(n11800), .Y(n5205) );
  AND2X2 U10702 ( .A(U0_U2_y1[24]), .B(U0_U2_y0[24]), .Y(n7559) );
  AND4XL U10703 ( .A(n11843), .B(n11842), .C(n11841), .D(n11840), .Y(n5213) );
  XOR2X1 U10704 ( .A(n11103), .B(n7010), .Y(U1_U1_z0[17]) );
  XOR2X2 U10705 ( .A(n6684), .B(n11300), .Y(U0_U1_z0[15]) );
  AND4XL U10706 ( .A(n11779), .B(n11778), .C(n11777), .D(n11776), .Y(n5233) );
  AND4XL U10707 ( .A(n11807), .B(n11806), .C(n11805), .D(n11804), .Y(n5219) );
  NOR2X1 U10708 ( .A(n12765), .B(n12764), .Y(n12786) );
  AND4XL U10709 ( .A(n11688), .B(n11687), .C(n11686), .D(n11685), .Y(n5229) );
  AND4XL U10710 ( .A(n11839), .B(n11838), .C(n11837), .D(n11836), .Y(n5221) );
  AND4XL U10711 ( .A(n11859), .B(n11858), .C(n11857), .D(n11856), .Y(n5225) );
  INVXL U10712 ( .A(n12472), .Y(n5902) );
  NAND2X2 U10713 ( .A(n6171), .B(n8690), .Y(U2_B_i[13]) );
  AND4XL U10714 ( .A(n11783), .B(n11782), .C(n11781), .D(n11780), .Y(n5223) );
  AND4XL U10715 ( .A(n11696), .B(n11695), .C(n11694), .D(n11693), .Y(n5231) );
  AND4XL U10716 ( .A(n11759), .B(n11758), .C(n11757), .D(n11756), .Y(n5237) );
  AND4XL U10717 ( .A(n11739), .B(n11738), .C(n11737), .D(n11736), .Y(n5227) );
  AND4XL U10718 ( .A(n11795), .B(n11794), .C(n11793), .D(n11792), .Y(n5235) );
  BUFX3 U10719 ( .A(n5750), .Y(n7119) );
  NAND2X1 U10720 ( .A(n12765), .B(n12764), .Y(n12788) );
  OAI21X1 U10721 ( .A0(n11296), .A1(n11348), .B0(n6685), .Y(n6684) );
  NOR2X2 U10722 ( .A(n13778), .B(n13777), .Y(n13837) );
  INVXL U10723 ( .A(n6578), .Y(n6571) );
  INVX1 U10724 ( .A(U2_B_i[16]), .Y(n11441) );
  OAI21X2 U10725 ( .A0(n6194), .A1(n11427), .B0(n11413), .Y(U2_B_i[21]) );
  AND4XL U10726 ( .A(n11811), .B(n11810), .C(n11809), .D(n11808), .Y(n5215) );
  AND4XL U10727 ( .A(n11671), .B(n11670), .C(n11669), .D(n11668), .Y(n5211) );
  AND4XL U10728 ( .A(n11815), .B(n11814), .C(n11813), .D(n11812), .Y(n5209) );
  AND4XL U10729 ( .A(n11863), .B(n11862), .C(n11861), .D(n11860), .Y(n5207) );
  AND4XL U10730 ( .A(n11868), .B(n11867), .C(n11866), .D(n11865), .Y(n5203) );
  AND4XL U10731 ( .A(n11714), .B(n11713), .C(n11712), .D(n11711), .Y(n5199) );
  AND4XL U10732 ( .A(n11743), .B(n11742), .C(n11741), .D(n11740), .Y(n5197) );
  AND4XL U10733 ( .A(n11835), .B(n11834), .C(n11833), .D(n11832), .Y(n5195) );
  AND4XL U10734 ( .A(n11791), .B(n11790), .C(n11789), .D(n11788), .Y(n5193) );
  AND4XL U10735 ( .A(n11727), .B(n11726), .C(n11725), .D(n11724), .Y(n5191) );
  AND4XL U10736 ( .A(n11718), .B(n11717), .C(n11716), .D(n11715), .Y(n5189) );
  AND4XL U10737 ( .A(n11823), .B(n11822), .C(n11821), .D(n11820), .Y(n5263) );
  AND4XL U10738 ( .A(n11763), .B(n11762), .C(n11761), .D(n11760), .Y(n5265) );
  AND4XL U10739 ( .A(n11675), .B(n11674), .C(n11673), .D(n11672), .Y(n5253) );
  ADDHXL U10740 ( .A(U2_U0_y1[13]), .B(n25800), .CO(n25846), .S(n24409) );
  AND4XL U10741 ( .A(n11751), .B(n11750), .C(n11749), .D(n11748), .Y(n5251) );
  AND4XL U10742 ( .A(n11708), .B(n11707), .C(n11706), .D(n11705), .Y(n5269) );
  AND4XL U10743 ( .A(n11855), .B(n11854), .C(n11853), .D(n11852), .Y(n5259) );
  AND4XL U10744 ( .A(n11831), .B(n11830), .C(n11829), .D(n11828), .Y(n5291) );
  NAND2X1 U10745 ( .A(n8416), .B(n8415), .Y(n8465) );
  INVX1 U10746 ( .A(n11886), .Y(n11887) );
  AND4XL U10747 ( .A(n11663), .B(n11662), .C(n11661), .D(n11660), .Y(n5261) );
  INVXL U10748 ( .A(U0_U1_y0[19]), .Y(n7772) );
  NOR2X1 U10749 ( .A(n12461), .B(n12460), .Y(n12518) );
  INVXL U10750 ( .A(n6763), .Y(n12109) );
  INVX2 U10751 ( .A(n13301), .Y(n5903) );
  CLKINVX3 U10752 ( .A(n27497), .Y(n27560) );
  NOR2X1 U10753 ( .A(n12123), .B(n12121), .Y(n12088) );
  NAND2X1 U10754 ( .A(n8742), .B(n8743), .Y(n8917) );
  NAND2X1 U10755 ( .A(n8741), .B(n8740), .Y(n8841) );
  NOR2X1 U10756 ( .A(n12760), .B(n12759), .Y(n12811) );
  INVX1 U10757 ( .A(n11875), .Y(n11876) );
  INVX1 U10758 ( .A(n7087), .Y(n7088) );
  NOR2XL U10759 ( .A(n5812), .B(U1_pipe7[26]), .Y(n7485) );
  INVXL U10760 ( .A(n25091), .Y(n6361) );
  NAND2X1 U10761 ( .A(n7550), .B(U2_B_i[1]), .Y(n6296) );
  NAND2X1 U10762 ( .A(U2_B_i[2]), .B(n6323), .Y(n11597) );
  INVXL U10763 ( .A(n5804), .Y(n6002) );
  NOR2X1 U10764 ( .A(n13249), .B(n13248), .Y(n13321) );
  INVX1 U10765 ( .A(n7604), .Y(n6486) );
  AOI21XL U10766 ( .A0(n9760), .A1(n6391), .B0(n9759), .Y(n9761) );
  NAND2XL U10767 ( .A(n13241), .B(n13334), .Y(n13243) );
  NAND2BX1 U10768 ( .AN(n13817), .B(n13819), .Y(n6065) );
  CLKINVX3 U10769 ( .A(n11107), .Y(n11172) );
  NAND2BXL U10770 ( .AN(n8859), .B(n8861), .Y(n6371) );
  NAND2X1 U10771 ( .A(n8739), .B(n8738), .Y(n8852) );
  OR2X1 U10772 ( .A(n5812), .B(U0_pipe12[27]), .Y(n7237) );
  NAND2BX1 U10773 ( .AN(n12826), .B(n12828), .Y(n6147) );
  NAND2X1 U10774 ( .A(n14219), .B(n14218), .Y(n14283) );
  INVXL U10775 ( .A(n5812), .Y(n6120) );
  NOR2XL U10776 ( .A(n7759), .B(n7757), .Y(n7756) );
  OR2X1 U10777 ( .A(n24784), .B(U0_pipe2[27]), .Y(n7577) );
  NAND3X2 U10778 ( .A(n11013), .B(n8316), .C(n6375), .Y(n6207) );
  OAI21XL U10779 ( .A0(n6867), .A1(n10650), .B0(n10651), .Y(n10649) );
  NAND2BXL U10780 ( .AN(U1_pipe9[26]), .B(n5837), .Y(n7490) );
  INVXL U10781 ( .A(U2_B_i[8]), .Y(n9628) );
  INVX4 U10782 ( .A(n5924), .Y(n5905) );
  INVXL U10783 ( .A(U2_B_r[13]), .Y(n6170) );
  NOR2X1 U10784 ( .A(n9290), .B(n9291), .Y(n9402) );
  INVXL U10785 ( .A(n9619), .Y(n7742) );
  AOI21X1 U10786 ( .A0(n6554), .A1(n10662), .B0(n10655), .Y(n10660) );
  INVX4 U10787 ( .A(n5924), .Y(n5906) );
  INVX4 U10788 ( .A(n5924), .Y(n5907) );
  INVX4 U10789 ( .A(n5924), .Y(n5908) );
  INVX1 U10790 ( .A(n12827), .Y(n6146) );
  NOR2X1 U10791 ( .A(n14214), .B(n14213), .Y(n14296) );
  INVX4 U10792 ( .A(n5924), .Y(n5910) );
  NOR2X1 U10793 ( .A(n14210), .B(n14209), .Y(n14329) );
  INVX4 U10794 ( .A(n11957), .Y(n5911) );
  NAND2X1 U10795 ( .A(n8409), .B(n8410), .Y(n8489) );
  INVX4 U10796 ( .A(n5924), .Y(n5912) );
  NOR2X1 U10797 ( .A(n8406), .B(n8405), .Y(n8513) );
  INVX4 U10798 ( .A(n5924), .Y(n5913) );
  INVX4 U10799 ( .A(n7126), .Y(n5914) );
  INVX1 U10800 ( .A(n13818), .Y(n6069) );
  AOI21X1 U10801 ( .A0(n9809), .A1(n9808), .B0(n9779), .Y(n9783) );
  BUFX3 U10802 ( .A(n11864), .Y(n11676) );
  XOR2X1 U10803 ( .A(n11041), .B(n11040), .Y(U0_U2_z0[2]) );
  INVX4 U10804 ( .A(n11891), .Y(n5916) );
  INVX4 U10805 ( .A(n5924), .Y(n5917) );
  XNOR2X1 U10806 ( .A(n10669), .B(n10668), .Y(U1_U0_z0[3]) );
  BUFX12 U10807 ( .A(n11929), .Y(n28252) );
  INVXL U10808 ( .A(n10191), .Y(n10192) );
  INVXL U10809 ( .A(n9380), .Y(n5919) );
  BUFX3 U10810 ( .A(T1_rom_addr[0]), .Y(n7121) );
  NAND2X1 U10811 ( .A(B_sel_reg[0]), .B(n11920), .Y(n11931) );
  BUFX3 U10812 ( .A(T1_rom_addr[1]), .Y(n7122) );
  NOR2X4 U10813 ( .A(n7354), .B(n27236), .Y(n11929) );
  INVX1 U10814 ( .A(n28638), .Y(n11885) );
  INVX1 U10815 ( .A(n10236), .Y(n10237) );
  XOR2X1 U10816 ( .A(n10865), .B(n10864), .Y(U1_U2_z0[2]) );
  INVXL U10817 ( .A(n25330), .Y(n6598) );
  INVX1 U10818 ( .A(n10150), .Y(n10151) );
  CLKBUFX8 U10819 ( .A(n16569), .Y(n7127) );
  INVX1 U10820 ( .A(n9920), .Y(n9877) );
  INVX1 U10821 ( .A(n10062), .Y(n10063) );
  INVX1 U10822 ( .A(n10073), .Y(n10074) );
  INVX1 U10823 ( .A(n10078), .Y(n10079) );
  INVX2 U10824 ( .A(n9868), .Y(n6336) );
  NAND2X1 U10825 ( .A(n6402), .B(n9794), .Y(n6401) );
  INVX1 U10826 ( .A(n9976), .Y(n10009) );
  INVX8 U10827 ( .A(n5836), .Y(n15963) );
  XOR2X1 U10828 ( .A(n11206), .B(n11205), .Y(U1_U1_z0[2]) );
  NAND2X1 U10829 ( .A(n11415), .B(n11410), .Y(n11421) );
  NAND2XL U10830 ( .A(n11415), .B(n28708), .Y(n6196) );
  INVXL U10831 ( .A(n7151), .Y(n10628) );
  INVXL U10832 ( .A(n20438), .Y(n6728) );
  INVX1 U10833 ( .A(n11415), .Y(n6206) );
  INVX1 U10834 ( .A(n28643), .Y(n15023) );
  INVX1 U10835 ( .A(n11080), .Y(n11070) );
  AND2X4 U10836 ( .A(buffer[15]), .B(n27236), .Y(n28452) );
  INVX1 U10837 ( .A(n11896), .Y(n28666) );
  INVX1 U10838 ( .A(n10329), .Y(n10330) );
  INVXL U10839 ( .A(n10334), .Y(n10335) );
  AND2X4 U10840 ( .A(buffer[31]), .B(n27236), .Y(n28625) );
  NAND2X1 U10841 ( .A(cnt[9]), .B(n11878), .Y(n14978) );
  NAND2X1 U10842 ( .A(n6826), .B(n10240), .Y(n10243) );
  BUFX3 U10843 ( .A(n10234), .Y(n10235) );
  INVXL U10844 ( .A(n11625), .Y(n7300) );
  NOR2XL U10845 ( .A(U0_U2_y1[13]), .B(n6364), .Y(n7970) );
  OR2XL U10846 ( .A(n11907), .B(n28674), .Y(n7299) );
  NAND2X1 U10847 ( .A(n9795), .B(n9794), .Y(n10084) );
  AND2X2 U10848 ( .A(n9798), .B(n9797), .Y(n10102) );
  CLKINVX8 U10849 ( .A(n5841), .Y(n16128) );
  INVX1 U10850 ( .A(n10292), .Y(n10293) );
  INVX4 U10851 ( .A(n27298), .Y(n5921) );
  AND2X2 U10852 ( .A(n11299), .B(n11298), .Y(n11300) );
  NAND2X1 U10853 ( .A(n9984), .B(n9983), .Y(n10236) );
  NAND2X1 U10854 ( .A(n9788), .B(n9787), .Y(n10055) );
  AND2X2 U10855 ( .A(n10544), .B(n10543), .Y(n10545) );
  AND2X2 U10856 ( .A(n8209), .B(n8317), .Y(n8210) );
  CLKINVX8 U10857 ( .A(n15633), .Y(n16354) );
  AND2XL U10858 ( .A(n13235), .B(U0_U0_y0[13]), .Y(n13236) );
  CLKINVX8 U10859 ( .A(n15495), .Y(n16143) );
  AND2X2 U10860 ( .A(n10589), .B(n10588), .Y(n10590) );
  NAND2X1 U10861 ( .A(n9861), .B(n9860), .Y(n10166) );
  NAND2X1 U10862 ( .A(n9808), .B(n9807), .Y(n10087) );
  AND2X1 U10863 ( .A(n10925), .B(n10924), .Y(n6975) );
  CLKBUFX8 U10864 ( .A(n16277), .Y(n15687) );
  INVX8 U10865 ( .A(n27236), .Y(n5922) );
  NAND2X1 U10866 ( .A(n9912), .B(n9911), .Y(n10322) );
  NAND2X1 U10867 ( .A(n9903), .B(n9902), .Y(n10337) );
  CLKINVX8 U10868 ( .A(n5841), .Y(n16158) );
  NAND2X1 U10869 ( .A(n9776), .B(n9775), .Y(n10048) );
  AND2X2 U10870 ( .A(n11155), .B(n11160), .Y(n11149) );
  NAND2BX1 U10871 ( .AN(out_sel), .B(n15027), .Y(n11654) );
  NAND2X2 U10872 ( .A(n11155), .B(n8284), .Y(n11140) );
  NAND2X1 U10873 ( .A(n11093), .B(n8290), .Y(n6223) );
  NOR2X1 U10874 ( .A(n11873), .B(n7305), .Y(n11896) );
  NAND2X1 U10875 ( .A(n9615), .B(n29104), .Y(n6390) );
  XOR2X2 U10876 ( .A(n8310), .B(n29103), .Y(n6324) );
  NAND2XL U10877 ( .A(cnt[7]), .B(n11633), .Y(n11618) );
  INVX1 U10878 ( .A(n11979), .Y(n14977) );
  NAND2X1 U10879 ( .A(n9990), .B(n9989), .Y(n10238) );
  AOI21X1 U10880 ( .A0(n10289), .A1(n10277), .B0(n7948), .Y(n10278) );
  INVX1 U10881 ( .A(n10289), .Y(n10290) );
  INVX2 U10882 ( .A(n11652), .Y(n14979) );
  NAND2X1 U10883 ( .A(n9909), .B(n9908), .Y(n10319) );
  NAND2X1 U10884 ( .A(n9933), .B(n9932), .Y(n10329) );
  NOR2XL U10885 ( .A(U1_U0_y1[13]), .B(n6654), .Y(n8141) );
  NAND2XL U10886 ( .A(n10458), .B(n10457), .Y(n10459) );
  NAND2X1 U10887 ( .A(n9740), .B(n9753), .Y(n10034) );
  INVX1 U10888 ( .A(n10070), .Y(n10086) );
  NAND2X1 U10889 ( .A(n9771), .B(n9770), .Y(n10078) );
  NAND2X1 U10890 ( .A(n9801), .B(n9800), .Y(n10104) );
  NAND2X1 U10891 ( .A(n10129), .B(n10121), .Y(n10180) );
  INVX1 U10892 ( .A(n11632), .Y(n11878) );
  XOR2X1 U10893 ( .A(n8265), .B(n7256), .Y(n15024) );
  AND2X2 U10894 ( .A(n10483), .B(n10482), .Y(n10484) );
  AND2X2 U10895 ( .A(n10584), .B(n10583), .Y(n10585) );
  AOI21XL U10896 ( .A0(n13734), .A1(n13733), .B0(n13732), .Y(n13742) );
  AND2XL U10897 ( .A(U0_U2_y1[12]), .B(U0_U2_y0[12]), .Y(n8733) );
  AND2XL U10898 ( .A(n11097), .B(n11096), .Y(n11098) );
  AND2X1 U10899 ( .A(n13773), .B(n13759), .Y(n13822) );
  AND2XL U10900 ( .A(n13771), .B(U1_U2_y0[13]), .Y(n7971) );
  INVX1 U10901 ( .A(n10480), .Y(n6329) );
  INVX1 U10902 ( .A(n10231), .Y(n6217) );
  NOR2X1 U10903 ( .A(n10023), .B(n10051), .Y(n10038) );
  NAND2BXL U10904 ( .AN(U1_U2_y0[13]), .B(U1_U2_y2[13]), .Y(n13773) );
  NOR2X1 U10905 ( .A(n29107), .B(n11976), .Y(n11979) );
  INVX1 U10906 ( .A(n9963), .Y(n9965) );
  AND2XL U10907 ( .A(U1_U1_y1[12]), .B(U1_U1_y0[12]), .Y(n14629) );
  INVX1 U10908 ( .A(n9968), .Y(n9970) );
  INVX1 U10909 ( .A(n9972), .Y(n9990) );
  AND2XL U10910 ( .A(n14170), .B(U0_U0_y0[13]), .Y(n8049) );
  INVX1 U10911 ( .A(n10994), .Y(n10987) );
  AND2XL U10912 ( .A(U1_U2_y2[12]), .B(U1_U2_y0[12]), .Y(n13772) );
  OR2X1 U10913 ( .A(n25330), .B(U0_pipe11[27]), .Y(n7754) );
  INVX1 U10914 ( .A(n11989), .Y(n29241) );
  INVX1 U10915 ( .A(n10241), .Y(n6827) );
  INVX1 U10916 ( .A(n9961), .Y(n9981) );
  INVX1 U10917 ( .A(n9820), .Y(n9822) );
  NAND2X1 U10918 ( .A(n11418), .B(BOPA[12]), .Y(n9620) );
  INVX1 U10919 ( .A(n14996), .Y(n11655) );
  BUFX4 U10920 ( .A(n25330), .Y(n20025) );
  INVX1 U10921 ( .A(n10224), .Y(n10225) );
  INVXL U10922 ( .A(U1_U2_y2[13]), .Y(n13771) );
  NAND2BX1 U10923 ( .AN(n7986), .B(n8000), .Y(n6180) );
  INVXL U10924 ( .A(U0_U0_y1[13]), .Y(n13235) );
  AND2XL U10925 ( .A(U0_U0_y1[12]), .B(U0_U0_y0[12]), .Y(n13237) );
  INVX1 U10926 ( .A(n10134), .Y(n10135) );
  INVX1 U10927 ( .A(n9842), .Y(n9838) );
  INVX1 U10928 ( .A(n9980), .Y(n9962) );
  INVX1 U10929 ( .A(n9989), .Y(n9973) );
  INVX4 U10930 ( .A(n7305), .Y(n11633) );
  INVX1 U10931 ( .A(n9837), .Y(n9843) );
  INVXL U10932 ( .A(n13745), .Y(n13752) );
  INVX1 U10933 ( .A(n9774), .Y(n9776) );
  AND2XL U10934 ( .A(U1_U0_y1[12]), .B(U1_U0_y0[12]), .Y(n9285) );
  NAND2X1 U10935 ( .A(n11418), .B(BOPA[21]), .Y(n11413) );
  INVX1 U10936 ( .A(n10512), .Y(n10349) );
  AND2XL U10937 ( .A(U0_U1_y1[12]), .B(U0_U1_y0[12]), .Y(n8793) );
  AND2XL U10938 ( .A(U1_U2_y1[12]), .B(U1_U2_y0[12]), .Y(n12748) );
  INVX1 U10939 ( .A(n9932), .Y(n9891) );
  AND2XL U10940 ( .A(U0_U2_y2[12]), .B(U0_U2_y0[12]), .Y(n12051) );
  NOR2X1 U10941 ( .A(n10370), .B(n10376), .Y(n10355) );
  INVX1 U10942 ( .A(n9905), .Y(n9912) );
  INVXL U10943 ( .A(n10559), .Y(n10561) );
  CLKINVX3 U10944 ( .A(n9916), .Y(n6162) );
  AND2X2 U10945 ( .A(n11410), .B(n28710), .Y(n6272) );
  CLKINVX2 U10946 ( .A(n7388), .Y(n10776) );
  INVX1 U10947 ( .A(n9886), .Y(n9888) );
  NAND2X1 U10948 ( .A(n11613), .B(n28706), .Y(n11873) );
  INVX1 U10949 ( .A(n9780), .Y(n9782) );
  INVX1 U10950 ( .A(n9890), .Y(n9933) );
  INVX1 U10951 ( .A(n9897), .Y(n9899) );
  INVX1 U10952 ( .A(n9892), .Y(n9894) );
  INVXL U10953 ( .A(n10359), .Y(n8229) );
  INVX1 U10954 ( .A(n10256), .Y(n10259) );
  INVX1 U10955 ( .A(n10257), .Y(n10258) );
  OAI21X2 U10956 ( .A0(n10200), .A1(n10224), .B0(n10199), .Y(n10216) );
  INVXL U10957 ( .A(n11024), .Y(n10876) );
  INVXL U10958 ( .A(n10808), .Y(n10810) );
  INVX1 U10959 ( .A(n11991), .Y(n11994) );
  INVXL U10960 ( .A(n13736), .Y(n13739) );
  NAND2X1 U10961 ( .A(W3[7]), .B(W3[23]), .Y(n9749) );
  NAND2BX1 U10962 ( .AN(ram_sel_reg[9]), .B(n28759), .Y(n14994) );
  NAND2X1 U10963 ( .A(n28677), .B(n28671), .Y(n16245) );
  NAND2X1 U10964 ( .A(n8191), .B(BOPC[36]), .Y(n11159) );
  NAND2X1 U10965 ( .A(n28758), .B(n29107), .Y(n11949) );
  NOR2X1 U10966 ( .A(BOPC[25]), .B(n8130), .Y(n11211) );
  NAND2X1 U10967 ( .A(n7052), .B(BOPC[42]), .Y(n11105) );
  NOR2X1 U10968 ( .A(n7059), .B(BOPC[44]), .Y(n11083) );
  NAND2X1 U10969 ( .A(n7059), .B(BOPC[44]), .Y(n11096) );
  AND2XL U10970 ( .A(U0_U0_y1[3]), .B(U0_U0_y0[3]), .Y(n13198) );
  OR2XL U10971 ( .A(U0_U0_y1[3]), .B(U0_U0_y0[3]), .Y(n13200) );
  NOR2X1 U10972 ( .A(cnt[9]), .B(n29107), .Y(n11613) );
  INVX1 U10973 ( .A(B1_q[42]), .Y(n16398) );
  XOR2X1 U10974 ( .A(n7959), .B(n7976), .Y(n7407) );
  AND2XL U10975 ( .A(U0_U0_y1[9]), .B(U0_U0_y0[9]), .Y(n13228) );
  AND2XL U10976 ( .A(U0_U0_y1[5]), .B(U0_U0_y0[5]), .Y(n13208) );
  NAND2X1 U10977 ( .A(n29106), .B(BOPA[0]), .Y(n7302) );
  INVX1 U10978 ( .A(B1_q[32]), .Y(n16439) );
  INVX1 U10979 ( .A(B1_q[34]), .Y(n16431) );
  AND2XL U10980 ( .A(U1_U1_y2[7]), .B(U1_U1_y0[7]), .Y(n12671) );
  OR2XL U10981 ( .A(U1_U1_y2[12]), .B(U1_U1_y0[12]), .Y(n12679) );
  AND2XL U10982 ( .A(U1_U1_y2[12]), .B(U1_U1_y0[12]), .Y(n12690) );
  INVX1 U10983 ( .A(B5_q[40]), .Y(n15819) );
  INVX1 U10984 ( .A(B5_q[30]), .Y(n15859) );
  INVX1 U10985 ( .A(B1_q[11]), .Y(n16527) );
  INVX1 U10986 ( .A(B1_q[1]), .Y(n16567) );
  XOR2X1 U10987 ( .A(n7986), .B(W3[15]), .Y(n6181) );
  INVX1 U10988 ( .A(B1_q[40]), .Y(n16406) );
  AND2XL U10989 ( .A(U1_U2_y2[11]), .B(U1_U2_y0[11]), .Y(n13767) );
  AND2XL U10990 ( .A(U1_U2_y1[1]), .B(U1_U2_y0[1]), .Y(n8142) );
  AND2XL U10991 ( .A(U1_U2_y1[2]), .B(U1_U2_y0[2]), .Y(n12713) );
  AND2XL U10992 ( .A(U1_U2_y1[3]), .B(U1_U2_y0[3]), .Y(n12712) );
  OR2XL U10993 ( .A(U1_U2_y1[5]), .B(U1_U2_y0[5]), .Y(n12723) );
  AND2XL U10994 ( .A(U1_U2_y1[4]), .B(U1_U2_y0[4]), .Y(n12722) );
  AND2XL U10995 ( .A(U1_U2_y1[5]), .B(U1_U2_y0[5]), .Y(n12721) );
  AND2XL U10996 ( .A(U1_U2_y1[6]), .B(U1_U2_y0[6]), .Y(n12725) );
  AND2XL U10997 ( .A(U1_U2_y1[7]), .B(U1_U2_y0[7]), .Y(n12724) );
  AND2XL U10998 ( .A(U0_U1_y2[12]), .B(U0_U1_y0[12]), .Y(n12447) );
  OR2XL U10999 ( .A(U1_U2_y1[8]), .B(U1_U2_y0[8]), .Y(n12734) );
  INVX1 U11000 ( .A(B1_q[30]), .Y(n16447) );
  AND2XL U11001 ( .A(U0_U1_y2[7]), .B(U0_U1_y0[7]), .Y(n12424) );
  AND2XL U11002 ( .A(U1_U2_y1[11]), .B(U1_U2_y0[11]), .Y(n12740) );
  NOR2X1 U11003 ( .A(BOPA[47]), .B(BOPA[46]), .Y(n11410) );
  AND2XL U11004 ( .A(U1_U0_y2[9]), .B(U1_U0_y0[9]), .Y(n8389) );
  OR2X1 U11005 ( .A(U1_U2_y2[5]), .B(U1_U2_y0[5]), .Y(n13743) );
  AND2XL U11006 ( .A(U1_U2_y2[1]), .B(U1_U2_y0[1]), .Y(n13732) );
  AND2XL U11007 ( .A(U1_U0_y2[5]), .B(U1_U0_y0[5]), .Y(n8374) );
  NOR2X1 U11008 ( .A(n6908), .B(W3[17]), .Y(n10011) );
  AND2XL U11009 ( .A(U0_U2_y2[5]), .B(U0_U2_y0[5]), .Y(n12024) );
  AND2XL U11010 ( .A(n7982), .B(W3[30]), .Y(n7983) );
  AND2XL U11011 ( .A(U0_U2_y2[7]), .B(U0_U2_y0[7]), .Y(n12027) );
  OR2XL U11012 ( .A(U0_U2_y2[8]), .B(U0_U2_y0[8]), .Y(n12038) );
  NOR2X1 U11013 ( .A(n8094), .B(AOPD[48]), .Y(n10900) );
  AND2XL U11014 ( .A(U0_U0_y2[12]), .B(U0_U0_y0[12]), .Y(n14171) );
  NAND2X1 U11015 ( .A(W0[11]), .B(W0[27]), .Y(n9827) );
  AND2XL U11016 ( .A(U0_U0_y2[9]), .B(U0_U0_y0[9]), .Y(n14162) );
  NAND2X1 U11017 ( .A(n6908), .B(W3[17]), .Y(n10010) );
  AND2XL U11018 ( .A(U0_U2_y2[3]), .B(U0_U2_y0[3]), .Y(n12013) );
  OR2XL U11019 ( .A(U0_U1_y1[8]), .B(U0_U1_y0[8]), .Y(n8780) );
  NAND2X1 U11020 ( .A(W3[5]), .B(W3[21]), .Y(n9781) );
  INVX1 U11021 ( .A(B1_q[7]), .Y(n16543) );
  NOR2X1 U11022 ( .A(BOPD[25]), .B(n8131), .Y(n10850) );
  NAND2X1 U11023 ( .A(n7955), .B(AOPB[38]), .Y(n10448) );
  NOR2X1 U11024 ( .A(n8045), .B(W3[25]), .Y(n10023) );
  NOR2X1 U11025 ( .A(W3[12]), .B(W3[28]), .Y(n9803) );
  OR2XL U11026 ( .A(U0_U1_y1[5]), .B(U0_U1_y0[5]), .Y(n8768) );
  OR2XL U11027 ( .A(U0_U1_y1[6]), .B(U0_U1_y0[6]), .Y(n8764) );
  AND2XL U11028 ( .A(U0_U1_y1[7]), .B(U0_U1_y0[7]), .Y(n8769) );
  NOR2X1 U11029 ( .A(W2[15]), .B(n7978), .Y(n10326) );
  NAND2X1 U11030 ( .A(n8031), .B(W2[29]), .Y(n10275) );
  AND2XL U11031 ( .A(U1_U1_y1[1]), .B(U1_U1_y0[1]), .Y(n14584) );
  AND2XL U11032 ( .A(n8012), .B(W2[30]), .Y(n7948) );
  INVX1 U11033 ( .A(B5_q[3]), .Y(n15972) );
  INVX2 U11034 ( .A(n25330), .Y(n5928) );
  BUFX1 U11035 ( .A(U2_A_r_d[14]), .Y(n6730) );
  NAND2X1 U11036 ( .A(n8050), .B(W1[25]), .Y(n10199) );
  INVXL U11037 ( .A(U2_A_r_d[14]), .Y(n6227) );
  AND2XL U11038 ( .A(U0_U0_y2[3]), .B(U0_U0_y0[3]), .Y(n14184) );
  AND2XL U11039 ( .A(U1_U1_y1[7]), .B(U1_U1_y0[7]), .Y(n14604) );
  INVX1 U11040 ( .A(B5_q[41]), .Y(n15815) );
  INVX1 U11041 ( .A(B5_q[33]), .Y(n15847) );
  AND2XL U11042 ( .A(U0_U0_y2[6]), .B(U0_U0_y0[6]), .Y(n14198) );
  AND2XL U11043 ( .A(U1_U1_y1[5]), .B(U1_U1_y0[5]), .Y(n14601) );
  NAND2X1 U11044 ( .A(n8042), .B(W2[23]), .Y(n10268) );
  AND2XL U11045 ( .A(U0_U0_y2[5]), .B(U0_U0_y0[5]), .Y(n14194) );
  AND2XL U11046 ( .A(U1_U1_y1[6]), .B(U1_U1_y0[6]), .Y(n14605) );
  INVX1 U11047 ( .A(B5_q[31]), .Y(n15855) );
  NAND2X1 U11048 ( .A(n28672), .B(D_sel_reg_4__0_), .Y(n15218) );
  NOR2X1 U11049 ( .A(D_sel_reg_4__0_), .B(n28672), .Y(n15214) );
  NAND2X1 U11050 ( .A(ram_sel_reg[9]), .B(n28759), .Y(n14998) );
  INVX4 U11051 ( .A(n15967), .Y(n5930) );
  NAND2X1 U11052 ( .A(cnt[9]), .B(cnt[8]), .Y(n11976) );
  CLKINVX3 U11053 ( .A(n16163), .Y(n5931) );
  INVX1 U11054 ( .A(B5_q[51]), .Y(n15775) );
  INVX1 U11055 ( .A(B1_q[5]), .Y(n16550) );
  NAND2X1 U11056 ( .A(cnt[0]), .B(cnt[2]), .Y(n11963) );
  AND2XL U11057 ( .A(U1_U0_y1[6]), .B(U1_U0_y0[6]), .Y(n9261) );
  NAND2X1 U11058 ( .A(ram_sel_reg[9]), .B(ram_sel_reg[8]), .Y(n14993) );
  AND2XL U11059 ( .A(U1_U0_y1[5]), .B(U1_U0_y0[5]), .Y(n9257) );
  INVX4 U11060 ( .A(n16154), .Y(n5933) );
  INVXL U11061 ( .A(U1_A_r_d0[10]), .Y(n6515) );
  INVX1 U11062 ( .A(B5_q[24]), .Y(n15883) );
  NOR2X2 U11063 ( .A(n8113), .B(AOPB[43]), .Y(n10404) );
  INVX1 U11064 ( .A(in_valid), .Y(n29099) );
  NAND2X1 U11065 ( .A(n13898), .B(n13899), .Y(n13910) );
  NOR2X2 U11066 ( .A(n13898), .B(n13899), .Y(n13909) );
  XOR2X2 U11067 ( .A(n5939), .B(n13933), .Y(n20014) );
  NAND3X1 U11068 ( .A(n20056), .B(n20101), .C(n7870), .Y(n7865) );
  AOI21X2 U11069 ( .A0(n13873), .A1(n13860), .B0(n13855), .Y(n5945) );
  NAND3X2 U11070 ( .A(n5947), .B(n7817), .C(n5946), .Y(n12970) );
  NAND3BX2 U11071 ( .AN(n12959), .B(n12957), .C(n7816), .Y(n5947) );
  NAND2X1 U11072 ( .A(n13553), .B(n17372), .Y(n5950) );
  OAI21X2 U11073 ( .A0(n5951), .A1(n13039), .B0(n13043), .Y(n6107) );
  XOR2X2 U11074 ( .A(n5951), .B(n13014), .Y(n19544) );
  AOI21X2 U11075 ( .A0(n6100), .A1(n7876), .B0(n7269), .Y(n7446) );
  NAND2X2 U11076 ( .A(n5954), .B(n5952), .Y(n6100) );
  NOR2X1 U11077 ( .A(n19579), .B(n19562), .Y(n5953) );
  NOR2X1 U11078 ( .A(n7270), .B(n19559), .Y(n19579) );
  NAND2X2 U11079 ( .A(n6101), .B(n6869), .Y(n19578) );
  OAI21X1 U11080 ( .A0(n5955), .A1(n17328), .B0(n17334), .Y(n17332) );
  XOR2X1 U11081 ( .A(n5955), .B(n17336), .Y(n17337) );
  NOR2X2 U11082 ( .A(n12952), .B(n12953), .Y(n12996) );
  NOR2X1 U11083 ( .A(n7873), .B(n7799), .Y(n6097) );
  AOI21X2 U11084 ( .A0(n7157), .A1(n7842), .B0(n20328), .Y(n7799) );
  NAND3BX4 U11085 ( .AN(n6680), .B(n5956), .C(n20315), .Y(n7157) );
  OAI21X4 U11086 ( .A0(n6055), .A1(n20319), .B0(n20318), .Y(n5956) );
  XOR2X4 U11087 ( .A(n7899), .B(n13937), .Y(n19998) );
  NAND2X4 U11088 ( .A(n7146), .B(n13960), .Y(n7200) );
  NOR2X4 U11089 ( .A(n13920), .B(n7871), .Y(n13960) );
  NAND3X2 U11090 ( .A(n6050), .B(n6049), .C(n13852), .Y(n7841) );
  NAND2X2 U11091 ( .A(n5970), .B(n6049), .Y(n7840) );
  NAND2BX2 U11092 ( .AN(n13888), .B(n5960), .Y(n5966) );
  NOR2X1 U11093 ( .A(n14008), .B(n13948), .Y(n5965) );
  AOI21X2 U11094 ( .A0(n5968), .A1(n6156), .B0(n5967), .Y(n17056) );
  OAI21X1 U11095 ( .A0(n17058), .A1(n16796), .B0(n16797), .Y(n5967) );
  XOR2X2 U11096 ( .A(n13908), .B(n13907), .Y(n14945) );
  INVX1 U11097 ( .A(n7867), .Y(n5970) );
  NAND4X2 U11098 ( .A(n6167), .B(n6168), .C(n7456), .D(n6710), .Y(n7470) );
  NOR2X1 U11099 ( .A(n5974), .B(n14924), .Y(n5982) );
  OR2X2 U11100 ( .A(n16872), .B(n14937), .Y(n5978) );
  AOI22X1 U11101 ( .A0(n6952), .A1(n14942), .B0(n19987), .B1(n14941), .Y(n5979) );
  INVX2 U11102 ( .A(n12970), .Y(n14941) );
  NOR2XL U11103 ( .A(n14943), .B(n16859), .Y(n5981) );
  NAND2X1 U11104 ( .A(n14939), .B(n14928), .Y(n16859) );
  NOR2XL U11105 ( .A(n14933), .B(n14934), .Y(n16871) );
  OAI21X2 U11106 ( .A0(n13808), .A1(n13813), .B0(n13809), .Y(n5983) );
  NAND2X1 U11107 ( .A(n13782), .B(n13781), .Y(n13809) );
  AOI21X1 U11108 ( .A0(n6100), .A1(n7881), .B0(n7906), .Y(n5984) );
  AOI21X4 U11109 ( .A0(n14850), .A1(n14681), .B0(n14684), .Y(n14862) );
  OAI21X4 U11110 ( .A0(n14848), .A1(n14846), .B0(n14847), .Y(n14850) );
  NAND2X4 U11111 ( .A(n5987), .B(n6124), .Y(n14848) );
  NAND2X4 U11112 ( .A(n7815), .B(n5988), .Y(n6130) );
  AOI21X2 U11113 ( .A0(n5988), .A1(n14775), .B0(n14774), .Y(n7420) );
  XOR2X1 U11114 ( .A(n5988), .B(n14765), .Y(n19978) );
  NAND4X4 U11115 ( .A(n6695), .B(n7307), .C(n7308), .D(n6693), .Y(n5988) );
  NAND2X2 U11116 ( .A(n6725), .B(n6722), .Y(n13983) );
  OAI21X4 U11117 ( .A0(n7721), .A1(n7871), .B0(n7154), .Y(n6048) );
  AND2X2 U11118 ( .A(n7814), .B(n7863), .Y(n6004) );
  AOI21X2 U11119 ( .A0(n19240), .A1(n14855), .B0(n5994), .Y(n19235) );
  XOR2X1 U11120 ( .A(n5995), .B(n7033), .Y(n19238) );
  AOI21X1 U11121 ( .A0(n19234), .A1(n5997), .B0(n5996), .Y(n5995) );
  INVXL U11122 ( .A(n19236), .Y(n5997) );
  OAI21X4 U11123 ( .A0(n19267), .A1(n7040), .B0(n7895), .Y(n19234) );
  XOR2X4 U11124 ( .A(n7874), .B(n13055), .Y(n7915) );
  XOR2X4 U11125 ( .A(n6137), .B(n5790), .Y(n20011) );
  NOR2X2 U11126 ( .A(n13004), .B(n13005), .Y(n13039) );
  INVX1 U11127 ( .A(n13854), .Y(n6056) );
  INVXL U11128 ( .A(n14944), .Y(n16838) );
  AOI21X1 U11129 ( .A0(n16809), .A1(n16855), .B0(n16808), .Y(n16823) );
  AOI21X1 U11130 ( .A0(n13954), .A1(n13955), .B0(n7473), .Y(n6000) );
  AOI2BB1X2 U11131 ( .A0N(n17056), .A1N(n7510), .B0(n7507), .Y(n6045) );
  NOR2X2 U11132 ( .A(n14648), .B(n14649), .Y(n14769) );
  OAI21X1 U11133 ( .A0(n19267), .A1(n19257), .B0(n19256), .Y(n19265) );
  AOI21X4 U11134 ( .A0(n19299), .A1(n7204), .B0(n7203), .Y(n19267) );
  NAND2X1 U11135 ( .A(n20007), .B(n5866), .Y(n14830) );
  AOI21X1 U11136 ( .A0(n12781), .A1(n12890), .B0(n12893), .Y(n12921) );
  NAND2X1 U11137 ( .A(n12796), .B(n7468), .Y(n12891) );
  NOR2X1 U11138 ( .A(n12697), .B(n12696), .Y(n12866) );
  NAND2X2 U11139 ( .A(n6009), .B(n14808), .Y(n7888) );
  NAND2X1 U11140 ( .A(n6009), .B(n14807), .Y(n6008) );
  NOR2X2 U11141 ( .A(n14809), .B(n14812), .Y(n6009) );
  AOI21X2 U11142 ( .A0(n6010), .A1(n7898), .B0(n7897), .Y(n6137) );
  AOI21X2 U11143 ( .A0(n20055), .A1(n7870), .B0(n6011), .Y(n6083) );
  OAI21X1 U11144 ( .A0(n20057), .A1(n6016), .B0(n6012), .Y(n6011) );
  NOR2X2 U11145 ( .A(n6015), .B(n6014), .Y(n20057) );
  AND2X2 U11146 ( .A(n20012), .B(n6901), .Y(n6015) );
  NOR2X1 U11147 ( .A(n6016), .B(n20058), .Y(n7870) );
  OAI21X2 U11148 ( .A0(n20080), .A1(n20010), .B0(n6017), .Y(n20055) );
  NOR2X2 U11149 ( .A(n20004), .B(n6018), .Y(n20080) );
  AOI21X1 U11150 ( .A0(n7866), .A1(n6022), .B0(n6021), .Y(n6020) );
  XOR2X2 U11151 ( .A(n6023), .B(n6905), .Y(n19994) );
  NOR2X1 U11152 ( .A(n7721), .B(n13913), .Y(n6025) );
  NAND3BX2 U11153 ( .AN(n13920), .B(n7841), .C(n7840), .Y(n6051) );
  NAND2X2 U11154 ( .A(n13891), .B(n13896), .Y(n13920) );
  OAI21X2 U11155 ( .A0(n13872), .A1(n13871), .B0(n13870), .Y(n13895) );
  NAND2X1 U11156 ( .A(n13853), .B(n13854), .Y(n13871) );
  XOR2X2 U11157 ( .A(U1_U2_y2[23]), .B(U1_U2_y0[23]), .Y(n13853) );
  NOR2X2 U11158 ( .A(n6028), .B(n6027), .Y(n6026) );
  NAND2XL U11159 ( .A(n12701), .B(n12700), .Y(n12803) );
  NOR2X4 U11160 ( .A(n12700), .B(n12701), .Y(n12802) );
  NAND2X1 U11161 ( .A(n6031), .B(n17666), .Y(n6030) );
  XOR2X4 U11162 ( .A(n13917), .B(n13916), .Y(n20002) );
  NAND2X1 U11163 ( .A(n13850), .B(n13849), .Y(n13866) );
  NAND2X1 U11164 ( .A(n13798), .B(n13797), .Y(n13862) );
  OAI21X2 U11165 ( .A0(n13795), .A1(n13794), .B0(n13793), .Y(n7469) );
  NOR2X2 U11166 ( .A(n13786), .B(n13785), .Y(n13795) );
  NOR2X2 U11167 ( .A(n13798), .B(n13797), .Y(n13863) );
  XOR2X2 U11168 ( .A(n13880), .B(n13879), .Y(n14930) );
  NAND2X4 U11169 ( .A(n13057), .B(n7927), .Y(n7788) );
  NOR2X2 U11170 ( .A(n13016), .B(n13026), .Y(n13057) );
  NOR2X2 U11171 ( .A(n12982), .B(n12983), .Y(n13026) );
  INVXL U11172 ( .A(n14503), .Y(n6038) );
  AOI21X1 U11173 ( .A0(n17633), .A1(n13070), .B0(n7967), .Y(n14504) );
  NOR2X2 U11174 ( .A(n6041), .B(n14499), .Y(n6040) );
  NAND2X1 U11175 ( .A(n17628), .B(n14503), .Y(n6041) );
  XOR2X2 U11176 ( .A(n7919), .B(n6927), .Y(n14959) );
  XOR2X4 U11177 ( .A(n7836), .B(n6978), .Y(n14948) );
  NAND3X2 U11178 ( .A(n7917), .B(n7918), .C(n7920), .Y(n14960) );
  NAND2BX2 U11179 ( .AN(n19996), .B(n5856), .Y(n16819) );
  NOR2X1 U11180 ( .A(n17074), .B(n6062), .Y(n6047) );
  AOI21X4 U11181 ( .A0(n13895), .A1(n13896), .B0(n7477), .Y(n7721) );
  AOI21X2 U11182 ( .A0(n20361), .A1(n14889), .B0(n14888), .Y(n20353) );
  OAI21X2 U11183 ( .A0(n14887), .A1(n20364), .B0(n14886), .Y(n20319) );
  NOR2BX2 U11184 ( .AN(n20310), .B(n20320), .Y(n6055) );
  NOR2BX2 U11185 ( .AN(n13860), .B(n13872), .Y(n13891) );
  XOR2X4 U11186 ( .A(n6057), .B(n6920), .Y(n14929) );
  AOI21X2 U11187 ( .A0(n13873), .A1(n13891), .B0(n13895), .Y(n13880) );
  NOR2X1 U11188 ( .A(n19998), .B(n14957), .Y(n6062) );
  OAI21X4 U11189 ( .A0(n13837), .A1(n13835), .B0(n13838), .Y(n13803) );
  NAND2X1 U11190 ( .A(n13777), .B(n13778), .Y(n13838) );
  NAND2X2 U11191 ( .A(n6071), .B(n13802), .Y(n13848) );
  NAND2X1 U11192 ( .A(n14927), .B(n14932), .Y(n17117) );
  NOR2X2 U11193 ( .A(n12783), .B(n12782), .Y(n12920) );
  NOR2BX2 U11194 ( .AN(n7830), .B(n6075), .Y(n6074) );
  OAI21X4 U11195 ( .A0(n6703), .A1(n7826), .B0(n7929), .Y(n7830) );
  NOR2X2 U11196 ( .A(n13894), .B(n13890), .Y(n13896) );
  NOR2X2 U11197 ( .A(n7839), .B(n13876), .Y(n13894) );
  NOR2X1 U11198 ( .A(n20006), .B(n14953), .Y(n16836) );
  AOI21X1 U11199 ( .A0(n7188), .A1(n7866), .B0(n7187), .Y(n6082) );
  NAND2X4 U11200 ( .A(n7865), .B(n6083), .Y(n7866) );
  NAND2X2 U11201 ( .A(n7867), .B(n7869), .Y(n6085) );
  NOR2X1 U11202 ( .A(n5845), .B(n14966), .Y(n16796) );
  AOI21X2 U11203 ( .A0(n13639), .A1(n13628), .B0(n13638), .Y(n13654) );
  AND2X2 U11204 ( .A(U1_U1_y0[32]), .B(U1_U1_y2[32]), .Y(n13084) );
  AOI21X4 U11205 ( .A0(n13609), .A1(n13595), .B0(n13608), .Y(n13627) );
  NAND2X4 U11206 ( .A(n6091), .B(n6087), .Y(n13609) );
  AOI21X4 U11207 ( .A0(n6089), .A1(n5884), .B0(n6088), .Y(n6087) );
  NAND2X1 U11208 ( .A(n13584), .B(n13583), .Y(n6090) );
  OAI21X2 U11209 ( .A0(n7940), .A1(n13593), .B0(n6092), .Y(n6091) );
  NOR2X1 U11210 ( .A(n13588), .B(n13591), .Y(n6092) );
  OAI21X2 U11211 ( .A0(n20030), .A1(n20022), .B0(n20021), .Y(n7187) );
  NOR2X2 U11212 ( .A(n6093), .B(n7960), .Y(n20030) );
  NAND2XL U11213 ( .A(n7489), .B(n6097), .Y(n6095) );
  OAI21XL U11214 ( .A0(n6098), .A1(n6097), .B0(n7490), .Y(n6096) );
  AOI21X2 U11215 ( .A0(n7463), .A1(n13908), .B0(n7460), .Y(n7459) );
  AOI21X1 U11216 ( .A0(n6099), .A1(n6719), .B0(n6718), .Y(n6717) );
  XOR2X1 U11217 ( .A(n7033), .B(n6100), .Y(n19577) );
  OAI21X2 U11218 ( .A0(n6103), .A1(n19594), .B0(n6102), .Y(n6101) );
  NOR2X4 U11219 ( .A(n19593), .B(n7804), .Y(n6103) );
  NOR2X4 U11220 ( .A(n6111), .B(n19536), .Y(n19593) );
  NAND2X1 U11221 ( .A(n14671), .B(n14670), .Y(n7159) );
  AND2X2 U11222 ( .A(U1_U1_y0[32]), .B(U1_U1_y1[32]), .Y(n14671) );
  NAND2BX1 U11223 ( .AN(n7807), .B(n6106), .Y(n6105) );
  AOI21XL U11224 ( .A0(n7886), .A1(n5882), .B0(n7802), .Y(n6106) );
  XOR2X4 U11225 ( .A(n6107), .B(n6977), .Y(n19282) );
  XOR2X4 U11226 ( .A(n6108), .B(n6968), .Y(n20007) );
  AOI21X1 U11227 ( .A0(n19548), .A1(n19547), .B0(n19546), .Y(n6109) );
  OAI21XL U11228 ( .A0(n7856), .A1(n6117), .B0(n6116), .Y(n6115) );
  INVXL U11229 ( .A(n7855), .Y(n6117) );
  NAND2BX1 U11230 ( .AN(n20040), .B(n7866), .Y(n6119) );
  MXI2X1 U11231 ( .A(n6121), .B(U1_pipe3[26]), .S0(n6120), .Y(n5066) );
  NOR2X2 U11232 ( .A(n14669), .B(n14668), .Y(n14801) );
  XOR2X4 U11233 ( .A(n14850), .B(n6966), .Y(n20033) );
  NOR2X1 U11234 ( .A(n20031), .B(n20022), .Y(n7188) );
  NOR2X1 U11235 ( .A(n20033), .B(n20020), .Y(n20022) );
  NOR2X2 U11236 ( .A(n14801), .B(n14804), .Y(n7894) );
  AOI21X4 U11237 ( .A0(n6127), .A1(n7866), .B0(n20024), .Y(n6126) );
  XOR2X4 U11238 ( .A(n6129), .B(n7189), .Y(n14852) );
  AND2X2 U11239 ( .A(n7370), .B(n7371), .Y(n6129) );
  NOR2X2 U11240 ( .A(n14662), .B(n14663), .Y(n14812) );
  NOR2X2 U11241 ( .A(n14664), .B(n14665), .Y(n14809) );
  NAND2BX4 U11242 ( .AN(n6130), .B(n5882), .Y(n7803) );
  AND2X2 U11243 ( .A(U1_U1_y1[25]), .B(U1_U1_y0[25]), .Y(n7044) );
  INVX1 U11244 ( .A(n14777), .Y(n6132) );
  NOR2X1 U11245 ( .A(n14809), .B(n14813), .Y(n6134) );
  NAND2X1 U11246 ( .A(n14663), .B(n14662), .Y(n14813) );
  OAI21X2 U11247 ( .A0(n14817), .A1(n14821), .B0(n14818), .Y(n14807) );
  NAND2X2 U11248 ( .A(n14659), .B(n14658), .Y(n14821) );
  INVX1 U11249 ( .A(n22930), .Y(n22949) );
  MXI2X1 U11250 ( .A(U0_pipe11[22]), .B(n22994), .S0(n22853), .Y(n4527) );
  NAND2X1 U11251 ( .A(n13531), .B(n24860), .Y(n13532) );
  OAI21X1 U11252 ( .A0(n18356), .A1(n18355), .B0(n18354), .Y(n18488) );
  OAI21X1 U11253 ( .A0(n18766), .A1(n18765), .B0(n18808), .Y(n18772) );
  BUFX3 U11254 ( .A(n11172), .Y(n11141) );
  OAI21XL U11255 ( .A0(n18492), .A1(n18491), .B0(n18490), .Y(n18493) );
  NOR2X2 U11256 ( .A(n8194), .B(BOPC[26]), .Y(n7293) );
  AOI21X2 U11257 ( .A0(n13476), .A1(n13285), .B0(n13288), .Y(n13481) );
  AOI21X1 U11258 ( .A0(n13282), .A1(n13430), .B0(n13281), .Y(n13467) );
  AOI21X1 U11259 ( .A0(n13485), .A1(n13291), .B0(n13294), .Y(n13498) );
  AOI21X2 U11260 ( .A0(n12175), .A1(n6762), .B0(n12174), .Y(n25677) );
  OAI21XL U11261 ( .A0(n8820), .A1(n8830), .B0(n8832), .Y(n8816) );
  NOR2X1 U11262 ( .A(n24582), .B(n13107), .Y(n25764) );
  AOI21X1 U11263 ( .A0(n25756), .A1(n12087), .B0(n12130), .Y(n12131) );
  NOR2X1 U11264 ( .A(n8879), .B(n8884), .Y(n8797) );
  INVX1 U11265 ( .A(n8938), .Y(n8909) );
  XNOR2X2 U11266 ( .A(n9732), .B(n9731), .Y(U1_U1_z2[14]) );
  NOR2X2 U11267 ( .A(n8070), .B(AOPC[31]), .Y(n11364) );
  AOI21X1 U11268 ( .A0(n11607), .A1(n11605), .B0(n11496), .Y(n11501) );
  OR2X2 U11269 ( .A(n11438), .B(U2_B_r[14]), .Y(n11540) );
  AOI21XL U11270 ( .A0(n10274), .A1(n10298), .B0(n10273), .Y(n10285) );
  OAI21X2 U11271 ( .A0(n6224), .A1(n11427), .B0(n9240), .Y(U2_B_i[14]) );
  AOI21X4 U11272 ( .A0(n13616), .A1(n13604), .B0(n13615), .Y(n13633) );
  NOR2X4 U11273 ( .A(n14223), .B(n14222), .Y(n14359) );
  XOR2X1 U11274 ( .A(U1_U2_y1[33]), .B(U1_U2_y0[33]), .Y(n7882) );
  INVX1 U11275 ( .A(n25188), .Y(n25497) );
  CLKINVX3 U11276 ( .A(n7861), .Y(n19568) );
  NOR2X1 U11277 ( .A(n13564), .B(n13568), .Y(n13570) );
  NOR2X1 U11278 ( .A(n13602), .B(n13601), .Y(n6139) );
  XNOR2X2 U11279 ( .A(n10408), .B(n10407), .Y(U0_U0_z0[17]) );
  XNOR2X2 U11280 ( .A(n8289), .B(n6955), .Y(U1_U1_z0[16]) );
  OAI21X2 U11281 ( .A0(n11150), .A1(n11159), .B0(n11151), .Y(n8283) );
  AOI21X1 U11282 ( .A0(n25592), .A1(n25552), .B0(n25551), .Y(n25567) );
  OAI21X1 U11283 ( .A0(n14330), .A1(n14276), .B0(n14275), .Y(n14289) );
  NOR2X2 U11284 ( .A(n8072), .B(AOPB[31]), .Y(n10492) );
  OAI21XL U11285 ( .A0(n25563), .A1(n25558), .B0(n25557), .Y(n25560) );
  OAI21XL U11286 ( .A0(n14286), .A1(n14282), .B0(n14283), .Y(n14281) );
  MXI2X1 U11287 ( .A(U0_pipe8[20]), .B(n25561), .S0(n25611), .Y(n4414) );
  NOR2XL U11288 ( .A(n25251), .B(U2_A_r_d[6]), .Y(n25468) );
  NOR2X1 U11289 ( .A(n14173), .B(U0_U0_y2[13]), .Y(n14317) );
  OAI21X1 U11290 ( .A0(n14801), .A1(n14805), .B0(n14802), .Y(n14793) );
  AND2X2 U11291 ( .A(n22975), .B(n22969), .Y(n6814) );
  AND2X2 U11292 ( .A(n19567), .B(n7861), .Y(n19571) );
  AOI21X1 U11293 ( .A0(n23043), .A1(n23041), .B0(n22940), .Y(n23027) );
  NAND2X1 U11294 ( .A(n6296), .B(n11600), .Y(n11602) );
  AOI21X1 U11295 ( .A0(n25129), .A1(n14490), .B0(n14489), .Y(n25127) );
  AOI21X1 U11296 ( .A0(n14455), .A1(n25160), .B0(n14454), .Y(n14456) );
  AOI21X2 U11297 ( .A0(n7238), .A1(n14424), .B0(n14423), .Y(n6488) );
  NAND2X1 U11298 ( .A(n12186), .B(n12185), .Y(n12209) );
  CLKINVX2 U11299 ( .A(n7426), .Y(n6739) );
  XOR2X1 U11300 ( .A(n13193), .B(n7430), .Y(n13194) );
  NOR2X2 U11301 ( .A(n12195), .B(n12199), .Y(n12206) );
  NAND2BX2 U11302 ( .AN(n12137), .B(n6786), .Y(n6212) );
  OAI21X2 U11303 ( .A0(n23480), .A1(n23479), .B0(n23478), .Y(n23935) );
  NAND2X4 U11304 ( .A(W0[6]), .B(W0[22]), .Y(n9834) );
  AOI21X2 U11305 ( .A0(n12194), .A1(n12206), .B0(n12211), .Y(n12193) );
  OAI21X1 U11306 ( .A0(n23794), .A1(n23793), .B0(n23792), .Y(n23869) );
  NOR2X1 U11307 ( .A(n23431), .B(n23430), .Y(n23474) );
  MXI2X1 U11308 ( .A(U2_pipe1[15]), .B(n23877), .S0(n21700), .Y(n4125) );
  OAI21X1 U11309 ( .A0(n22338), .A1(n6754), .B0(n6753), .Y(n22317) );
  OAI21X1 U11310 ( .A0(n12081), .A1(n12080), .B0(n12079), .Y(n12138) );
  AOI21X2 U11311 ( .A0(n11488), .A1(n11455), .B0(n11454), .Y(n11472) );
  NAND2X4 U11312 ( .A(n28681), .B(n28713), .Y(n7777) );
  XOR2X2 U11313 ( .A(n8268), .B(n28748), .Y(n7339) );
  AOI21X2 U11314 ( .A0(n24868), .A1(n24866), .B0(n13530), .Y(n24862) );
  AOI21X1 U11315 ( .A0(n9639), .A1(n11545), .B0(n7185), .Y(n9640) );
  NOR2X1 U11316 ( .A(n24523), .B(n24529), .Y(n13510) );
  AOI21X2 U11317 ( .A0(n6854), .A1(n13318), .B0(n7230), .Y(n13302) );
  NOR2X2 U11318 ( .A(n6759), .B(n6756), .Y(n7430) );
  OAI21X1 U11319 ( .A0(n22304), .A1(n21961), .B0(n21962), .Y(n13170) );
  MXI2X1 U11320 ( .A(U0_pipe1[22]), .B(n25000), .S0(n25101), .Y(n4262) );
  INVX1 U11321 ( .A(n6277), .Y(n25004) );
  NOR2X1 U11322 ( .A(n22601), .B(n22602), .Y(n14127) );
  NAND2X1 U11323 ( .A(n6318), .B(n9146), .Y(n9148) );
  AOI21X2 U11324 ( .A0(n13140), .A1(n13139), .B0(n6244), .Y(n13151) );
  NOR2X2 U11325 ( .A(n8060), .B(AOPD[35]), .Y(n10989) );
  XOR2X2 U11326 ( .A(n9944), .B(n10334), .Y(U1_U2_z2[12]) );
  INVX1 U11327 ( .A(n10966), .Y(n10955) );
  XNOR2X2 U11328 ( .A(n10878), .B(n10877), .Y(U0_U2_z0[25]) );
  NAND2X1 U11329 ( .A(n12161), .B(n12162), .Y(n12177) );
  OAI21XL U11330 ( .A0(n6878), .A1(n10755), .B0(n10754), .Y(n10760) );
  OAI21XL U11331 ( .A0(n25317), .A1(n25301), .B0(n25300), .Y(n25306) );
  MXI2X1 U11332 ( .A(U0_pipe13[23]), .B(n25307), .S0(n25318), .Y(n4669) );
  NOR2BX1 U11333 ( .AN(n25362), .B(n6382), .Y(n6381) );
  NOR2X1 U11334 ( .A(n12389), .B(n6381), .Y(n25348) );
  NAND2X2 U11335 ( .A(n7324), .B(n7322), .Y(n10839) );
  AOI21X2 U11336 ( .A0(n11607), .A1(n11489), .B0(n11488), .Y(n11494) );
  NAND2X2 U11337 ( .A(n7226), .B(n11430), .Y(n7758) );
  XOR2X2 U11338 ( .A(n9985), .B(n10236), .Y(U1_U1_z2[6]) );
  INVX1 U11339 ( .A(n10478), .Y(n10500) );
  XOR2X1 U11340 ( .A(n7191), .B(n6974), .Y(n14851) );
  NAND2X1 U11341 ( .A(n20051), .B(n19557), .Y(n19588) );
  AND2X2 U11342 ( .A(n19560), .B(n7271), .Y(n7270) );
  INVX1 U11343 ( .A(n9073), .Y(n9149) );
  NOR2X1 U11344 ( .A(n9153), .B(n9149), .Y(n9155) );
  NOR2X1 U11345 ( .A(n22978), .B(n7755), .Y(n22967) );
  NOR2X2 U11346 ( .A(W0[27]), .B(W0[11]), .Y(n9826) );
  OAI2BB1X2 U11347 ( .A0N(n9870), .A1N(n9871), .B0(n6337), .Y(n9872) );
  NAND2X1 U11348 ( .A(n8137), .B(BOPD[29]), .Y(n10842) );
  NAND2X1 U11349 ( .A(n11567), .B(n9631), .Y(n9633) );
  OAI21X1 U11350 ( .A0(n11555), .A1(n11548), .B0(n11552), .Y(n11551) );
  INVX4 U11351 ( .A(n10309), .Y(n10324) );
  INVX4 U11352 ( .A(n10761), .Y(n10817) );
  OR2X2 U11353 ( .A(n13185), .B(n6757), .Y(n6756) );
  OAI21X2 U11354 ( .A0(n9520), .A1(n9497), .B0(n9498), .Y(n9496) );
  NAND3X1 U11355 ( .A(n7350), .B(n9721), .C(n7349), .Y(n7676) );
  AOI21X1 U11356 ( .A0(n19117), .A1(n7679), .B0(n9702), .Y(n19104) );
  INVX1 U11357 ( .A(n13699), .Y(n9701) );
  NOR2X2 U11358 ( .A(n12220), .B(n12219), .Y(n12245) );
  INVX1 U11359 ( .A(n9723), .Y(n9724) );
  CLKINVX2 U11360 ( .A(n14579), .Y(n6761) );
  OAI21X1 U11361 ( .A0(n9464), .A1(n9469), .B0(n9465), .Y(n7328) );
  OAI21X2 U11362 ( .A0(n9461), .A1(n9323), .B0(n7327), .Y(n9479) );
  NAND3X2 U11363 ( .A(n6215), .B(n6700), .C(n10233), .Y(n6214) );
  NAND2X1 U11364 ( .A(BOPA[1]), .B(n11428), .Y(n8302) );
  OAI21X1 U11365 ( .A0(n7681), .A1(n9353), .B0(n9354), .Y(n9360) );
  XOR2X4 U11366 ( .A(n6606), .B(n6913), .Y(n8675) );
  ADDHX2 U11367 ( .A(U1_U0_y2[27]), .B(U1_U0_y0[27]), .CO(n8433), .S(n8430) );
  NAND2X2 U11368 ( .A(n8085), .B(AOPB[28]), .Y(n10508) );
  INVX1 U11369 ( .A(n22736), .Y(n22737) );
  AOI21X1 U11370 ( .A0(n22744), .A1(n14157), .B0(n14156), .Y(n22742) );
  NOR2X1 U11371 ( .A(n8678), .B(n16658), .Y(n8680) );
  NOR2X2 U11372 ( .A(n8069), .B(AOPB[32]), .Y(n10485) );
  OAI21X2 U11373 ( .A0(n8576), .A1(n8582), .B0(n8577), .Y(n7544) );
  CLKINVX3 U11374 ( .A(n14102), .Y(n14103) );
  XOR2X1 U11375 ( .A(n16631), .B(n16630), .Y(n16632) );
  NAND2X1 U11376 ( .A(n13486), .B(U2_A_r_d[21]), .Y(n24439) );
  XOR2X2 U11377 ( .A(n7573), .B(n13473), .Y(n14146) );
  OAI21X1 U11378 ( .A0(n10481), .A1(n10486), .B0(n10482), .Y(n8213) );
  NOR2X1 U11379 ( .A(n9287), .B(U1_U0_y1[13]), .Y(n9389) );
  OAI2BB1XL U11380 ( .A0N(n9381), .A1N(n9288), .B0(n9390), .Y(n6514) );
  AOI21X1 U11381 ( .A0(n9379), .A1(n9377), .B0(n9371), .Y(n6716) );
  XNOR2X2 U11382 ( .A(n10473), .B(n10472), .Y(U0_U0_z0[9]) );
  NOR2X1 U11383 ( .A(n6192), .B(n7745), .Y(n19387) );
  NAND2X1 U11384 ( .A(n19450), .B(n6184), .Y(n6183) );
  MXI2X1 U11385 ( .A(n6191), .B(U1_pipe0[26]), .S0(n7096), .Y(n5129) );
  INVX1 U11386 ( .A(n9914), .Y(n9947) );
  NAND2BX1 U11387 ( .AN(n8618), .B(n16993), .Y(n7619) );
  OAI21X4 U11388 ( .A0(n11032), .A1(n11035), .B0(n11033), .Y(n11014) );
  NOR2X1 U11389 ( .A(n7535), .B(n7534), .Y(n7533) );
  AOI21X2 U11390 ( .A0(n8345), .A1(n11277), .B0(n8344), .Y(n11261) );
  NAND2X1 U11391 ( .A(n8114), .B(AOPC[42]), .Y(n11289) );
  OAI21X1 U11392 ( .A0(n9826), .A1(n9857), .B0(n9827), .Y(n9813) );
  XNOR2X1 U11393 ( .A(n17310), .B(n17613), .Y(n17311) );
  NOR2X2 U11394 ( .A(n9748), .B(n9799), .Y(n6395) );
  NAND2X1 U11395 ( .A(n12533), .B(n12532), .Y(n12555) );
  NOR2X2 U11396 ( .A(n8065), .B(AOPD[33]), .Y(n8318) );
  MXI2X1 U11397 ( .A(U0_pipe15[23]), .B(n22607), .S0(n22620), .Y(n4613) );
  XNOR2X4 U11398 ( .A(n9745), .B(n10067), .Y(U2_U0_z2[13]) );
  MXI2X1 U11399 ( .A(U0_pipe15[22]), .B(n22611), .S0(n22620), .Y(n4614) );
  AOI21X2 U11400 ( .A0(n6391), .A1(n9737), .B0(n9736), .Y(n9806) );
  NAND3X1 U11401 ( .A(n22655), .B(n14123), .C(n14113), .Y(n6242) );
  OAI21X1 U11402 ( .A0(n12596), .A1(n12618), .B0(n12622), .Y(n6740) );
  NAND2BX1 U11403 ( .AN(n25006), .B(n6318), .Y(n7753) );
  XNOR2X1 U11404 ( .A(n8849), .B(n8848), .Y(n24595) );
  XOR2X1 U11405 ( .A(n6365), .B(n25012), .Y(n25013) );
  XOR2X2 U11406 ( .A(n7028), .B(n13616), .Y(n19248) );
  NAND2X4 U11407 ( .A(n6140), .B(n6138), .Y(n13616) );
  NOR2X2 U11408 ( .A(n6139), .B(n7277), .Y(n6138) );
  OAI21X2 U11409 ( .A0(n6142), .A1(n13603), .B0(n6141), .Y(n6140) );
  NOR2X1 U11410 ( .A(n19243), .B(n14966), .Y(n17307) );
  XOR2X4 U11411 ( .A(n13633), .B(n13620), .Y(n19243) );
  AOI22XL U11412 ( .A0(n6143), .A1(n7784), .B0(n19568), .B1(n14976), .Y(n7783)
         );
  XOR2X1 U11413 ( .A(n6143), .B(n7931), .Y(n6707) );
  NAND3X1 U11414 ( .A(n6705), .B(n17597), .C(n6704), .Y(n6143) );
  XOR2X2 U11415 ( .A(n13609), .B(n6144), .Y(n14963) );
  AND2X2 U11416 ( .A(n13595), .B(n13607), .Y(n6144) );
  NOR2BX2 U11417 ( .AN(n13589), .B(n13594), .Y(n7940) );
  INVX1 U11418 ( .A(U1_U1_y2[13]), .Y(n12689) );
  XOR2X2 U11419 ( .A(n6148), .B(n12899), .Y(n14935) );
  NAND2X2 U11420 ( .A(n6150), .B(n6149), .Y(n7178) );
  NAND3X2 U11421 ( .A(n6151), .B(n7497), .C(n7496), .Y(n17304) );
  OAI21X1 U11422 ( .A0(n17305), .A1(n17307), .B0(n17308), .Y(n13623) );
  NAND2BX4 U11423 ( .AN(n13593), .B(n7786), .Y(n13082) );
  OAI21X1 U11424 ( .A0(n17632), .A1(n14499), .B0(n14504), .Y(n17630) );
  OAI21X2 U11425 ( .A0(n13012), .A1(n13056), .B0(n13060), .Y(n6154) );
  XOR2X4 U11426 ( .A(n10246), .B(n6999), .Y(U1_U1_z1[10]) );
  INVX8 U11427 ( .A(n6157), .Y(U1_U1_z1[9]) );
  XNOR2X4 U11428 ( .A(n6218), .B(n10228), .Y(n6157) );
  NAND2X1 U11429 ( .A(n8258), .B(n10747), .Y(n6159) );
  OAI21X1 U11430 ( .A0(n10756), .A1(n10754), .B0(n10757), .Y(n10747) );
  NAND2X1 U11431 ( .A(n8177), .B(BOPD[43]), .Y(n10757) );
  NOR2X1 U11432 ( .A(n8177), .B(BOPD[43]), .Y(n10756) );
  NAND2X1 U11433 ( .A(n5869), .B(n19994), .Y(n16849) );
  NAND2X4 U11434 ( .A(n6164), .B(n6161), .Y(n9913) );
  NOR2X4 U11435 ( .A(n6163), .B(n6162), .Y(n6161) );
  NOR2X2 U11436 ( .A(n9915), .B(n9946), .Y(n6163) );
  NAND2X4 U11437 ( .A(n9914), .B(n6165), .Y(n6164) );
  NOR2X2 U11438 ( .A(n9915), .B(n9945), .Y(n6165) );
  NOR2X4 U11439 ( .A(W2[2]), .B(W2[18]), .Y(n9945) );
  NOR2X4 U11440 ( .A(W2[3]), .B(W2[19]), .Y(n9915) );
  OAI21X4 U11441 ( .A0(n9935), .A1(n9937), .B0(n9936), .Y(n9914) );
  NAND2X4 U11442 ( .A(W2[1]), .B(W2[17]), .Y(n9936) );
  NAND2X4 U11443 ( .A(W2[16]), .B(W2[0]), .Y(n9937) );
  NOR2X4 U11444 ( .A(W2[17]), .B(W2[1]), .Y(n9935) );
  XOR2X4 U11445 ( .A(n6166), .B(n10807), .Y(U1_U2_z0[10]) );
  AOI21X1 U11446 ( .A0(n10761), .A1(n10803), .B0(n10804), .Y(n6166) );
  NAND3BX4 U11447 ( .AN(n7239), .B(n6423), .C(n6422), .Y(n10761) );
  NAND2X1 U11448 ( .A(n16808), .B(n7455), .Y(n6168) );
  NOR2X4 U11449 ( .A(n8168), .B(BOPD[27]), .Y(n10857) );
  AOI21X2 U11450 ( .A0(n7830), .A1(n5878), .B0(n7514), .Y(n13030) );
  OAI21X1 U11451 ( .A0(n11297), .A1(n11306), .B0(n11298), .Y(n8337) );
  NAND2X1 U11452 ( .A(n8195), .B(AOPC[41]), .Y(n11298) );
  NAND2X1 U11453 ( .A(n7992), .B(AOPC[40]), .Y(n11306) );
  XOR2X1 U11454 ( .A(n10703), .B(n10702), .Y(U1_U2_z0[25]) );
  NOR2X1 U11455 ( .A(n21268), .B(n21267), .Y(n21307) );
  INVX2 U11456 ( .A(n26646), .Y(n21309) );
  NAND2X2 U11457 ( .A(n21614), .B(n6172), .Y(n6175) );
  NOR2X1 U11458 ( .A(n21657), .B(n6173), .Y(n6172) );
  NAND2X2 U11459 ( .A(n7343), .B(n21572), .Y(n21614) );
  AOI21XL U11460 ( .A0(n21614), .A1(n21575), .B0(n21613), .Y(n21658) );
  NAND2BX1 U11461 ( .AN(n21657), .B(n21613), .Y(n6174) );
  AND4X4 U11462 ( .A(n8356), .B(n8355), .C(n8354), .D(n8240), .Y(n7576) );
  OAI21X4 U11463 ( .A0(n6176), .A1(n11427), .B0(n11405), .Y(U2_B_i[16]) );
  XOR2X1 U11464 ( .A(n11422), .B(n28712), .Y(n6176) );
  NAND2X4 U11465 ( .A(n9607), .B(n7576), .Y(n11422) );
  NOR3X4 U11466 ( .A(n7777), .B(n7332), .C(n7331), .Y(n9607) );
  AOI21X2 U11467 ( .A0(n6178), .A1(n11529), .B0(n11528), .Y(n11533) );
  AOI2BB1X2 U11468 ( .A0N(n11502), .A1N(n6177), .B0(n11534), .Y(n11538) );
  AOI21X1 U11469 ( .A0(n6178), .A1(n11513), .B0(n11512), .Y(n11518) );
  AOI21X2 U11470 ( .A0(n11521), .A1(n6178), .B0(n11520), .Y(n11525) );
  XOR2X2 U11471 ( .A(n11502), .B(n11541), .Y(U2_U0_z0[14]) );
  INVX4 U11472 ( .A(n11502), .Y(n6178) );
  XNOR2X4 U11473 ( .A(n10100), .B(n6181), .Y(U2_U0_z1[15]) );
  OAI21X2 U11474 ( .A0(n9422), .A1(n9427), .B0(n9423), .Y(n9437) );
  NAND2X1 U11475 ( .A(n9311), .B(n9310), .Y(n9423) );
  NOR2X2 U11476 ( .A(n9311), .B(n9310), .Y(n9422) );
  NAND2BX2 U11477 ( .AN(n19451), .B(n6186), .Y(n6185) );
  NOR2X1 U11478 ( .A(n6187), .B(n7747), .Y(n6192) );
  OAI21XL U11479 ( .A0(n6187), .A1(n19075), .B0(n19076), .Y(n14896) );
  XOR2X1 U11480 ( .A(n6187), .B(n19390), .Y(n19391) );
  AOI21X2 U11481 ( .A0(n19392), .A1(n13715), .B0(n13714), .Y(n6187) );
  NOR2X1 U11482 ( .A(n19410), .B(n13706), .Y(n13708) );
  INVX1 U11483 ( .A(n9936), .Y(n6193) );
  NOR2X1 U11484 ( .A(n6193), .B(n9935), .Y(n14992) );
  XOR2X2 U11485 ( .A(n9491), .B(n9500), .Y(n9700) );
  XOR2X2 U11486 ( .A(U1_U0_y0[28]), .B(U1_U0_y1[28]), .Y(n9318) );
  OAI21X4 U11487 ( .A0(n9774), .A1(n9777), .B0(n9775), .Y(n9763) );
  NAND2X2 U11488 ( .A(W3[1]), .B(W3[17]), .Y(n9775) );
  NOR2X4 U11489 ( .A(W3[17]), .B(W3[1]), .Y(n9774) );
  NAND2X1 U11490 ( .A(n28711), .B(n11401), .Y(n7767) );
  NOR2X1 U11491 ( .A(BOPA[42]), .B(BOPA[43]), .Y(n11401) );
  XOR2X1 U11492 ( .A(n6195), .B(BOPA[47]), .Y(n6194) );
  NOR2X1 U11493 ( .A(n11422), .B(n6196), .Y(n6195) );
  OAI21X4 U11494 ( .A0(n6197), .A1(n10301), .B0(n10300), .Y(n10302) );
  XOR2X1 U11495 ( .A(n6197), .B(n10333), .Y(U1_U2_z1[10]) );
  AOI21X4 U11496 ( .A0(n10331), .A1(n10299), .B0(n10298), .Y(n6197) );
  NOR2X2 U11497 ( .A(n11150), .B(n11146), .Y(n8284) );
  NOR2X2 U11498 ( .A(n8188), .B(BOPC[37]), .Y(n11150) );
  NOR2X4 U11499 ( .A(n7947), .B(W2[18]), .Y(n10341) );
  NOR2X4 U11500 ( .A(n8027), .B(W2[19]), .Y(n10266) );
  NAND2X1 U11501 ( .A(n8188), .B(BOPC[37]), .Y(n11151) );
  OAI21X4 U11502 ( .A0(n6198), .A1(n10214), .B0(n10213), .Y(n7582) );
  OAI21X2 U11503 ( .A0(n6198), .A1(n10250), .B0(n10249), .Y(n10254) );
  XOR2X1 U11504 ( .A(n10245), .B(n6198), .Y(U1_U1_z1[12]) );
  AOI21X4 U11505 ( .A0(n6823), .A1(n7584), .B0(n7583), .Y(n6198) );
  NAND2BX1 U11506 ( .AN(n21955), .B(n21956), .Y(n22300) );
  INVX1 U11507 ( .A(n21953), .Y(n6202) );
  INVXL U11508 ( .A(n21954), .Y(n6203) );
  XOR2X2 U11509 ( .A(n6751), .B(n12190), .Y(n14555) );
  NAND2BX1 U11510 ( .AN(n7346), .B(n13125), .Y(n7016) );
  NOR2X2 U11511 ( .A(n12084), .B(n12083), .Y(n12149) );
  NAND2X1 U11512 ( .A(n6204), .B(n11401), .Y(n6340) );
  INVX1 U11513 ( .A(n11422), .Y(n6204) );
  NAND2X1 U11514 ( .A(n6272), .B(n6205), .Y(n6271) );
  NOR2X2 U11515 ( .A(n11422), .B(n6206), .Y(n6205) );
  INVX4 U11516 ( .A(n10988), .Y(n10997) );
  NAND2X4 U11517 ( .A(n6208), .B(n6207), .Y(n10988) );
  AOI21X4 U11518 ( .A0(n8319), .A1(n6375), .B0(n6374), .Y(n6208) );
  XOR2X2 U11519 ( .A(n10997), .B(n10996), .Y(U0_U2_z0[8]) );
  OAI21X4 U11520 ( .A0(n12258), .A1(n12207), .B0(n12212), .Y(n12194) );
  AOI21X4 U11521 ( .A0(n6210), .A1(n12180), .B0(n6209), .Y(n12212) );
  OAI21X2 U11522 ( .A0(n12179), .A1(n12178), .B0(n12177), .Y(n6209) );
  NAND2BX2 U11523 ( .AN(n6785), .B(n6210), .Y(n12207) );
  NOR2X4 U11524 ( .A(n6212), .B(n6211), .Y(n12258) );
  AOI21X4 U11525 ( .A0(n6788), .A1(n7429), .B0(n6787), .Y(n6211) );
  NAND2X2 U11526 ( .A(n6733), .B(n10231), .Y(n6220) );
  NOR2X2 U11527 ( .A(n10256), .B(n10196), .Y(n10231) );
  NOR2X4 U11528 ( .A(n10232), .B(n10198), .Y(n6733) );
  NAND2BX4 U11529 ( .AN(n11443), .B(n11531), .Y(n11444) );
  INVX1 U11530 ( .A(U2_B_r[16]), .Y(n6213) );
  NOR2X2 U11531 ( .A(U2_B_r[17]), .B(n5824), .Y(n11443) );
  OAI21X2 U11532 ( .A0(n8249), .A1(n11427), .B0(n8248), .Y(U2_B_i[17]) );
  XOR2X4 U11533 ( .A(n6214), .B(n10235), .Y(U1_U1_z1[7]) );
  INVX4 U11534 ( .A(n10229), .Y(n10260) );
  AOI21X2 U11535 ( .A0(n6823), .A1(n10226), .B0(n10225), .Y(n6218) );
  OAI21X4 U11536 ( .A0(n10229), .A1(n6220), .B0(n6219), .Y(n6823) );
  AOI21X4 U11537 ( .A0(n10230), .A1(n6733), .B0(n7360), .Y(n6219) );
  AOI21X4 U11538 ( .A0(n6820), .A1(n6735), .B0(n6734), .Y(n10229) );
  NOR2X1 U11539 ( .A(n7061), .B(BOPC[45]), .Y(n11087) );
  NOR2X1 U11540 ( .A(n8176), .B(BOPC[43]), .Y(n11100) );
  NOR2X1 U11541 ( .A(n11104), .B(n11100), .Y(n11092) );
  NOR2X1 U11542 ( .A(n7052), .B(BOPC[42]), .Y(n11104) );
  NOR2X1 U11543 ( .A(n11083), .B(n11087), .Y(n8290) );
  NAND2X4 U11544 ( .A(n8246), .B(n7576), .Y(n9619) );
  NAND2X2 U11545 ( .A(W0[18]), .B(n6876), .Y(n9851) );
  XOR2X1 U11546 ( .A(n10477), .B(n6916), .Y(U0_U0_z0[8]) );
  NOR2X2 U11547 ( .A(n10435), .B(n10441), .Y(n10427) );
  NOR2X2 U11548 ( .A(n8198), .B(AOPB[39]), .Y(n10441) );
  INVX1 U11549 ( .A(n14816), .Y(n14823) );
  NAND2BX4 U11550 ( .AN(n7886), .B(n6130), .Y(n14816) );
  NAND2X1 U11551 ( .A(n14826), .B(n7434), .Y(n20379) );
  XOR2X1 U11552 ( .A(U2_U0_y2[36]), .B(U2_U0_y0[36]), .Y(n24290) );
  OR2X2 U11553 ( .A(n6228), .B(n6730), .Y(n24495) );
  OR2X2 U11554 ( .A(n6228), .B(U2_A_i_d[14]), .Y(n22515) );
  NAND2XL U11555 ( .A(n6228), .B(U2_A_r_d[14]), .Y(n24494) );
  NOR2X1 U11556 ( .A(n6228), .B(n5781), .Y(n14089) );
  NAND2XL U11557 ( .A(n6228), .B(U2_A_i_d[14]), .Y(n22514) );
  NAND2X1 U11558 ( .A(n6228), .B(n5781), .Y(n14090) );
  NAND2X1 U11559 ( .A(n6228), .B(n6227), .Y(n13451) );
  OAI21X4 U11560 ( .A0(n24871), .A1(n24424), .B0(n24425), .Y(n24868) );
  AOI21X4 U11561 ( .A0(n7272), .A1(n24873), .B0(n6229), .Y(n24871) );
  NAND3BX1 U11562 ( .AN(n19598), .B(n7177), .C(n6231), .Y(n6230) );
  XOR2X1 U11563 ( .A(n6232), .B(n19614), .Y(n19615) );
  XOR2X2 U11564 ( .A(n6233), .B(n14778), .Y(n14791) );
  OAI21X1 U11565 ( .A0(n7420), .A1(n14779), .B0(n14780), .Y(n6233) );
  OAI21X2 U11566 ( .A0(n6234), .A1(n11418), .B0(n9608), .Y(U2_B_i[22]) );
  NOR2X1 U11567 ( .A(n11421), .B(n11422), .Y(n6235) );
  NAND2X1 U11568 ( .A(n8198), .B(AOPB[39]), .Y(n10442) );
  INVX4 U11569 ( .A(n13427), .Y(n13402) );
  INVX2 U11570 ( .A(n13415), .Y(n13425) );
  NAND2X4 U11571 ( .A(n6236), .B(n13400), .Y(n13415) );
  NAND2BX4 U11572 ( .AN(n13401), .B(n13427), .Y(n6236) );
  NAND2X4 U11573 ( .A(n6523), .B(n6412), .Y(n13427) );
  NAND2X2 U11574 ( .A(n13383), .B(n6565), .Y(n13401) );
  NOR2X2 U11575 ( .A(W0[18]), .B(n6875), .Y(n10155) );
  XOR2X1 U11576 ( .A(n24336), .B(n6237), .Y(n24337) );
  AOI21X4 U11577 ( .A0(n24330), .A1(n24329), .B0(n24328), .Y(n6237) );
  NOR2X2 U11578 ( .A(n13250), .B(n13251), .Y(n13323) );
  AOI21X4 U11579 ( .A0(n14127), .A1(n22599), .B0(n6241), .Y(n22597) );
  OAI21X1 U11580 ( .A0(n22600), .A1(n22602), .B0(n22603), .Y(n6241) );
  AOI21X1 U11581 ( .A0(n14124), .A1(n14126), .B0(n14125), .Y(n22600) );
  NAND2X1 U11582 ( .A(n14123), .B(n14122), .Y(n6243) );
  XOR2X1 U11583 ( .A(n11099), .B(n11098), .Y(U1_U1_z0[18]) );
  OAI21X1 U11584 ( .A0(n13138), .A1(n13137), .B0(n13136), .Y(n6244) );
  OAI21X2 U11585 ( .A0(n12640), .A1(n12639), .B0(n12638), .Y(n13139) );
  NOR2X2 U11586 ( .A(n12644), .B(n12645), .Y(n13138) );
  OAI21X4 U11587 ( .A0(n6245), .A1(n13173), .B0(n13172), .Y(n13181) );
  AOI21X4 U11588 ( .A0(n13161), .A1(n13155), .B0(n13160), .Y(n6245) );
  NAND2X1 U11589 ( .A(n8136), .B(BOPC[29]), .Y(n11198) );
  NOR2X2 U11590 ( .A(n11202), .B(n11197), .Y(n6295) );
  NOR2X2 U11591 ( .A(n8136), .B(BOPC[29]), .Y(n11197) );
  NOR2X2 U11592 ( .A(n8138), .B(BOPC[28]), .Y(n11202) );
  OAI21X4 U11593 ( .A0(n11187), .A1(n11192), .B0(n11188), .Y(n11174) );
  NAND2X1 U11594 ( .A(n8127), .B(BOPC[31]), .Y(n11188) );
  NAND2X2 U11595 ( .A(n8133), .B(BOPC[30]), .Y(n11192) );
  XOR2X4 U11596 ( .A(n6246), .B(n6816), .Y(n22973) );
  AOI21X4 U11597 ( .A0(n22967), .A1(n6795), .B0(n6247), .Y(n22975) );
  OAI21X2 U11598 ( .A0(n22977), .A1(n7755), .B0(n22966), .Y(n6247) );
  OAI21X4 U11599 ( .A0(n22999), .A1(n22956), .B0(n22955), .Y(n6795) );
  OAI21X2 U11600 ( .A0(n11364), .A1(n11369), .B0(n11365), .Y(n11350) );
  NAND2X1 U11601 ( .A(n8070), .B(AOPC[31]), .Y(n11365) );
  NAND2X1 U11602 ( .A(n8074), .B(AOPC[30]), .Y(n11369) );
  OAI21X1 U11603 ( .A0(n27031), .A1(n27030), .B0(n27029), .Y(n27039) );
  AOI21X2 U11604 ( .A0(n26989), .A1(n26988), .B0(n26987), .Y(n27031) );
  OAI2BB1X4 U11605 ( .A0N(n7539), .A1N(n26907), .B0(n6248), .Y(n26989) );
  AND2X4 U11606 ( .A(n7538), .B(n26946), .Y(n6248) );
  NOR2X1 U11607 ( .A(n12640), .B(n12637), .Y(n13135) );
  NOR2X1 U11608 ( .A(n12628), .B(n12629), .Y(n12637) );
  NOR2X2 U11609 ( .A(n12631), .B(n12630), .Y(n12640) );
  NOR2X1 U11610 ( .A(n22990), .B(n6249), .Y(n22983) );
  OAI21X1 U11611 ( .A0(n6249), .A1(n22989), .B0(n22963), .Y(n22984) );
  NOR2X1 U11612 ( .A(n22962), .B(n24680), .Y(n6249) );
  AOI21X1 U11613 ( .A0(n6391), .A1(n9768), .B0(n9767), .Y(n9792) );
  OAI21X4 U11614 ( .A0(n6393), .A1(n9746), .B0(n6250), .Y(n6391) );
  AOI21X4 U11615 ( .A0(n9763), .A1(n6397), .B0(n6396), .Y(n9746) );
  NAND3BXL U11616 ( .AN(n6419), .B(n6258), .C(n18986), .Y(n6257) );
  MXI2X1 U11617 ( .A(n6260), .B(U2_pipe3[25]), .S0(n5929), .Y(n4249) );
  NAND2XL U11618 ( .A(n6261), .B(n23923), .Y(n23931) );
  AOI21X1 U11619 ( .A0(n23929), .A1(n6261), .B0(n23928), .Y(n23930) );
  NOR2X1 U11620 ( .A(n23922), .B(n23927), .Y(n6261) );
  OAI2BB1X4 U11621 ( .A0N(n6264), .A1N(n24247), .B0(n6263), .Y(n24330) );
  AOI21X4 U11622 ( .A0(n9991), .A1(n9967), .B0(n9966), .Y(n9985) );
  NAND2X4 U11623 ( .A(n6266), .B(n6265), .Y(n9991) );
  AOI2BB1X4 U11624 ( .A0N(n9977), .A1N(n10007), .B0(n7276), .Y(n6265) );
  NAND2X4 U11625 ( .A(n9976), .B(n6267), .Y(n6266) );
  NOR2X2 U11626 ( .A(n9977), .B(n10006), .Y(n6267) );
  OAI21X4 U11627 ( .A0(n10002), .A1(n10005), .B0(n10003), .Y(n9976) );
  XOR2X2 U11628 ( .A(n11079), .B(n11078), .Y(U1_U1_z0[21]) );
  AOI21X1 U11629 ( .A0(n18816), .A1(n18701), .B0(n18706), .Y(n18649) );
  NAND2X1 U11630 ( .A(n8176), .B(BOPC[43]), .Y(n11101) );
  XOR2X1 U11631 ( .A(n6271), .B(n28684), .Y(n6270) );
  OAI21X2 U11632 ( .A0(n6273), .A1(n8294), .B0(n8293), .Y(n11214) );
  OAI21X1 U11633 ( .A0(n8289), .A1(n11080), .B0(n6273), .Y(n7562) );
  NAND2BX2 U11634 ( .AN(n8948), .B(n8953), .Y(n7183) );
  NOR2X2 U11635 ( .A(n8900), .B(n8898), .Y(n6368) );
  NOR2X2 U11636 ( .A(n8744), .B(n8745), .Y(n8900) );
  NOR2X2 U11637 ( .A(n8740), .B(n8741), .Y(n8840) );
  NAND2X1 U11638 ( .A(n24664), .B(n24663), .Y(n24738) );
  XOR2X2 U11639 ( .A(n9077), .B(n9076), .Y(n24663) );
  AOI21X2 U11640 ( .A0(n7727), .A1(n9163), .B0(n9167), .Y(n9077) );
  XOR2X4 U11641 ( .A(n6274), .B(n9111), .Y(n24644) );
  AOI21X4 U11642 ( .A0(n9118), .A1(n9096), .B0(n9095), .Y(n9107) );
  CLKINVX2 U11643 ( .A(n6278), .Y(n6276) );
  NOR2X1 U11644 ( .A(n9148), .B(n25006), .Y(n6278) );
  NAND3BX2 U11645 ( .AN(n9061), .B(n6774), .C(n9062), .Y(n6311) );
  NAND2X2 U11646 ( .A(n9059), .B(n9096), .Y(n9061) );
  NOR2X4 U11647 ( .A(n9108), .B(n9106), .Y(n9059) );
  AND2X2 U11648 ( .A(U0_U1_y1[29]), .B(U0_U1_y0[29]), .Y(n9057) );
  XOR2X4 U11649 ( .A(n6279), .B(n10308), .Y(U1_U2_z1[9]) );
  AOI21X2 U11650 ( .A0(n10331), .A1(n10306), .B0(n10305), .Y(n6279) );
  OAI21X4 U11651 ( .A0(n10309), .A1(n6281), .B0(n6280), .Y(n10331) );
  AOI21X4 U11652 ( .A0(n10310), .A1(n7193), .B0(n7192), .Y(n6280) );
  NAND2X2 U11653 ( .A(n10311), .B(n7193), .Y(n6281) );
  AOI21X4 U11654 ( .A0(n7196), .A1(n10339), .B0(n7194), .Y(n10309) );
  AOI21X2 U11655 ( .A0(n9934), .A1(n9885), .B0(n6755), .Y(n6831) );
  NAND2X4 U11656 ( .A(n6284), .B(n6282), .Y(n9934) );
  AOI21X4 U11657 ( .A0(n7391), .A1(n6285), .B0(n6283), .Y(n6282) );
  OAI21X4 U11658 ( .A0(n9907), .A1(n9911), .B0(n9908), .Y(n7391) );
  NAND3X4 U11659 ( .A(n9913), .B(n6285), .C(n9896), .Y(n6284) );
  NOR2X2 U11660 ( .A(n9907), .B(n9905), .Y(n9896) );
  NOR2X2 U11661 ( .A(n9897), .B(n9901), .Y(n6285) );
  OAI21X4 U11662 ( .A0(n6286), .A1(n9856), .B0(n9857), .Y(n7267) );
  XOR2X4 U11663 ( .A(n6286), .B(n10175), .Y(U0_U0_z2[10]) );
  NOR2X4 U11664 ( .A(n7265), .B(n7263), .Y(n6286) );
  XOR2X1 U11665 ( .A(n9615), .B(BOPA[30]), .Y(n6287) );
  NOR2X4 U11666 ( .A(n8309), .B(n6288), .Y(n9615) );
  NAND2X2 U11667 ( .A(n29103), .B(n29102), .Y(n6288) );
  NAND2X4 U11668 ( .A(n28751), .B(n28682), .Y(n8309) );
  OAI2BB2X4 U11669 ( .B0(n10266), .B1(n10340), .A0N(n8027), .A1N(W2[19]), .Y(
        n7194) );
  XOR2X1 U11670 ( .A(n10338), .B(n6289), .Y(U1_U2_z1[6]) );
  AOI21X4 U11671 ( .A0(n10324), .A1(n10311), .B0(n10310), .Y(n6289) );
  NOR2X2 U11672 ( .A(n6944), .B(BOPB[40]), .Y(n10600) );
  XOR2X2 U11673 ( .A(n9074), .B(n6973), .Y(n24664) );
  NAND3X2 U11674 ( .A(n7336), .B(n9033), .C(n7335), .Y(n9074) );
  AOI21X2 U11675 ( .A0(n6535), .A1(n13135), .B0(n13139), .Y(n6290) );
  OAI21X4 U11676 ( .A0(n11173), .A1(n6292), .B0(n6291), .Y(n11107) );
  AOI21X4 U11677 ( .A0(n6293), .A1(n11174), .B0(n7286), .Y(n6291) );
  NAND2X2 U11678 ( .A(n11175), .B(n6293), .Y(n6292) );
  NOR2X4 U11679 ( .A(n11176), .B(n11181), .Y(n6293) );
  AOI21X4 U11680 ( .A0(n11196), .A1(n6295), .B0(n6294), .Y(n11173) );
  OAI21X2 U11681 ( .A0(n11197), .A1(n11203), .B0(n11198), .Y(n6294) );
  OAI21X4 U11682 ( .A0(n11218), .A1(n7293), .B0(n11219), .Y(n11196) );
  CLKINVX8 U11683 ( .A(U2_factor_reg), .Y(n8242) );
  NOR2X1 U11684 ( .A(n9175), .B(n9178), .Y(n6297) );
  AOI21X1 U11685 ( .A0(n6528), .A1(n6301), .B0(n5842), .Y(n6300) );
  INVX1 U11686 ( .A(n24987), .Y(n6301) );
  NAND2XL U11687 ( .A(n25289), .B(n12403), .Y(n6308) );
  NAND3X2 U11688 ( .A(n6303), .B(n6302), .C(n12405), .Y(n7733) );
  NAND2X1 U11689 ( .A(n6305), .B(n12402), .Y(n6303) );
  NAND2XL U11690 ( .A(n6308), .B(n6304), .Y(n6307) );
  XOR2X1 U11691 ( .A(n6307), .B(n6306), .Y(n25288) );
  NOR2X4 U11692 ( .A(n9119), .B(n9127), .Y(n9096) );
  NOR2X2 U11693 ( .A(n9050), .B(n9051), .Y(n9127) );
  NOR2X4 U11694 ( .A(n9054), .B(n9055), .Y(n9106) );
  XOR2X2 U11695 ( .A(U0_U1_y1[29]), .B(U0_U1_y0[29]), .Y(n9054) );
  NOR2X4 U11696 ( .A(n9056), .B(n9057), .Y(n9108) );
  NAND3X2 U11697 ( .A(n6311), .B(n9060), .C(n6310), .Y(n7727) );
  NAND2X2 U11698 ( .A(n6772), .B(n6773), .Y(n6310) );
  AOI2BB2X1 U11699 ( .B0(n14562), .B1(n24642), .A0N(n6385), .A1N(n6312), .Y(
        n25323) );
  INVX1 U11700 ( .A(n12394), .Y(n6312) );
  NAND3X1 U11701 ( .A(n6435), .B(n9060), .C(n6316), .Y(n6315) );
  NAND2X1 U11702 ( .A(n9051), .B(n9050), .Y(n9128) );
  AOI22X1 U11703 ( .A0(n7733), .A1(n6317), .B0(n5815), .B1(n7729), .Y(n25287)
         );
  NOR2X1 U11704 ( .A(n9140), .B(n25027), .Y(n6318) );
  NAND2X1 U11705 ( .A(n8104), .B(AOPB[27]), .Y(n10525) );
  OAI21X4 U11706 ( .A0(n6319), .A1(n11427), .B0(n9553), .Y(U2_B_i[7]) );
  XNOR2X2 U11707 ( .A(n6320), .B(n29100), .Y(n6319) );
  NOR2X2 U11708 ( .A(n9552), .B(BOPA[32]), .Y(n6320) );
  XOR2X4 U11709 ( .A(n6321), .B(n9122), .Y(n24646) );
  AOI21X2 U11710 ( .A0(n9118), .A1(n5895), .B0(n6322), .Y(n6321) );
  NAND2X4 U11711 ( .A(n6478), .B(n9093), .Y(n9118) );
  INVXL U11712 ( .A(U2_B_r[2]), .Y(n6323) );
  OR2X2 U11713 ( .A(n11608), .B(U2_B_r[3]), .Y(n11593) );
  AOI21X4 U11714 ( .A0(n6324), .A1(n11428), .B0(n6937), .Y(n11608) );
  NAND2X2 U11715 ( .A(n6325), .B(n11600), .Y(n11599) );
  NAND2X1 U11716 ( .A(n8308), .B(U2_B_r[1]), .Y(n11600) );
  XOR2X2 U11717 ( .A(n6327), .B(n10484), .Y(U0_U0_z0[7]) );
  OAI21X1 U11718 ( .A0(n10489), .A1(n10485), .B0(n10486), .Y(n6327) );
  NOR2X2 U11719 ( .A(n6328), .B(n10479), .Y(n10489) );
  NOR2X1 U11720 ( .A(n10478), .B(n6329), .Y(n6328) );
  XOR2X1 U11721 ( .A(n11425), .B(n28687), .Y(n6330) );
  NOR2X1 U11722 ( .A(n11422), .B(n6407), .Y(n6331) );
  OAI21X4 U11723 ( .A0(n21950), .A1(n14581), .B0(n14580), .Y(n6805) );
  AOI21X4 U11724 ( .A0(n6446), .A1(n21952), .B0(n6332), .Y(n21950) );
  OAI21X4 U11725 ( .A0(n21953), .A1(n6447), .B0(n14578), .Y(n6332) );
  NAND3X2 U11726 ( .A(n6539), .B(n6540), .C(n6537), .Y(n21952) );
  NOR2X4 U11727 ( .A(n12064), .B(n12065), .Y(n12094) );
  AOI21X1 U11728 ( .A0(n14514), .A1(n22059), .B0(n14528), .Y(n6333) );
  OAI21XL U11729 ( .A0(n22067), .A1(n22073), .B0(n22068), .Y(n22059) );
  NAND2XL U11730 ( .A(n14525), .B(n22886), .Y(n22073) );
  NOR2X1 U11731 ( .A(n14526), .B(n22885), .Y(n22067) );
  AOI21X4 U11732 ( .A0(n5923), .A1(n6336), .B0(n6335), .Y(n6337) );
  NAND2X1 U11733 ( .A(n9866), .B(n9863), .Y(n9868) );
  AOI21X2 U11734 ( .A0(n9814), .A1(n9824), .B0(n9813), .Y(n9869) );
  OAI21X4 U11735 ( .A0(n9829), .A1(n7281), .B0(n7280), .Y(n9870) );
  AOI21X4 U11736 ( .A0(n9830), .A1(n7373), .B0(n7372), .Y(n7280) );
  NAND3X4 U11737 ( .A(n5839), .B(n5932), .C(n7374), .Y(n7281) );
  AOI21X4 U11738 ( .A0(n9845), .A1(n7261), .B0(n7260), .Y(n9829) );
  NOR2X4 U11739 ( .A(n7974), .B(W2[26]), .Y(n10301) );
  XOR2X2 U11740 ( .A(n6338), .B(n24378), .Y(n24379) );
  OAI21X4 U11741 ( .A0(n6339), .A1(n11427), .B0(n11402), .Y(U2_B_i[18]) );
  XOR2X2 U11742 ( .A(n6340), .B(n28711), .Y(n6339) );
  NOR2X1 U11743 ( .A(n23745), .B(n23744), .Y(n23791) );
  XOR2X4 U11744 ( .A(n6342), .B(n24698), .Y(n6341) );
  OAI21X2 U11745 ( .A0(n7284), .A1(n24704), .B0(n24705), .Y(n6342) );
  AOI21X2 U11746 ( .A0(n9203), .A1(n9190), .B0(n9202), .Y(n6846) );
  NAND2X4 U11747 ( .A(n6348), .B(n6347), .Y(n9203) );
  AOI2BB1X2 U11748 ( .A0N(n9187), .A1N(n9186), .B0(n6358), .Y(n6347) );
  INVX4 U11749 ( .A(n6351), .Y(n24633) );
  NOR2X4 U11750 ( .A(n6819), .B(n6818), .Y(n9189) );
  OAI21X2 U11751 ( .A0(n6844), .A1(n9013), .B0(n9015), .Y(n6354) );
  OAI2BB1X2 U11752 ( .A0N(n5891), .A1N(n6376), .B0(n6352), .Y(n6844) );
  NAND3BX2 U11753 ( .AN(n6819), .B(n6353), .C(n5891), .Y(n6352) );
  INVX1 U11754 ( .A(n6818), .Y(n6353) );
  XNOR2X4 U11755 ( .A(n6354), .B(n8998), .Y(n6351) );
  NOR2BX1 U11756 ( .AN(U0_U2_y1[16]), .B(n6355), .Y(n8743) );
  NAND2X1 U11757 ( .A(n5881), .B(n6357), .Y(n6356) );
  NAND2X2 U11758 ( .A(n9203), .B(n6851), .Y(n6850) );
  XOR2X4 U11759 ( .A(n12350), .B(n9237), .Y(n24693) );
  AOI21X4 U11760 ( .A0(n9233), .A1(n9221), .B0(n9232), .Y(n12350) );
  AOI21X1 U11761 ( .A0(n25046), .A1(n25030), .B0(n25029), .Y(n25036) );
  INVX1 U11762 ( .A(U0_U2_y1[13]), .Y(n8732) );
  NAND2X1 U11763 ( .A(n8744), .B(n8745), .Y(n8901) );
  NAND2BX2 U11764 ( .AN(n8736), .B(n6369), .Y(n8953) );
  OAI21X1 U11765 ( .A0(n6370), .A1(n8860), .B0(n8737), .Y(n6369) );
  OAI21X2 U11766 ( .A0(n7284), .A1(n6531), .B0(n6530), .Y(n6528) );
  OAI21X4 U11767 ( .A0(n9189), .A1(n9100), .B0(n9099), .Y(n9123) );
  OAI21X2 U11768 ( .A0(n8318), .A1(n10999), .B0(n8317), .Y(n6374) );
  NAND2X1 U11769 ( .A(n6373), .B(n10995), .Y(n10993) );
  NAND2XL U11770 ( .A(n10988), .B(n10987), .Y(n6373) );
  OAI21X2 U11771 ( .A0(n11010), .A1(n11005), .B0(n11006), .Y(n8319) );
  NOR2X2 U11772 ( .A(n8318), .B(n10998), .Y(n6375) );
  NAND2X4 U11773 ( .A(n7206), .B(n7205), .Y(n11013) );
  XOR2X1 U11774 ( .A(n8825), .B(n8817), .Y(n24606) );
  OAI21X1 U11775 ( .A0(n22597), .A1(n22595), .B0(n22596), .Y(n7419) );
  OAI21X4 U11776 ( .A0(n11015), .A1(n11038), .B0(n11016), .Y(n7144) );
  NAND2X2 U11777 ( .A(AOPD[28]), .B(n5777), .Y(n11038) );
  NOR2X4 U11778 ( .A(n8080), .B(AOPD[29]), .Y(n11015) );
  AOI21X1 U11779 ( .A0(n22655), .A1(n14113), .B0(n14122), .Y(n22623) );
  NAND2X1 U11780 ( .A(n12580), .B(n22657), .Y(n6377) );
  NAND2BX1 U11781 ( .AN(n10973), .B(n10988), .Y(n6378) );
  AOI21X4 U11782 ( .A0(n9934), .A1(n9877), .B0(n9876), .Y(n9944) );
  OR2X2 U11783 ( .A(n25348), .B(n12393), .Y(n6380) );
  INVXL U11784 ( .A(n25364), .Y(n6382) );
  OAI21X1 U11785 ( .A0(n25323), .A1(n12396), .B0(n12395), .Y(n6384) );
  INVXL U11786 ( .A(n6942), .Y(n6385) );
  OAI21X2 U11787 ( .A0(n12203), .A1(n12199), .B0(n12200), .Y(n6386) );
  NAND2BX2 U11788 ( .AN(n12134), .B(n12139), .Y(n6788) );
  NOR2X1 U11789 ( .A(n12058), .B(n12059), .Y(n12121) );
  NOR2X1 U11790 ( .A(n12061), .B(n12060), .Y(n12123) );
  NOR2X4 U11791 ( .A(n12094), .B(n12092), .Y(n12067) );
  XOR2X4 U11792 ( .A(n6387), .B(n12145), .Y(n13114) );
  AOI21X2 U11793 ( .A0(n5875), .A1(n12146), .B0(n12142), .Y(n6387) );
  AOI21X1 U11794 ( .A0(n25334), .A1(n25326), .B0(n25325), .Y(n6388) );
  OAI21X1 U11795 ( .A0(n25336), .A1(n25324), .B0(n25323), .Y(n25334) );
  AOI21X1 U11796 ( .A0(n25370), .A1(n25322), .B0(n25321), .Y(n25336) );
  NOR2X2 U11797 ( .A(n7992), .B(AOPC[40]), .Y(n11305) );
  OAI21X2 U11798 ( .A0(n6389), .A1(n29106), .B0(n9616), .Y(U2_B_i[5]) );
  XOR2X4 U11799 ( .A(n6390), .B(n29105), .Y(n6389) );
  NOR2X4 U11800 ( .A(n10315), .B(n10267), .Y(n10311) );
  NOR2X4 U11801 ( .A(n7942), .B(W2[21]), .Y(n10267) );
  AOI21X1 U11802 ( .A0(n6391), .A1(n9798), .B0(n9785), .Y(n6405) );
  XOR2X1 U11803 ( .A(n6391), .B(n10102), .Y(U2_U0_z2[8]) );
  NOR2X4 U11804 ( .A(W3[19]), .B(W3[3]), .Y(n9764) );
  NOR2X2 U11805 ( .A(n9764), .B(n9793), .Y(n6397) );
  NOR2X2 U11806 ( .A(W3[2]), .B(W3[18]), .Y(n9793) );
  BUFX2 U11807 ( .A(n9806), .Y(n6398) );
  OAI21X2 U11808 ( .A0(n9802), .A1(n9799), .B0(n9800), .Y(n6399) );
  NOR2X1 U11809 ( .A(n11422), .B(n7767), .Y(n6404) );
  NAND2X2 U11810 ( .A(n6406), .B(n10043), .Y(n10021) );
  NOR2X1 U11811 ( .A(n11425), .B(BOPA[50]), .Y(n7769) );
  XOR2X4 U11812 ( .A(n6408), .B(n8210), .Y(U0_U2_z0[7]) );
  AOI21X1 U11813 ( .A0(n11013), .A1(n8316), .B0(n8319), .Y(n11002) );
  OAI21X4 U11814 ( .A0(n10295), .A1(n10276), .B0(n10275), .Y(n10289) );
  NOR2X2 U11815 ( .A(n8031), .B(W2[29]), .Y(n10276) );
  NAND2X2 U11816 ( .A(n7988), .B(W2[28]), .Y(n10295) );
  INVX2 U11817 ( .A(n10328), .Y(U1_U2_z1[16]) );
  NAND2X4 U11818 ( .A(W0[17]), .B(W0[1]), .Y(n10160) );
  INVX8 U11819 ( .A(n6409), .Y(U0_U0_z2[9]) );
  XNOR2X4 U11820 ( .A(n6410), .B(n10137), .Y(n6409) );
  AOI21X2 U11821 ( .A0(n9870), .A1(n9855), .B0(n8352), .Y(n6410) );
  OAI21X4 U11822 ( .A0(n11399), .A1(n11396), .B0(n11397), .Y(n11373) );
  NOR2X2 U11823 ( .A(n8102), .B(AOPC[27]), .Y(n11396) );
  NOR2X2 U11824 ( .A(n8206), .B(AOPC[26]), .Y(n11399) );
  OAI21X2 U11825 ( .A0(n13303), .A1(n5903), .B0(n13302), .Y(n6413) );
  NAND2X2 U11826 ( .A(n6854), .B(n13317), .Y(n13303) );
  AOI21X1 U11827 ( .A0(n24421), .A1(n13493), .B0(n13492), .Y(n6414) );
  OAI21X1 U11828 ( .A0(n6414), .A1(n24416), .B0(n24417), .Y(n24413) );
  XOR2XL U11829 ( .A(n24419), .B(n6414), .Y(n24420) );
  NOR2X4 U11830 ( .A(n8187), .B(BOPB[37]), .Y(n10624) );
  AOI21X4 U11831 ( .A0(n13415), .A1(n13404), .B0(n13403), .Y(n13413) );
  NOR2X4 U11832 ( .A(BOPA[26]), .B(BOPA[28]), .Y(n8356) );
  XOR2X1 U11833 ( .A(n6419), .B(n6418), .Y(n18946) );
  XOR2XL U11834 ( .A(n18980), .B(n18979), .Y(n6418) );
  OAI21X2 U11835 ( .A0(n6420), .A1(n11427), .B0(n9620), .Y(U2_B_i[12]) );
  OAI21X4 U11836 ( .A0(n10857), .A1(n6421), .B0(n10858), .Y(n10840) );
  XOR2X1 U11837 ( .A(n10860), .B(n6421), .Y(U1_U2_z0[1]) );
  NOR2X4 U11838 ( .A(n7991), .B(BOPD[26]), .Y(n6421) );
  OAI21X1 U11839 ( .A0(n10817), .A1(n10797), .B0(n10796), .Y(n10802) );
  NAND3X2 U11840 ( .A(n10839), .B(n8251), .C(n10819), .Y(n6423) );
  INVX1 U11841 ( .A(n10373), .Y(n10381) );
  AOI21X1 U11842 ( .A0(n10519), .A1(n10349), .B0(n10348), .Y(n10350) );
  NAND2BX1 U11843 ( .AN(n8235), .B(n10373), .Y(n6424) );
  NAND2X2 U11844 ( .A(n7057), .B(AOPB[42]), .Y(n10410) );
  INVX2 U11845 ( .A(n26515), .Y(n21190) );
  XOR2X4 U11846 ( .A(n6426), .B(n21699), .Y(n21701) );
  NOR2X1 U11847 ( .A(n10387), .B(n10391), .Y(n8226) );
  AOI21X1 U11848 ( .A0(n10373), .A1(n10355), .B0(n10357), .Y(n8227) );
  NOR2X1 U11849 ( .A(n6430), .B(n6431), .Y(n12144) );
  XNOR2X1 U11850 ( .A(U0_U2_y2[23]), .B(n6431), .Y(n12140) );
  NAND2BX1 U11851 ( .AN(n22934), .B(n14547), .Y(n22010) );
  AOI21XL U11852 ( .A0(n21988), .A1(n21983), .B0(n21982), .Y(n21985) );
  OAI21XL U11853 ( .A0(n21990), .A1(n21981), .B0(n21980), .Y(n21988) );
  AOI21X1 U11854 ( .A0(n22022), .A1(n21979), .B0(n21978), .Y(n21990) );
  NOR2X1 U11855 ( .A(n14559), .B(n22000), .Y(n21979) );
  AOI2BB1X2 U11856 ( .A0N(n9179), .A1N(n9178), .B0(n6433), .Y(n6432) );
  AOI21X1 U11857 ( .A0(n9167), .A1(n9168), .B0(n6434), .Y(n9179) );
  OAI21XL U11858 ( .A0(n9166), .A1(n9165), .B0(n9164), .Y(n6434) );
  OAI21X1 U11859 ( .A0(n9084), .A1(n9091), .B0(n9085), .Y(n9167) );
  AOI21X4 U11860 ( .A0(n9048), .A1(n9049), .B0(n9047), .Y(n9093) );
  NAND3X1 U11861 ( .A(n6438), .B(n12343), .C(n6437), .Y(n6436) );
  INVXL U11862 ( .A(n9214), .Y(n6439) );
  NOR2XL U11863 ( .A(n9214), .B(n6444), .Y(n6440) );
  NOR2XL U11864 ( .A(n6444), .B(n12344), .Y(n6441) );
  NOR2X4 U11865 ( .A(n6445), .B(n6448), .Y(n21953) );
  NOR2X2 U11866 ( .A(n22960), .B(n14577), .Y(n6447) );
  CLKINVX3 U11867 ( .A(n22965), .Y(n22960) );
  NAND2X1 U11868 ( .A(n12642), .B(n12641), .Y(n13137) );
  NAND2X2 U11869 ( .A(n6455), .B(n12242), .Y(n12252) );
  NAND2BX1 U11870 ( .AN(n12256), .B(n7244), .Y(n6453) );
  AOI21X1 U11871 ( .A0(n6455), .A1(n12246), .B0(n6454), .Y(n12256) );
  OAI21XL U11872 ( .A0(n12245), .A1(n12244), .B0(n12243), .Y(n6454) );
  OAI21X2 U11873 ( .A0(n12225), .A1(n12230), .B0(n12226), .Y(n12246) );
  NOR2X2 U11874 ( .A(n12245), .B(n7240), .Y(n6455) );
  NAND2XL U11875 ( .A(n14579), .B(n22968), .Y(n21948) );
  XOR2X2 U11876 ( .A(n13188), .B(n6536), .Y(n22968) );
  AOI21X2 U11877 ( .A0(n13181), .A1(n13174), .B0(n13180), .Y(n13188) );
  XOR2X2 U11878 ( .A(n12357), .B(n12284), .Y(n14579) );
  AOI21X2 U11879 ( .A0(n12280), .A1(n12274), .B0(n12279), .Y(n12357) );
  OAI21X2 U11880 ( .A0(n12273), .A1(n12272), .B0(n12271), .Y(n12280) );
  AND2X2 U11881 ( .A(U0_U2_y0[27]), .B(U0_U2_y2[27]), .Y(n12184) );
  XOR2X1 U11882 ( .A(U0_U2_y2[27]), .B(U0_U2_y0[27]), .Y(n12181) );
  NOR2BX2 U11883 ( .AN(n12253), .B(n12258), .Y(n7243) );
  NOR2X2 U11884 ( .A(n12207), .B(n6745), .Y(n12253) );
  NAND2X2 U11885 ( .A(n6466), .B(n12206), .Y(n6745) );
  NOR2X2 U11886 ( .A(n12205), .B(n12210), .Y(n6466) );
  OAI21X1 U11887 ( .A0(n12357), .A1(n12356), .B0(n12355), .Y(n12361) );
  NOR2X1 U11888 ( .A(n25286), .B(n24696), .Y(n6457) );
  OAI21X1 U11889 ( .A0(n6459), .A1(n9987), .B0(n9958), .Y(n6834) );
  XOR2X2 U11890 ( .A(n10586), .B(n10585), .Y(U1_U0_z0[18]) );
  OAI22X4 U11891 ( .A0(n10117), .A1(n10134), .B0(n6461), .B1(n6460), .Y(n10128) );
  INVX1 U11892 ( .A(W0[25]), .Y(n6460) );
  NOR2X4 U11893 ( .A(n8048), .B(W0[25]), .Y(n10117) );
  OAI21X4 U11894 ( .A0(n7406), .A1(n6933), .B0(n6462), .Y(n10001) );
  OAI21X4 U11895 ( .A0(n7976), .A1(n7959), .B0(n7408), .Y(n6462) );
  NAND2BX4 U11896 ( .AN(n10000), .B(n6463), .Y(n7408) );
  NAND3BX2 U11897 ( .AN(n9998), .B(n5772), .C(n7397), .Y(n6463) );
  NAND2X4 U11898 ( .A(n7395), .B(n7396), .Y(n7397) );
  OAI21X4 U11899 ( .A0(n6745), .A1(n12212), .B0(n6464), .Y(n12257) );
  AOI21X2 U11900 ( .A0(n6466), .A1(n12211), .B0(n6465), .Y(n6464) );
  OAI21X1 U11901 ( .A0(n12209), .A1(n12210), .B0(n12208), .Y(n6465) );
  OAI21X4 U11902 ( .A0(n12158), .A1(n12159), .B0(n12157), .Y(n12180) );
  NOR2X2 U11903 ( .A(n12143), .B(n12144), .Y(n12159) );
  NAND2X1 U11904 ( .A(n12141), .B(n12140), .Y(n12158) );
  NOR2X4 U11905 ( .A(n12162), .B(n12161), .Y(n12179) );
  NAND2X1 U11906 ( .A(n9885), .B(n9875), .Y(n9920) );
  OR2X4 U11907 ( .A(n9473), .B(n9476), .Y(n7693) );
  NOR2X2 U11908 ( .A(n9317), .B(n9316), .Y(n9476) );
  XOR2X2 U11909 ( .A(U1_U0_y1[27]), .B(U1_U0_y0[27]), .Y(n9316) );
  NOR2X4 U11910 ( .A(n9318), .B(n9319), .Y(n9473) );
  INVX1 U11911 ( .A(U1_U0_y1[27]), .Y(n6467) );
  NAND2XL U11912 ( .A(n6468), .B(n25308), .Y(n25313) );
  NAND2X1 U11913 ( .A(n25289), .B(n6469), .Y(n6468) );
  NAND3BX2 U11914 ( .AN(n25320), .B(n12397), .C(n25322), .Y(n6470) );
  NAND2X4 U11915 ( .A(n6744), .B(n6471), .Y(n12224) );
  NAND2X2 U11916 ( .A(n12253), .B(n5875), .Y(n6471) );
  CLKINVX3 U11917 ( .A(n13128), .Y(n14560) );
  XOR2X4 U11918 ( .A(n12247), .B(n6472), .Y(n13128) );
  NAND2BX1 U11919 ( .AN(n12229), .B(n12230), .Y(n6472) );
  NAND2X2 U11920 ( .A(n7341), .B(n7639), .Y(n9490) );
  INVX1 U11921 ( .A(n13702), .Y(n9512) );
  NAND2X1 U11922 ( .A(n13702), .B(n5760), .Y(n19107) );
  XOR2X4 U11923 ( .A(n9490), .B(n9489), .Y(n13702) );
  OAI21X1 U11924 ( .A0(n11331), .A1(n11340), .B0(n11332), .Y(n8335) );
  NOR2X2 U11925 ( .A(n8200), .B(AOPC[37]), .Y(n11331) );
  NOR2X4 U11926 ( .A(n8026), .B(W0[19]), .Y(n10108) );
  OAI21XL U11927 ( .A0(n25661), .A1(n25292), .B0(n25293), .Y(n25653) );
  AOI2BB1X2 U11928 ( .A0N(n25661), .A1N(n6475), .B0(n6473), .Y(n25658) );
  NOR2X2 U11929 ( .A(n11327), .B(n11331), .Y(n8336) );
  NOR2X1 U11930 ( .A(n8203), .B(AOPC[36]), .Y(n11327) );
  OAI21X2 U11931 ( .A0(n12234), .A1(n25700), .B0(n12233), .Y(n25678) );
  NOR2X1 U11932 ( .A(n24646), .B(n13123), .Y(n6477) );
  NOR2X1 U11933 ( .A(n8910), .B(n8912), .Y(n8809) );
  NOR2X1 U11934 ( .A(n8807), .B(n8806), .Y(n8912) );
  NOR2X1 U11935 ( .A(n8805), .B(n8804), .Y(n8910) );
  OAI21X2 U11936 ( .A0(n8982), .A1(n8981), .B0(n8980), .Y(n9048) );
  NAND2X1 U11937 ( .A(n8943), .B(n8942), .Y(n8980) );
  NAND2BX2 U11938 ( .AN(n9094), .B(n9062), .Y(n6478) );
  NAND2X4 U11939 ( .A(n6479), .B(n6770), .Y(n9062) );
  OAI2BB1X2 U11940 ( .A0N(n8937), .A1N(n7290), .B0(n7036), .Y(n6479) );
  XNOR2X1 U11941 ( .A(n10323), .B(n10324), .Y(U1_U2_z1[4]) );
  NAND2X2 U11942 ( .A(n6482), .B(n6481), .Y(n6480) );
  OAI22X4 U11943 ( .A0(n10267), .A1(n10316), .B0(W2[5]), .B1(n5758), .Y(n10310) );
  NAND2X2 U11944 ( .A(n7980), .B(W2[20]), .Y(n10316) );
  INVXL U11945 ( .A(n14898), .Y(n19386) );
  NAND2X1 U11946 ( .A(n9065), .B(n9066), .Y(n9085) );
  NAND2X1 U11947 ( .A(n9064), .B(n9063), .Y(n9091) );
  AND2X2 U11948 ( .A(n9341), .B(n7666), .Y(n6484) );
  NOR2X1 U11949 ( .A(n7667), .B(n9528), .Y(n7666) );
  NOR2X1 U11950 ( .A(n9338), .B(n9527), .Y(n7667) );
  NAND3X4 U11951 ( .A(n7725), .B(n9526), .C(n7668), .Y(n7622) );
  NOR2X2 U11952 ( .A(n14240), .B(n14239), .Y(n14410) );
  AOI21X4 U11953 ( .A0(n13313), .A1(n7231), .B0(n6485), .Y(n6523) );
  OAI21X2 U11954 ( .A0(n13373), .A1(n13376), .B0(n13377), .Y(n6485) );
  NAND2X1 U11955 ( .A(n13258), .B(n13257), .Y(n13377) );
  NOR2X4 U11956 ( .A(n13374), .B(n13376), .Y(n7231) );
  NOR2X4 U11957 ( .A(n13257), .B(n13258), .Y(n13376) );
  NOR2BX1 U11958 ( .AN(n14031), .B(U2_A_i_d[10]), .Y(n14078) );
  XOR2X4 U11959 ( .A(n6487), .B(n13369), .Y(n14031) );
  AOI2BB1X2 U11960 ( .A0N(n7084), .A1N(n13402), .B0(n13365), .Y(n6487) );
  NOR2XL U11961 ( .A(n25166), .B(U2_A_i_d[19]), .Y(n22205) );
  XOR2X4 U11962 ( .A(n6488), .B(n14432), .Y(n25166) );
  NAND2BX2 U11963 ( .AN(n14422), .B(n7592), .Y(n7238) );
  XNOR2XL U11964 ( .A(n22180), .B(n22181), .Y(n22182) );
  AOI21X4 U11965 ( .A0(n22185), .A1(n22173), .B0(n22172), .Y(n6697) );
  NAND2X2 U11966 ( .A(n6493), .B(n22163), .Y(n22185) );
  XOR2X2 U11967 ( .A(n10283), .B(n10327), .Y(U1_U2_z1[15]) );
  OAI21X4 U11968 ( .A0(n6542), .A1(n10304), .B0(n10270), .Y(n10298) );
  NAND2X2 U11969 ( .A(n8011), .B(W2[24]), .Y(n10304) );
  NOR2X4 U11970 ( .A(n8047), .B(W2[25]), .Y(n6542) );
  NAND2BX2 U11971 ( .AN(n14259), .B(n6489), .Y(n14472) );
  NAND2X2 U11972 ( .A(n6492), .B(n6490), .Y(n6489) );
  NAND2BX2 U11973 ( .AN(n14422), .B(n6491), .Y(n6490) );
  NAND3X1 U11974 ( .A(n14369), .B(n7594), .C(n7593), .Y(n6491) );
  NOR2X1 U11975 ( .A(n14465), .B(n14463), .Y(n6492) );
  NAND2X1 U11976 ( .A(n14256), .B(n14424), .Y(n14463) );
  NAND2BX2 U11977 ( .AN(n22164), .B(n22236), .Y(n6493) );
  OR2X4 U11978 ( .A(n22138), .B(n22139), .Y(n22236) );
  AOI21X4 U11979 ( .A0(n14226), .A1(n6499), .B0(n6494), .Y(n14421) );
  OAI21X2 U11980 ( .A0(n6500), .A1(n14275), .B0(n6495), .Y(n6494) );
  AOI21X2 U11981 ( .A0(n14287), .A1(n6501), .B0(n6496), .Y(n6495) );
  OAI21X1 U11982 ( .A0(n14277), .A1(n14283), .B0(n14278), .Y(n14287) );
  AOI21X2 U11983 ( .A0(n14217), .A1(n14293), .B0(n6497), .Y(n14275) );
  NAND2X1 U11984 ( .A(n14332), .B(n6498), .Y(n14293) );
  OR2X2 U11985 ( .A(n14331), .B(n14328), .Y(n6498) );
  NOR2X2 U11986 ( .A(n6500), .B(n14276), .Y(n6499) );
  NAND2X2 U11987 ( .A(n14288), .B(n6501), .Y(n6500) );
  NOR2X4 U11988 ( .A(n14361), .B(n14359), .Y(n6501) );
  NOR2X1 U11989 ( .A(n14282), .B(n14277), .Y(n14288) );
  NOR2XL U11990 ( .A(n25212), .B(U2_A_i_d[12]), .Y(n21886) );
  OAI21X2 U11991 ( .A0(n14379), .A1(n14375), .B0(n14376), .Y(n6502) );
  AOI21X2 U11992 ( .A0(n14369), .A1(n14368), .B0(n14367), .Y(n14379) );
  XOR2X1 U11993 ( .A(n6504), .B(n22206), .Y(n6503) );
  OAI21XL U11994 ( .A0(n22208), .A1(n22205), .B0(n22204), .Y(n6504) );
  AOI2BB1X2 U11995 ( .A0N(n22212), .A1N(n22201), .B0(n22203), .Y(n22208) );
  AOI21X1 U11996 ( .A0(n14423), .A1(n14256), .B0(n6505), .Y(n14462) );
  OAI21XL U11997 ( .A0(n14425), .A1(n14430), .B0(n14426), .Y(n6505) );
  NAND2X1 U11998 ( .A(n14255), .B(n14254), .Y(n14426) );
  NOR2X2 U11999 ( .A(n14255), .B(n14254), .Y(n14425) );
  NOR2X4 U12000 ( .A(n14251), .B(n14250), .Y(n14434) );
  CLKINVX3 U12001 ( .A(n14482), .Y(n25147) );
  XOR2X1 U12002 ( .A(n14471), .B(n14472), .Y(n14482) );
  NAND2X2 U12003 ( .A(n8047), .B(W2[25]), .Y(n10270) );
  OAI21X2 U12004 ( .A0(n9711), .A1(n6506), .B0(n9710), .Y(n19072) );
  INVX1 U12005 ( .A(n19150), .Y(n6506) );
  NAND2X1 U12006 ( .A(n9686), .B(n19152), .Y(n6507) );
  AOI21X1 U12007 ( .A0(n14486), .A1(n6508), .B0(n14485), .Y(n25130) );
  AOI21X1 U12008 ( .A0(n14132), .A1(n22805), .B0(n14141), .Y(n22773) );
  NAND3X2 U12009 ( .A(n6510), .B(n14084), .C(n6509), .Y(n22805) );
  OR2X2 U12010 ( .A(n22808), .B(n14085), .Y(n6509) );
  NOR2X1 U12011 ( .A(n22809), .B(n14085), .Y(n6511) );
  CLKINVX2 U12012 ( .A(n22805), .Y(n14144) );
  INVX1 U12013 ( .A(n13683), .Y(n9450) );
  NOR2X1 U12014 ( .A(n9676), .B(n19168), .Y(n9679) );
  NOR2XL U12015 ( .A(n9449), .B(U1_A_r_d0[9]), .Y(n19168) );
  INVX1 U12016 ( .A(n13682), .Y(n9449) );
  AND2X2 U12017 ( .A(n6515), .B(n13683), .Y(n9676) );
  NAND2X1 U12018 ( .A(n14242), .B(n14241), .Y(n14404) );
  NAND2XL U12019 ( .A(n6602), .B(n8689), .Y(n6516) );
  AOI21X1 U12020 ( .A0(n16641), .A1(n8686), .B0(n8685), .Y(n7167) );
  NOR2XL U12021 ( .A(n19782), .B(U1_A_i_d0[24]), .Y(n6519) );
  CLKINVX3 U12022 ( .A(n7238), .Y(n14464) );
  NAND2X1 U12023 ( .A(n6520), .B(n14462), .Y(n14469) );
  NAND2X1 U12024 ( .A(n7238), .B(n6521), .Y(n6520) );
  NOR2X1 U12025 ( .A(n10276), .B(n10296), .Y(n10288) );
  NOR2X2 U12026 ( .A(n7988), .B(W2[28]), .Y(n10296) );
  NAND2X1 U12027 ( .A(U1_U0_y1[13]), .B(n6654), .Y(n9286) );
  XOR2X2 U12028 ( .A(U0_U1_y0[30]), .B(U0_U1_y2[30]), .Y(n12597) );
  AND2X2 U12029 ( .A(U0_U1_y2[30]), .B(U0_U1_y0[30]), .Y(n12629) );
  NOR2X2 U12030 ( .A(n9028), .B(n9100), .Y(n9184) );
  NAND2X2 U12031 ( .A(n7726), .B(n7180), .Y(n9100) );
  NOR2X2 U12032 ( .A(n9013), .B(n9016), .Y(n7180) );
  NOR2X2 U12033 ( .A(n7559), .B(n8994), .Y(n9013) );
  NAND2X2 U12034 ( .A(n9026), .B(n9102), .Y(n9028) );
  NOR2X2 U12035 ( .A(n9124), .B(n9131), .Y(n9102) );
  NOR2X2 U12036 ( .A(n9021), .B(n9020), .Y(n9124) );
  NOR2X2 U12037 ( .A(n9115), .B(n9113), .Y(n9026) );
  NOR2X2 U12038 ( .A(n9022), .B(n9023), .Y(n9113) );
  NOR2X4 U12039 ( .A(n9025), .B(n9024), .Y(n9115) );
  INVXL U12040 ( .A(n6524), .Y(n12556) );
  NOR2X2 U12041 ( .A(n6524), .B(n12553), .Y(n12536) );
  NOR2X2 U12042 ( .A(n12533), .B(n12532), .Y(n6524) );
  NOR2BXL U12043 ( .AN(n6532), .B(U0_pipe1[26]), .Y(n6526) );
  NOR3BX1 U12044 ( .AN(n24988), .B(n6532), .C(n24987), .Y(n6527) );
  NAND2BXL U12045 ( .AN(n24704), .B(n12342), .Y(n6531) );
  NAND2X1 U12046 ( .A(n5814), .B(n5815), .Y(n24988) );
  NAND2X1 U12047 ( .A(n25018), .B(n8033), .Y(n25008) );
  XOR2X4 U12048 ( .A(n6533), .B(n9087), .Y(n24642) );
  XOR2X4 U12049 ( .A(n6534), .B(n9083), .Y(n24662) );
  AOI21X2 U12050 ( .A0(n7738), .A1(n5793), .B0(n9079), .Y(n6534) );
  INVX2 U12051 ( .A(n6535), .Y(n13141) );
  NAND2X4 U12052 ( .A(n6817), .B(n6790), .Y(n6535) );
  AOI21X2 U12053 ( .A0(n6535), .A1(n5886), .B0(n6789), .Y(n6750) );
  INVX1 U12054 ( .A(n23982), .Y(n18596) );
  NAND2X1 U12055 ( .A(n6761), .B(n5847), .Y(n21949) );
  NAND2X1 U12056 ( .A(n13186), .B(n13184), .Y(n6536) );
  NOR2X1 U12057 ( .A(n21980), .B(n14568), .Y(n6538) );
  NAND3X1 U12058 ( .A(n22022), .B(n21979), .C(n14569), .Y(n6539) );
  NAND2BX4 U12059 ( .AN(n14545), .B(n7152), .Y(n22022) );
  NAND2X1 U12060 ( .A(n21978), .B(n14569), .Y(n6540) );
  NAND2X1 U12061 ( .A(n18549), .B(n18548), .Y(n18592) );
  NAND2X1 U12062 ( .A(n9946), .B(n6541), .Y(n10345) );
  INVX1 U12063 ( .A(n9945), .Y(n6541) );
  NOR2X2 U12064 ( .A(n10303), .B(n6542), .Y(n10299) );
  AOI21X2 U12065 ( .A0(n12625), .A1(n12624), .B0(n6543), .Y(n6811) );
  OAI21X1 U12066 ( .A0(n12623), .A1(n12622), .B0(n12621), .Y(n6543) );
  NAND2X1 U12067 ( .A(n12597), .B(n12598), .Y(n12621) );
  NAND2X1 U12068 ( .A(n12592), .B(n12593), .Y(n12622) );
  OAI21X1 U12069 ( .A0(n12602), .A1(n12608), .B0(n12603), .Y(n12624) );
  NAND2X1 U12070 ( .A(n12590), .B(n12591), .Y(n12603) );
  NAND2X1 U12071 ( .A(n12589), .B(n12588), .Y(n12608) );
  NOR2X2 U12072 ( .A(n12591), .B(n12590), .Y(n12602) );
  NOR2X2 U12073 ( .A(n12623), .B(n12618), .Y(n12625) );
  NOR2X2 U12074 ( .A(n12593), .B(n12592), .Y(n12618) );
  NAND2BX1 U12075 ( .AN(n24874), .B(n5860), .Y(n6544) );
  NAND2X1 U12076 ( .A(n13996), .B(n13526), .Y(n6545) );
  NAND3X2 U12077 ( .A(n24917), .B(n13526), .C(n13997), .Y(n6546) );
  NAND2BX1 U12078 ( .AN(n22931), .B(n24664), .Y(n23009) );
  NAND2XL U12079 ( .A(n6548), .B(U2_A_r_d[6]), .Y(n24954) );
  INVX1 U12080 ( .A(n14066), .Y(n6548) );
  NOR2XL U12081 ( .A(n14066), .B(U2_A_r_d[6]), .Y(n24547) );
  NOR2X1 U12082 ( .A(n14066), .B(U2_A_i_d[6]), .Y(n22848) );
  AND2X2 U12083 ( .A(n14066), .B(n5776), .Y(n24953) );
  AND2X1 U12084 ( .A(n14066), .B(n5773), .Y(n22558) );
  AOI2BB1X2 U12085 ( .A0N(n13312), .A1N(n6549), .B0(n13313), .Y(n13375) );
  NOR2BX2 U12086 ( .AN(n13302), .B(n6550), .Y(n13312) );
  NOR2X1 U12087 ( .A(n5903), .B(n13303), .Y(n6550) );
  NAND2X1 U12088 ( .A(n24917), .B(n13997), .Y(n6551) );
  XOR2X2 U12089 ( .A(n10546), .B(n10545), .Y(U1_U0_z0[23]) );
  NAND2X2 U12090 ( .A(n7051), .B(BOPB[28]), .Y(n10687) );
  INVX1 U12091 ( .A(n10644), .Y(n6554) );
  NOR2X2 U12092 ( .A(n6555), .B(n10645), .Y(n6867) );
  NOR2X1 U12093 ( .A(n10644), .B(n6556), .Y(n6555) );
  INVX1 U12094 ( .A(n10646), .Y(n6556) );
  XOR2X1 U12095 ( .A(n10663), .B(n10644), .Y(U1_U0_z0[4]) );
  NOR2X2 U12096 ( .A(n8204), .B(AOPD[36]), .Y(n10970) );
  NAND2X4 U12097 ( .A(n6559), .B(n6557), .Y(n10957) );
  NOR2X4 U12098 ( .A(n6558), .B(n6560), .Y(n6557) );
  NOR2X2 U12099 ( .A(n10983), .B(n10974), .Y(n6558) );
  NAND2X4 U12100 ( .A(n8320), .B(n10980), .Y(n6559) );
  OAI21X4 U12101 ( .A0(n10989), .A1(n10995), .B0(n10990), .Y(n10980) );
  INVX1 U12102 ( .A(n10957), .Y(n10965) );
  NAND2X2 U12103 ( .A(n8204), .B(AOPD[36]), .Y(n10983) );
  NAND2X1 U12104 ( .A(n8060), .B(AOPD[35]), .Y(n10990) );
  NAND2X2 U12105 ( .A(n8063), .B(AOPD[34]), .Y(n10995) );
  NAND2X1 U12106 ( .A(W2[9]), .B(W2[25]), .Y(n9893) );
  AOI21X2 U12107 ( .A0(n22466), .A1(n22464), .B0(n22455), .Y(n22461) );
  OAI21X4 U12108 ( .A0(n22471), .A1(n22468), .B0(n22469), .Y(n22466) );
  AOI21X4 U12109 ( .A0(n22473), .A1(n7285), .B0(n6563), .Y(n22471) );
  NAND2X1 U12110 ( .A(n7611), .B(n22477), .Y(n6563) );
  NAND2X2 U12111 ( .A(n22444), .B(n6564), .Y(n22473) );
  NAND2BX2 U12112 ( .AN(n22445), .B(n5854), .Y(n6564) );
  NAND2X1 U12113 ( .A(n8322), .B(n10946), .Y(n8324) );
  NOR2X1 U12114 ( .A(n7989), .B(AOPD[39]), .Y(n10960) );
  NOR2X1 U12115 ( .A(n8199), .B(AOPD[38]), .Y(n10954) );
  NOR2X1 U12116 ( .A(n10940), .B(n10949), .Y(n8322) );
  NOR2X1 U12117 ( .A(n8196), .B(AOPD[41]), .Y(n10940) );
  AOI21X4 U12118 ( .A0(n13382), .A1(n6565), .B0(n7572), .Y(n13400) );
  OAI21X4 U12119 ( .A0(n13370), .A1(n13366), .B0(n13367), .Y(n13382) );
  NAND2X2 U12120 ( .A(n13259), .B(n13260), .Y(n13370) );
  NOR2X2 U12121 ( .A(n13384), .B(n13388), .Y(n6565) );
  NOR2X2 U12122 ( .A(n6911), .B(n13262), .Y(n13388) );
  NOR2X1 U12123 ( .A(n13259), .B(n13260), .Y(n13364) );
  AND2X2 U12124 ( .A(U1_U0_y2[32]), .B(U1_U0_y0[32]), .Y(n8443) );
  XOR2X2 U12125 ( .A(U1_U0_y2[32]), .B(U1_U0_y0[32]), .Y(n8440) );
  NOR2X1 U12126 ( .A(n6567), .B(n6566), .Y(n19789) );
  NOR2X1 U12127 ( .A(n6649), .B(n19793), .Y(n6567) );
  CLKINVX3 U12128 ( .A(n6568), .Y(n8449) );
  NAND3X1 U12129 ( .A(n8446), .B(n5890), .C(n8588), .Y(n6568) );
  CLKINVX3 U12130 ( .A(n6666), .Y(n6643) );
  NAND3X2 U12131 ( .A(n8449), .B(n8542), .C(n8586), .Y(n6666) );
  NAND2X4 U12132 ( .A(n8541), .B(n8429), .Y(n8563) );
  NOR2X4 U12133 ( .A(n8543), .B(n8548), .Y(n8429) );
  NOR2X4 U12134 ( .A(n8427), .B(n8428), .Y(n8543) );
  NAND2X4 U12135 ( .A(n7531), .B(n8564), .Y(n7400) );
  NOR2X4 U12136 ( .A(n8568), .B(n8570), .Y(n7531) );
  NOR2X4 U12137 ( .A(n8436), .B(n8437), .Y(n8570) );
  NOR2X4 U12138 ( .A(n8435), .B(n8434), .Y(n8568) );
  NAND2X1 U12139 ( .A(n19767), .B(n5782), .Y(n16665) );
  XOR2X2 U12140 ( .A(n8595), .B(n8594), .Y(n19767) );
  NAND3X1 U12141 ( .A(n6572), .B(n6570), .C(n6569), .Y(n5094) );
  NAND2BXL U12142 ( .AN(U1_pipe4[26]), .B(n6578), .Y(n6569) );
  NAND3X1 U12143 ( .A(n6634), .B(n6635), .C(n6571), .Y(n6570) );
  NAND2X1 U12144 ( .A(n6575), .B(n6577), .Y(n6635) );
  NOR2X1 U12145 ( .A(n6574), .B(n6578), .Y(n6573) );
  INVX1 U12146 ( .A(n6575), .Y(n6574) );
  AOI21X2 U12147 ( .A0(n7536), .A1(n16629), .B0(n6576), .Y(n6575) );
  NAND2X1 U12148 ( .A(n7533), .B(n16629), .Y(n6577) );
  INVXL U12149 ( .A(n17187), .Y(n6578) );
  OAI21X1 U12150 ( .A0(n8514), .A1(n8463), .B0(n8462), .Y(n8475) );
  AOI21X2 U12151 ( .A0(n8479), .A1(n6592), .B0(n6581), .Y(n8462) );
  NOR2X2 U12152 ( .A(n8412), .B(n8411), .Y(n8484) );
  NOR2X1 U12153 ( .A(n8513), .B(n8515), .Y(n8478) );
  NOR2X1 U12154 ( .A(n8408), .B(n8407), .Y(n8515) );
  OAI21XL U12155 ( .A0(n17024), .A1(n6583), .B0(n16748), .Y(n17019) );
  OAI21XL U12156 ( .A0(n8472), .A1(n8468), .B0(n8469), .Y(n6584) );
  OAI22X1 U12157 ( .A0(n6589), .A1(n6587), .B0(n5816), .B1(U1_A_r_d0[25]), .Y(
        n12335) );
  XOR2X2 U12158 ( .A(n6589), .B(n6588), .Y(n20188) );
  XNOR2X1 U12159 ( .A(n5851), .B(n29007), .Y(n6588) );
  AOI21X4 U12160 ( .A0(n20190), .A1(n12333), .B0(n6590), .Y(n6589) );
  INVX1 U12161 ( .A(n19791), .Y(n6590) );
  NAND3X2 U12162 ( .A(n6630), .B(n7303), .C(n19798), .Y(n20190) );
  OAI21X1 U12163 ( .A0(n8514), .A1(n8463), .B0(n8462), .Y(n6638) );
  NAND2X1 U12164 ( .A(n8516), .B(n6591), .Y(n8479) );
  OR2X2 U12165 ( .A(n8515), .B(n8512), .Y(n6591) );
  NOR2X2 U12166 ( .A(n8482), .B(n8484), .Y(n6592) );
  NOR2X1 U12167 ( .A(n8410), .B(n8409), .Y(n8482) );
  XOR2X2 U12168 ( .A(n6593), .B(n8546), .Y(n19745) );
  OAI21X1 U12169 ( .A0(n8552), .A1(n8548), .B0(n8549), .Y(n6593) );
  AOI21X4 U12170 ( .A0(n8542), .A1(n8541), .B0(n8540), .Y(n8552) );
  AOI21X1 U12171 ( .A0(n8680), .A1(n16655), .B0(n8679), .Y(n6676) );
  OR2X2 U12172 ( .A(n8674), .B(n16679), .Y(n6594) );
  AOI21X4 U12173 ( .A0(n8575), .A1(n8564), .B0(n7544), .Y(n8569) );
  NAND2X2 U12174 ( .A(n8542), .B(n6596), .Y(n6595) );
  CLKINVX3 U12175 ( .A(n8563), .Y(n6596) );
  NAND2X4 U12176 ( .A(n6608), .B(n6607), .Y(n8542) );
  NAND2X1 U12177 ( .A(n19751), .B(n7069), .Y(n8672) );
  NAND2X1 U12178 ( .A(n16633), .B(n16640), .Y(n6601) );
  XOR2X1 U12179 ( .A(n7165), .B(n7166), .Y(n7141) );
  OAI21X4 U12180 ( .A0(n7400), .A1(n8562), .B0(n6603), .Y(n8585) );
  OAI21X2 U12181 ( .A0(n8567), .A1(n8570), .B0(n8571), .Y(n6604) );
  NAND2X2 U12182 ( .A(n8434), .B(n8435), .Y(n8567) );
  AOI21X4 U12183 ( .A0(n8540), .A1(n8429), .B0(n6605), .Y(n8562) );
  OAI21X2 U12184 ( .A0(n8543), .A1(n8549), .B0(n8544), .Y(n6605) );
  OAI21X4 U12185 ( .A0(n8527), .A1(n8531), .B0(n8528), .Y(n8540) );
  NAND2X2 U12186 ( .A(n8421), .B(n8422), .Y(n8531) );
  INVX1 U12187 ( .A(n8675), .Y(n7301) );
  OAI21X2 U12188 ( .A0(n8595), .A1(n8592), .B0(n6665), .Y(n6606) );
  AOI21X4 U12189 ( .A0(n6633), .A1(n8588), .B0(n8587), .Y(n8595) );
  CLKINVX3 U12190 ( .A(n19777), .Y(n19773) );
  AOI21X1 U12191 ( .A0(n8629), .A1(n8148), .B0(n8628), .Y(n16945) );
  NAND2X1 U12192 ( .A(n19777), .B(n5757), .Y(n8148) );
  XOR2X4 U12193 ( .A(n7162), .B(n8625), .Y(n19777) );
  AOI21X1 U12194 ( .A0(n8542), .A1(n5899), .B0(n8526), .Y(n8530) );
  NAND3X2 U12195 ( .A(n6638), .B(n6637), .C(n8474), .Y(n6607) );
  AOI21X4 U12196 ( .A0(n8473), .A1(n6637), .B0(n6636), .Y(n6608) );
  NAND2X1 U12197 ( .A(n8419), .B(n8420), .Y(n8537) );
  OAI21XL U12198 ( .A0(n6665), .A1(n8589), .B0(n8590), .Y(n6612) );
  AOI21X2 U12199 ( .A0(n8446), .A1(n8587), .B0(n6612), .Y(n8619) );
  OAI21X4 U12200 ( .A0(n8596), .A1(n8602), .B0(n8597), .Y(n8587) );
  NOR2X2 U12201 ( .A(n8448), .B(n8447), .Y(n8621) );
  XOR2X1 U12202 ( .A(n6614), .B(n16940), .Y(n6613) );
  NOR2X1 U12203 ( .A(n7533), .B(n7536), .Y(n6614) );
  NAND2X2 U12204 ( .A(n8430), .B(n8431), .Y(n8582) );
  INVX1 U12205 ( .A(n19765), .Y(n19756) );
  NAND2X1 U12206 ( .A(n19765), .B(n5783), .Y(n16674) );
  XOR2X2 U12207 ( .A(n6633), .B(n8604), .Y(n19765) );
  NOR2X4 U12208 ( .A(n8440), .B(n8441), .Y(n8596) );
  XOR2X2 U12209 ( .A(n6616), .B(n6615), .Y(n19775) );
  NOR2BX1 U12210 ( .AN(n8627), .B(n8626), .Y(n6615) );
  NAND2X1 U12211 ( .A(n6648), .B(n6646), .Y(n6616) );
  NOR2X1 U12212 ( .A(n6617), .B(U1_A_r_d0[19]), .Y(n20216) );
  NAND2XL U12213 ( .A(n6617), .B(U1_A_i_d0[19]), .Y(n16961) );
  NAND2X1 U12214 ( .A(n6617), .B(U1_A_r_d0[19]), .Y(n20215) );
  NAND3X1 U12215 ( .A(n6627), .B(n6624), .C(n6618), .Y(n4721) );
  AOI2BB1XL U12216 ( .A0N(n7527), .A1N(n6622), .B0(n6619), .Y(n6618) );
  NOR2XL U12217 ( .A(n19787), .B(n5928), .Y(n6621) );
  NAND2XL U12218 ( .A(n6623), .B(n19788), .Y(n6622) );
  NOR2XL U12219 ( .A(n7527), .B(n6626), .Y(n6625) );
  NAND2X1 U12220 ( .A(n5810), .B(n19787), .Y(n6626) );
  OR2X2 U12221 ( .A(n19793), .B(n6628), .Y(n6627) );
  NAND2XL U12222 ( .A(n7527), .B(n6629), .Y(n6628) );
  NOR2XL U12223 ( .A(n19788), .B(n5928), .Y(n6629) );
  NAND2BX2 U12224 ( .AN(n12324), .B(n6631), .Y(n20194) );
  NOR2BXL U12225 ( .AN(n20210), .B(n20208), .Y(n6632) );
  OAI21X1 U12226 ( .A0(n6632), .A1(n20209), .B0(n12325), .Y(n6631) );
  NAND2X4 U12227 ( .A(n7398), .B(n7399), .Y(n6633) );
  XOR2X1 U12228 ( .A(n5851), .B(n29008), .Y(n6634) );
  OAI21X2 U12229 ( .A0(n8536), .A1(n8533), .B0(n8537), .Y(n6636) );
  NOR2X1 U12230 ( .A(n8468), .B(n8464), .Y(n8474) );
  NOR2X4 U12231 ( .A(n8536), .B(n8534), .Y(n6637) );
  INVX1 U12232 ( .A(n12313), .Y(n19760) );
  NAND2X1 U12233 ( .A(n12313), .B(U1_A_i_d0[15]), .Y(n16979) );
  NAND2X1 U12234 ( .A(n6639), .B(n8627), .Y(n8634) );
  NAND2X1 U12235 ( .A(n6648), .B(n6644), .Y(n6639) );
  NAND2X1 U12236 ( .A(n6667), .B(n6666), .Y(n7162) );
  NAND2XL U12237 ( .A(n7526), .B(n6650), .Y(n6649) );
  AOI2BB1XL U12238 ( .A0N(n19752), .A1N(n19851), .B0(n19762), .Y(n6651) );
  NAND2X1 U12239 ( .A(n6659), .B(n6660), .Y(n6652) );
  NAND3X1 U12240 ( .A(n6664), .B(n19770), .C(n6653), .Y(n6663) );
  NAND2X1 U12241 ( .A(n8402), .B(n8495), .Y(n8404) );
  NOR2X1 U12242 ( .A(n8503), .B(n8498), .Y(n8402) );
  NAND2X1 U12243 ( .A(n8399), .B(n8385), .Y(n8498) );
  NOR2X1 U12244 ( .A(n8400), .B(U1_U0_y2[13]), .Y(n8503) );
  AOI21X1 U12245 ( .A0(n8575), .A1(n5900), .B0(n6656), .Y(n6655) );
  XOR2X2 U12246 ( .A(U1_U0_y0[21]), .B(U1_U0_y2[21]), .Y(n8417) );
  NAND3X1 U12247 ( .A(n19870), .B(n19772), .C(n19823), .Y(n6660) );
  NOR2X1 U12248 ( .A(n19771), .B(n19825), .Y(n19772) );
  NAND2X1 U12249 ( .A(n6657), .B(n8683), .Y(n16641) );
  NOR2X1 U12250 ( .A(n19784), .B(n19796), .Y(n19785) );
  NAND2X1 U12251 ( .A(n19802), .B(n19781), .Y(n19796) );
  NAND2BX1 U12252 ( .AN(n19775), .B(n7074), .Y(n19781) );
  NOR2X1 U12253 ( .A(n19779), .B(n19812), .Y(n19802) );
  NOR2X1 U12254 ( .A(n19777), .B(U1_A_r_d0[22]), .Y(n19779) );
  NAND2X1 U12255 ( .A(n8426), .B(n8425), .Y(n8549) );
  OAI21X1 U12256 ( .A0(n19795), .A1(n19784), .B0(n19783), .Y(n6658) );
  NAND2BX2 U12257 ( .AN(n6663), .B(n6660), .Y(n6661) );
  NAND2X1 U12258 ( .A(n6662), .B(n19778), .Y(n19803) );
  OR2X2 U12259 ( .A(n19779), .B(n19811), .Y(n6662) );
  OR2X2 U12260 ( .A(n19771), .B(n19824), .Y(n6664) );
  OR2X2 U12261 ( .A(n8675), .B(U1_A_r_d0[20]), .Y(n19769) );
  NAND2X1 U12262 ( .A(n16628), .B(n16629), .Y(n16940) );
  NOR2X4 U12263 ( .A(n8527), .B(n8525), .Y(n8541) );
  NOR2X2 U12264 ( .A(n8421), .B(n8422), .Y(n8525) );
  NOR2X4 U12265 ( .A(n8423), .B(n8424), .Y(n8527) );
  NAND2X1 U12266 ( .A(n8436), .B(n8437), .Y(n8571) );
  NOR2BX4 U12267 ( .AN(U1_U0_y2[29]), .B(n6670), .Y(n8437) );
  INVXL U12268 ( .A(n6888), .Y(n6671) );
  XOR2X1 U12269 ( .A(n6673), .B(n16649), .Y(n6672) );
  AOI21X1 U12270 ( .A0(n16633), .A1(n6674), .B0(n16646), .Y(n6673) );
  NAND2X1 U12271 ( .A(n8414), .B(n8413), .Y(n8469) );
  NOR2X2 U12272 ( .A(n8416), .B(n8415), .Y(n8464) );
  CLKINVX3 U12273 ( .A(n6661), .Y(n19820) );
  NAND2X1 U12274 ( .A(n6661), .B(n19802), .Y(n6677) );
  OAI21X2 U12275 ( .A0(n8569), .A1(n8568), .B0(n8567), .Y(n6678) );
  NOR2X2 U12276 ( .A(n8404), .B(n8493), .Y(n6679) );
  NOR2X1 U12277 ( .A(n13964), .B(n13965), .Y(n13963) );
  NOR2X1 U12278 ( .A(n20317), .B(n20316), .Y(n6680) );
  AOI21X2 U12279 ( .A0(n14971), .A1(n7470), .B0(n6683), .Y(n16785) );
  NOR2X1 U12280 ( .A(n16785), .B(n16781), .Y(n7487) );
  NOR2X1 U12281 ( .A(n11295), .B(n6686), .Y(n6685) );
  NOR2BXL U12282 ( .AN(n11293), .B(n11321), .Y(n6686) );
  AOI21X2 U12283 ( .A0(n7448), .A1(n12904), .B0(n6687), .Y(n7447) );
  OAI21X1 U12284 ( .A0(n12927), .A1(n12930), .B0(n12931), .Y(n6687) );
  NAND2X1 U12285 ( .A(n12792), .B(n12791), .Y(n12927) );
  OAI21X1 U12286 ( .A0(n12789), .A1(n12788), .B0(n12787), .Y(n12904) );
  NAND2X1 U12287 ( .A(n12766), .B(n12767), .Y(n12787) );
  NOR2X1 U12288 ( .A(n12766), .B(n12767), .Y(n12789) );
  NOR2X2 U12289 ( .A(n12903), .B(n12902), .Y(n12930) );
  NOR2X2 U12290 ( .A(n12792), .B(n12791), .Y(n12928) );
  AOI21X1 U12291 ( .A0(n19870), .A1(n19823), .B0(n19822), .Y(n19835) );
  OAI21X1 U12292 ( .A0(n8535), .A1(n8534), .B0(n8533), .Y(n6689) );
  NOR2X2 U12293 ( .A(n6690), .B(n8473), .Y(n8535) );
  AND2X2 U12294 ( .A(n8475), .B(n8474), .Y(n6690) );
  NOR2BX1 U12295 ( .AN(U1_U0_y0[13]), .B(U1_U0_y2[13]), .Y(n6691) );
  NOR2X1 U12296 ( .A(n14963), .B(n5850), .Y(n14965) );
  AND2X2 U12297 ( .A(n13969), .B(n13967), .Y(n6692) );
  OAI2BB1X4 U12298 ( .A0N(n13048), .A1N(n7172), .B0(n13047), .Y(n13019) );
  NOR2BX2 U12299 ( .AN(n14770), .B(n6694), .Y(n6693) );
  NOR2X1 U12300 ( .A(n14766), .B(n14769), .Y(n6694) );
  NAND3X2 U12301 ( .A(n6696), .B(n14703), .C(n7797), .Y(n6695) );
  NAND2X1 U12302 ( .A(n7310), .B(n7309), .Y(n6696) );
  NAND3X2 U12303 ( .A(n7800), .B(n7796), .C(n7795), .Y(n7310) );
  NOR2X1 U12304 ( .A(n7062), .B(AOPC[38]), .Y(n11310) );
  XOR2X4 U12305 ( .A(n9884), .B(n5759), .Y(U1_U2_z2[13]) );
  XOR2X1 U12306 ( .A(n22183), .B(n6697), .Y(n22184) );
  NOR2X4 U12307 ( .A(n14225), .B(n14224), .Y(n14361) );
  OAI21X4 U12308 ( .A0(n10661), .A1(n10656), .B0(n10657), .Y(n10645) );
  NOR2X2 U12309 ( .A(n8126), .B(BOPB[31]), .Y(n10656) );
  NAND2X1 U12310 ( .A(n8132), .B(BOPB[30]), .Y(n10661) );
  AOI21X1 U12311 ( .A0(n7708), .A1(n6699), .B0(n6698), .Y(n22178) );
  NOR2XL U12312 ( .A(n7707), .B(U2_A_i_d[25]), .Y(n6698) );
  NAND2X2 U12313 ( .A(n7709), .B(n22176), .Y(n7708) );
  AOI21X1 U12314 ( .A0(n10260), .A1(n10231), .B0(n10230), .Y(n6701) );
  NAND2BX1 U12315 ( .AN(n10232), .B(n10230), .Y(n6700) );
  XOR2X2 U12316 ( .A(n6701), .B(n10237), .Y(U1_U1_z1[6]) );
  OAI21XL U12317 ( .A0(n13953), .A1(n13952), .B0(n13951), .Y(n7473) );
  NAND2X1 U12318 ( .A(n13928), .B(n13929), .Y(n13952) );
  NOR2X1 U12319 ( .A(n13931), .B(n13930), .Y(n13953) );
  AOI21X1 U12320 ( .A0(n13970), .A1(n13969), .B0(n13968), .Y(n13977) );
  OAI21X2 U12321 ( .A0(n12919), .A1(n12922), .B0(n12923), .Y(n7828) );
  NAND2X1 U12322 ( .A(n12782), .B(n12783), .Y(n12919) );
  NOR2BXL U12323 ( .AN(n17355), .B(n17358), .Y(n7517) );
  NAND2X1 U12324 ( .A(n5866), .B(n13037), .Y(n17355) );
  INVXL U12325 ( .A(n7826), .Y(n7521) );
  NOR2X2 U12326 ( .A(n7522), .B(n7825), .Y(n6703) );
  NAND2BX1 U12327 ( .AN(n17596), .B(n7932), .Y(n6704) );
  NAND2X1 U12328 ( .A(n6706), .B(n17602), .Y(n6705) );
  NOR2BX2 U12329 ( .AN(n7829), .B(n17596), .Y(n6706) );
  MXI2X1 U12330 ( .A(n6707), .B(U1_pipe11[26]), .S0(n6708), .Y(n4892) );
  AOI21XL U12331 ( .A0(n17602), .A1(n7829), .B0(n7932), .Y(n17600) );
  INVXL U12332 ( .A(n5812), .Y(n6708) );
  CLKINVX3 U12333 ( .A(n13035), .Y(n14950) );
  NAND2XL U12334 ( .A(n19541), .B(n13035), .Y(n17662) );
  CLKINVX3 U12335 ( .A(n20014), .Y(n19996) );
  INVX1 U12336 ( .A(n7433), .Y(n6710) );
  NAND2X4 U12337 ( .A(W1[17]), .B(W1[1]), .Y(n10003) );
  NAND2X1 U12338 ( .A(n8190), .B(BOPB[36]), .Y(n10630) );
  AOI21X4 U12339 ( .A0(n6713), .A1(n7934), .B0(n6711), .Y(n7148) );
  OAI21X2 U12340 ( .A0(n10616), .A1(n9559), .B0(n9558), .Y(n6711) );
  OAI21X4 U12341 ( .A0(n10644), .A1(n7568), .B0(n7566), .Y(n7934) );
  BUFX8 U12342 ( .A(n7148), .Y(n6712) );
  OAI21X1 U12343 ( .A0(n6712), .A1(n10592), .B0(n10593), .Y(n10591) );
  NOR2X2 U12344 ( .A(n9559), .B(n10617), .Y(n6713) );
  INVX8 U12345 ( .A(n6714), .Y(U1_U1_z2[9]) );
  NAND2X4 U12346 ( .A(n5770), .B(n9991), .Y(n7395) );
  XNOR2X4 U12347 ( .A(n6715), .B(n10227), .Y(n6714) );
  AOI21X4 U12348 ( .A0(n7397), .A1(n9981), .B0(n9962), .Y(n6715) );
  AOI21X4 U12349 ( .A0(n7393), .A1(n9966), .B0(n7392), .Y(n7396) );
  NAND2X1 U12350 ( .A(n7454), .B(n16837), .Y(n16808) );
  NOR2X1 U12351 ( .A(n9384), .B(n9389), .Y(n9288) );
  NAND2X1 U12352 ( .A(n9286), .B(n9270), .Y(n9384) );
  NAND2X1 U12353 ( .A(n14950), .B(n20002), .Y(n16853) );
  XOR2X1 U12354 ( .A(n7863), .B(n7814), .Y(n7938) );
  NOR2X1 U12355 ( .A(n13972), .B(n13971), .Y(n13976) );
  NOR2X1 U12356 ( .A(n13957), .B(n13956), .Y(n13962) );
  MXI2X1 U12357 ( .A(n6717), .B(U1_pipe13[27]), .S0(n5811), .Y(n4750) );
  NOR2XL U12358 ( .A(n5843), .B(n7814), .Y(n6718) );
  AND2X2 U12359 ( .A(n13982), .B(n13980), .Y(n6720) );
  NAND2BX1 U12360 ( .AN(n13979), .B(n6721), .Y(n13982) );
  NOR2X1 U12361 ( .A(n6724), .B(n6723), .Y(n6722) );
  NOR2BX1 U12362 ( .AN(n13968), .B(n13976), .Y(n6724) );
  NAND2X1 U12363 ( .A(n13970), .B(n7474), .Y(n6725) );
  AOI21X4 U12364 ( .A0(n6726), .A1(n10129), .B0(n10128), .Y(n10177) );
  AOI21X1 U12365 ( .A0(n6726), .A1(n10136), .B0(n10135), .Y(n6862) );
  AOI21X2 U12366 ( .A0(n7580), .A1(n6726), .B0(n7579), .Y(n7273) );
  XNOR2X1 U12367 ( .A(n10165), .B(n6726), .Y(U0_U0_z1[8]) );
  OAI2BB1X2 U12368 ( .A0N(n10186), .A1N(n6726), .B0(n7362), .Y(n7766) );
  OAI21X4 U12369 ( .A0(n10139), .A1(n6864), .B0(n6863), .Y(n6726) );
  NOR2X1 U12370 ( .A(n14215), .B(n14216), .Y(n14298) );
  NAND2X1 U12371 ( .A(n25174), .B(n5780), .Y(n21783) );
  XOR2X4 U12372 ( .A(n6729), .B(n14437), .Y(n25174) );
  NOR2X1 U12373 ( .A(n13959), .B(n13962), .Y(n7453) );
  NAND2X1 U12374 ( .A(n13955), .B(n13950), .Y(n13959) );
  NOR2X2 U12375 ( .A(n13934), .B(n13938), .Y(n13950) );
  NOR2X2 U12376 ( .A(n13926), .B(n13927), .Y(n13934) );
  NOR2X1 U12377 ( .A(n13953), .B(n13949), .Y(n13955) );
  NOR2X1 U12378 ( .A(n13928), .B(n13929), .Y(n13949) );
  OAI22X4 U12379 ( .A0(n6731), .A1(n13429), .B0(n13430), .B1(n13431), .Y(
        n13441) );
  OAI21X4 U12380 ( .A0(n13400), .A1(n7283), .B0(n7282), .Y(n13429) );
  NAND2X2 U12381 ( .A(n13428), .B(n6732), .Y(n6731) );
  INVX1 U12382 ( .A(n13430), .Y(n6732) );
  NAND2X4 U12383 ( .A(n13426), .B(n13427), .Y(n13428) );
  NOR2X4 U12384 ( .A(n13401), .B(n7283), .Y(n13426) );
  XOR2X2 U12385 ( .A(U0_U0_y1[24]), .B(U0_U0_y0[24]), .Y(n13261) );
  OAI21X4 U12386 ( .A0(n10196), .A1(n10257), .B0(n10195), .Y(n10230) );
  NOR2X4 U12387 ( .A(n7996), .B(W1[19]), .Y(n6736) );
  OAI2BB2X4 U12388 ( .B0(n12005), .B1(n6737), .A0N(n8040), .A1N(W1[17]), .Y(
        n6820) );
  NOR2X4 U12389 ( .A(n8009), .B(W1[16]), .Y(n12005) );
  NAND2X1 U12390 ( .A(n12477), .B(n12478), .Y(n12552) );
  XOR2X1 U12391 ( .A(n6738), .B(n22298), .Y(n22299) );
  OAI21XL U12392 ( .A0(n22301), .A1(n21955), .B0(n21956), .Y(n6738) );
  AOI21X4 U12393 ( .A0(n22303), .A1(n13171), .B0(n13170), .Y(n22301) );
  NAND3X2 U12394 ( .A(n6747), .B(n6746), .C(n6739), .Y(n22303) );
  XOR2X2 U12395 ( .A(n6740), .B(n6971), .Y(n7346) );
  AOI21X1 U12396 ( .A0(n12601), .A1(n12619), .B0(n12624), .Y(n12596) );
  OAI21X1 U12397 ( .A0(n13154), .A1(n12620), .B0(n12627), .Y(n12601) );
  OAI21X2 U12398 ( .A0(n8993), .A1(n8992), .B0(n8991), .Y(n9017) );
  NAND2X1 U12399 ( .A(n8957), .B(n6741), .Y(n8991) );
  XNOR2X1 U12400 ( .A(U0_U2_y1[24]), .B(n6742), .Y(n6741) );
  NAND2X1 U12401 ( .A(n6988), .B(n22347), .Y(n6754) );
  AOI21X1 U12402 ( .A0(n22351), .A1(n22353), .B0(n13124), .Y(n22338) );
  NOR2X1 U12403 ( .A(n22935), .B(n13123), .Y(n6743) );
  AND2X2 U12404 ( .A(U0_U2_y2[29]), .B(U0_U2_y0[29]), .Y(n12188) );
  XOR2X2 U12405 ( .A(U0_U2_y0[29]), .B(U0_U2_y2[29]), .Y(n12185) );
  INVX4 U12406 ( .A(n12257), .Y(n6744) );
  INVX1 U12407 ( .A(n22303), .Y(n22315) );
  NAND3X1 U12408 ( .A(n22318), .B(n6748), .C(n22359), .Y(n6746) );
  NAND2BX4 U12409 ( .AN(n7425), .B(n7424), .Y(n22359) );
  NAND2X1 U12410 ( .A(n22317), .B(n6748), .Y(n6747) );
  NOR2X1 U12411 ( .A(n22319), .B(n7428), .Y(n6748) );
  NAND2BX1 U12412 ( .AN(n22932), .B(n14562), .Y(n21992) );
  XOR2X4 U12413 ( .A(n6749), .B(n12228), .Y(n14562) );
  OAI21X4 U12414 ( .A0(n12247), .A1(n12229), .B0(n12230), .Y(n6749) );
  OAI21X1 U12415 ( .A0(n12193), .A1(n12205), .B0(n12209), .Y(n6751) );
  XOR2X2 U12416 ( .A(U0_U2_y0[24]), .B(U0_U2_y2[24]), .Y(n12143) );
  NOR2X1 U12417 ( .A(n22331), .B(n22319), .Y(n6843) );
  AOI21X1 U12418 ( .A0(n13127), .A1(n6988), .B0(n13126), .Y(n6753) );
  NOR2X1 U12419 ( .A(n22337), .B(n6754), .Y(n22318) );
  NAND2X2 U12420 ( .A(n12160), .B(n6752), .Y(n12178) );
  NOR2X1 U12421 ( .A(n6758), .B(n21956), .Y(n6757) );
  NAND2BX1 U12422 ( .AN(n21955), .B(n21949), .Y(n6760) );
  NOR2X1 U12423 ( .A(n25654), .B(n5815), .Y(n25656) );
  NOR2X2 U12424 ( .A(n12182), .B(n12181), .Y(n12199) );
  NOR2X2 U12425 ( .A(n12183), .B(n12184), .Y(n12195) );
  NAND2X1 U12426 ( .A(n12052), .B(n12037), .Y(n6763) );
  NOR2X1 U12427 ( .A(n6763), .B(n12111), .Y(n12055) );
  NAND2X2 U12428 ( .A(n6782), .B(n6764), .Y(n14564) );
  OAI21X1 U12429 ( .A0(n7248), .A1(n5874), .B0(n6765), .Y(n6764) );
  OAI2BB1X1 U12430 ( .A0N(n12222), .A1N(n7245), .B0(n7248), .Y(n6765) );
  NAND2BX1 U12431 ( .AN(n22930), .B(n14564), .Y(n6934) );
  XOR2X2 U12432 ( .A(n6766), .B(n6923), .Y(n22930) );
  NOR2X1 U12433 ( .A(n24586), .B(n13103), .Y(n25427) );
  AOI21X1 U12434 ( .A0(n12101), .A1(n12099), .B0(n12093), .Y(n6768) );
  OAI21X1 U12435 ( .A0(n12122), .A1(n12091), .B0(n12090), .Y(n12101) );
  XOR2X2 U12436 ( .A(n6769), .B(n6893), .Y(n14532) );
  OAI21X4 U12437 ( .A0(n12166), .A1(n12176), .B0(n12178), .Y(n6769) );
  AOI2BB1X4 U12438 ( .A0N(n12258), .A1N(n6785), .B0(n12180), .Y(n12166) );
  AND2X2 U12439 ( .A(n25650), .B(n25652), .Y(n7006) );
  OR2X2 U12440 ( .A(n24692), .B(n14579), .Y(n25652) );
  NAND4X1 U12441 ( .A(n6779), .B(n6780), .C(n12239), .D(n6784), .Y(n25663) );
  NAND2X1 U12442 ( .A(n12071), .B(n12070), .Y(n12079) );
  NAND2X1 U12443 ( .A(n12068), .B(n12069), .Y(n12080) );
  NOR2X2 U12444 ( .A(n12071), .B(n12070), .Y(n12081) );
  XOR2X1 U12445 ( .A(U0_U1_y1[19]), .B(U0_U1_y0[19]), .Y(n8810) );
  AOI21X1 U12446 ( .A0(n8936), .A1(n8935), .B0(n8934), .Y(n6770) );
  OAI21X1 U12447 ( .A0(n9001), .A1(n9042), .B0(n9045), .Y(n8989) );
  AOI21X1 U12448 ( .A0(n9062), .A1(n9043), .B0(n9048), .Y(n9001) );
  NAND2BX4 U12449 ( .AN(n24638), .B(n6771), .Y(n24773) );
  NAND2X1 U12450 ( .A(n24639), .B(n24775), .Y(n6771) );
  INVX2 U12451 ( .A(n9093), .Y(n6773) );
  INVX1 U12452 ( .A(n9061), .Y(n6772) );
  NOR2X1 U12453 ( .A(n9061), .B(n9094), .Y(n9176) );
  INVX1 U12454 ( .A(n9094), .Y(n6774) );
  INVX1 U12455 ( .A(n24701), .Y(n24727) );
  NAND2BX2 U12456 ( .AN(n24673), .B(n24773), .Y(n6777) );
  INVX1 U12457 ( .A(n24744), .Y(n6778) );
  NAND2BX1 U12458 ( .AN(n24642), .B(n24662), .Y(n24744) );
  AND2X2 U12459 ( .A(U0_U1_y1[24]), .B(U0_U1_y0[24]), .Y(n8984) );
  NOR2X2 U12460 ( .A(n12215), .B(n12216), .Y(n12225) );
  NAND3BX2 U12461 ( .AN(n25677), .B(n12241), .C(n25679), .Y(n6779) );
  NAND2X1 U12462 ( .A(n25678), .B(n12241), .Y(n6780) );
  NAND2X1 U12463 ( .A(n12182), .B(n12181), .Y(n12200) );
  NAND2X1 U12464 ( .A(n25339), .B(n25343), .Y(n25680) );
  OR2X2 U12465 ( .A(n13128), .B(n24643), .Y(n25343) );
  XOR2X2 U12466 ( .A(n9169), .B(n9092), .Y(n24643) );
  NAND2BX1 U12467 ( .AN(n24642), .B(n14562), .Y(n25339) );
  NAND2X2 U12468 ( .A(n6781), .B(n12133), .Y(n6787) );
  NOR2X2 U12469 ( .A(n12151), .B(n12149), .Y(n6781) );
  NAND2X1 U12470 ( .A(n6783), .B(n14564), .Y(n25328) );
  INVX1 U12471 ( .A(n25663), .Y(n25675) );
  OR2X2 U12472 ( .A(n25681), .B(n12240), .Y(n6784) );
  NOR2X2 U12473 ( .A(n12240), .B(n25680), .Y(n12241) );
  NAND2X1 U12474 ( .A(n12183), .B(n12184), .Y(n12196) );
  NOR2X2 U12475 ( .A(n12135), .B(n12136), .Y(n12151) );
  NAND2BX1 U12476 ( .AN(n24645), .B(n14547), .Y(n25358) );
  NAND2BX1 U12477 ( .AN(n24644), .B(n13125), .Y(n25353) );
  NAND2BX2 U12478 ( .AN(n12156), .B(n5898), .Y(n6785) );
  NOR2X1 U12479 ( .A(n12393), .B(n25347), .Y(n25322) );
  NAND2X1 U12480 ( .A(n25364), .B(n12385), .Y(n25347) );
  NAND2X1 U12481 ( .A(n13123), .B(n5820), .Y(n25364) );
  NAND2X1 U12482 ( .A(n12084), .B(n12083), .Y(n12148) );
  NAND2BX1 U12483 ( .AN(n24619), .B(n14532), .Y(n25377) );
  INVX2 U12484 ( .A(n25320), .Y(n25370) );
  NOR2X1 U12485 ( .A(n12626), .B(n12620), .Y(n13148) );
  NAND2X1 U12486 ( .A(n12143), .B(n12144), .Y(n12157) );
  AOI21XL U12487 ( .A0(n13139), .A1(n5885), .B0(n6792), .Y(n6791) );
  INVXL U12488 ( .A(n13135), .Y(n6794) );
  AOI21X1 U12489 ( .A0(n6795), .A1(n22983), .B0(n22984), .Y(n6803) );
  NOR2X2 U12490 ( .A(n12477), .B(n12478), .Y(n12553) );
  NAND2X1 U12491 ( .A(n6799), .B(n6797), .Y(n6796) );
  XOR2X1 U12492 ( .A(n6799), .B(n6798), .Y(n7736) );
  INVX1 U12493 ( .A(n7209), .Y(n6800) );
  NOR2X1 U12494 ( .A(n22670), .B(n22672), .Y(n12575) );
  NOR2X1 U12495 ( .A(n7565), .B(n22913), .Y(n22672) );
  XOR2X4 U12496 ( .A(n6801), .B(n12548), .Y(n22913) );
  OAI2BB1X2 U12497 ( .A0N(n12549), .A1N(n12551), .B0(n12561), .Y(n6801) );
  NAND2X1 U12498 ( .A(n22916), .B(n6802), .Y(n23053) );
  INVX1 U12499 ( .A(n22913), .Y(n22922) );
  XOR2X1 U12500 ( .A(n6803), .B(n22987), .Y(n22988) );
  NAND2X1 U12501 ( .A(n13135), .B(n13140), .Y(n13147) );
  NOR2X2 U12502 ( .A(n12642), .B(n12641), .Y(n13134) );
  NAND2X1 U12503 ( .A(n25654), .B(n21946), .Y(n22295) );
  OAI21X1 U12504 ( .A0(n13188), .A1(n13187), .B0(n13186), .Y(n6804) );
  AOI2BB1X2 U12505 ( .A0N(n13151), .A1N(n13150), .B0(n6807), .Y(n6806) );
  INVX1 U12506 ( .A(n13149), .Y(n6807) );
  NAND2X1 U12507 ( .A(n13148), .B(n6810), .Y(n6809) );
  INVXL U12508 ( .A(n13154), .Y(n6810) );
  OAI22X1 U12509 ( .A0(n6814), .A1(n6812), .B0(n22884), .B1(n6815), .Y(n22971)
         );
  OAI2BB1XL U12510 ( .A0N(n22969), .A1N(n22970), .B0(n6813), .Y(n6812) );
  XOR2X1 U12511 ( .A(n5814), .B(n22972), .Y(n6816) );
  NOR2X2 U12512 ( .A(n8950), .B(n8949), .Y(n8967) );
  NAND2X1 U12513 ( .A(n13148), .B(n12551), .Y(n6817) );
  AOI21X4 U12514 ( .A0(n9017), .A1(n7180), .B0(n7179), .Y(n9099) );
  NOR2X1 U12515 ( .A(n8993), .B(n8990), .Y(n7726) );
  NAND2BX2 U12516 ( .AN(n7739), .B(n7181), .Y(n6818) );
  AOI21X2 U12517 ( .A0(n7183), .A1(n8952), .B0(n7182), .Y(n6819) );
  NAND2X1 U12518 ( .A(n12464), .B(n12465), .Y(n12474) );
  NAND2X1 U12519 ( .A(n6820), .B(n6827), .Y(n6826) );
  XNOR2X1 U12520 ( .A(n10265), .B(n6820), .Y(U1_U1_z1[2]) );
  INVX1 U12521 ( .A(n10255), .Y(n6821) );
  NAND2BX4 U12522 ( .AN(n10209), .B(n6825), .Y(n6856) );
  XNOR2X4 U12523 ( .A(n7403), .B(n6999), .Y(n6909) );
  OAI21X4 U12524 ( .A0(n9956), .A1(n9957), .B0(n6822), .Y(n7403) );
  NAND3X2 U12525 ( .A(n7395), .B(n7396), .C(n7394), .Y(n6822) );
  NAND2X1 U12526 ( .A(n10210), .B(n6823), .Y(n6825) );
  AOI21X2 U12527 ( .A0(n6823), .A1(n10217), .B0(n10216), .Y(n10246) );
  XOR2X1 U12528 ( .A(n6824), .B(n6823), .Y(U1_U1_z1[8]) );
  NOR2X4 U12529 ( .A(W1[5]), .B(W1[21]), .Y(n9974) );
  XOR2X4 U12530 ( .A(n6829), .B(n10261), .Y(U1_U1_z2[5]) );
  NAND2X1 U12531 ( .A(n6830), .B(n10007), .Y(n9979) );
  NAND2BX1 U12532 ( .AN(n10006), .B(n9976), .Y(n6830) );
  NAND2X4 U12533 ( .A(W1[16]), .B(W1[0]), .Y(n10005) );
  NOR2X4 U12534 ( .A(W1[17]), .B(W1[1]), .Y(n10002) );
  NOR2X4 U12535 ( .A(W1[19]), .B(W1[3]), .Y(n9977) );
  NOR2X1 U12536 ( .A(n7985), .B(W3[26]), .Y(n10077) );
  OAI21X2 U12537 ( .A0(n6831), .A1(n9938), .B0(n9939), .Y(n9889) );
  OAI21XL U12538 ( .A0(n7430), .A1(n22296), .B0(n22295), .Y(n6832) );
  NOR2X1 U12539 ( .A(n22931), .B(n14550), .Y(n22323) );
  XOR2X2 U12540 ( .A(n6833), .B(n12223), .Y(n14550) );
  AOI21X1 U12541 ( .A0(n12224), .A1(n12242), .B0(n12246), .Y(n6833) );
  AOI21X2 U12542 ( .A0(n9956), .A1(n9726), .B0(n6834), .Y(n9999) );
  NAND2X1 U12543 ( .A(W1[11]), .B(W1[27]), .Y(n9958) );
  NOR2X1 U12544 ( .A(n8015), .B(W3[23]), .Y(n6835) );
  OAI21X1 U12545 ( .A0(n6836), .A1(n10077), .B0(n10076), .Y(n10080) );
  XOR2X1 U12546 ( .A(n6836), .B(n10040), .Y(U2_U0_z1[10]) );
  AOI21X2 U12547 ( .A0(n10103), .A1(n10038), .B0(n10037), .Y(n6836) );
  NOR2X2 U12548 ( .A(n8967), .B(n8966), .Y(n7740) );
  NOR2X1 U12549 ( .A(n8827), .B(n8826), .Y(n8966) );
  INVX2 U12550 ( .A(n23049), .Y(n22999) );
  INVX1 U12551 ( .A(n22929), .Y(n6838) );
  NAND2X1 U12552 ( .A(n6841), .B(n23051), .Y(n6839) );
  NAND2X1 U12553 ( .A(n6840), .B(n22911), .Y(n23051) );
  OR2X2 U12554 ( .A(n22912), .B(n23083), .Y(n6840) );
  NOR2X1 U12555 ( .A(n23053), .B(n22929), .Y(n6841) );
  OAI21XL U12556 ( .A0(n22327), .A1(n22323), .B0(n22322), .Y(n6842) );
  NOR2X1 U12557 ( .A(n6843), .B(n22321), .Y(n22327) );
  OAI2BB1XL U12558 ( .A0N(n5902), .A1N(n12476), .B0(n12474), .Y(n12470) );
  XOR2X1 U12559 ( .A(n12476), .B(n12471), .Y(n22886) );
  XNOR2X4 U12560 ( .A(n12004), .B(n12005), .Y(n29097) );
  NAND2X2 U12561 ( .A(n10003), .B(n10004), .Y(n12004) );
  INVXL U12562 ( .A(U0_U1_y2[13]), .Y(n12446) );
  NOR2X1 U12563 ( .A(n12502), .B(n12497), .Y(n12451) );
  NAND2X1 U12564 ( .A(n12433), .B(n12448), .Y(n12497) );
  NAND2BX1 U12565 ( .AN(U0_U1_y0[13]), .B(U0_U1_y2[13]), .Y(n12448) );
  NOR2X1 U12566 ( .A(n12449), .B(U0_U1_y2[13]), .Y(n12502) );
  INVXL U12567 ( .A(n13192), .Y(n22296) );
  NAND2XL U12568 ( .A(n22972), .B(n25286), .Y(n13192) );
  AOI21X2 U12569 ( .A0(n9026), .A1(n9101), .B0(n6845), .Y(n9027) );
  OAI21X1 U12570 ( .A0(n9115), .A1(n9112), .B0(n9116), .Y(n6845) );
  NAND2X1 U12571 ( .A(n9025), .B(n9024), .Y(n9116) );
  NAND2X1 U12572 ( .A(n9022), .B(n9023), .Y(n9112) );
  OAI21X2 U12573 ( .A0(n9124), .A1(n9132), .B0(n9125), .Y(n9101) );
  NAND2X1 U12574 ( .A(n9019), .B(n9018), .Y(n9132) );
  NAND2X1 U12575 ( .A(n22983), .B(n22986), .Y(n22978) );
  NAND2BX1 U12576 ( .AN(n24684), .B(n22959), .Y(n22986) );
  XOR2X2 U12577 ( .A(n9207), .B(n6846), .Y(n24684) );
  OAI21XL U12578 ( .A0(n9153), .A1(n9152), .B0(n9151), .Y(n6847) );
  NAND2X1 U12579 ( .A(n9039), .B(n9038), .Y(n9151) );
  NAND2X1 U12580 ( .A(n9032), .B(n9031), .Y(n9081) );
  NAND2X1 U12581 ( .A(n9029), .B(n9030), .Y(n9088) );
  NOR2X1 U12582 ( .A(n9032), .B(n9031), .Y(n9080) );
  NAND2X4 U12583 ( .A(n6850), .B(n6848), .Y(n9233) );
  NOR2X1 U12584 ( .A(n9220), .B(n6852), .Y(n6851) );
  XOR2X2 U12585 ( .A(n7763), .B(n6853), .Y(n24697) );
  XOR2X1 U12586 ( .A(n22884), .B(n5815), .Y(n6853) );
  XOR2X2 U12587 ( .A(n12354), .B(n12353), .Y(n22884) );
  NOR2X2 U12588 ( .A(n13323), .B(n13321), .Y(n6854) );
  NOR2X4 U12589 ( .A(n8008), .B(W2[16]), .Y(n14991) );
  OR2X2 U12590 ( .A(n24666), .B(n24665), .Y(n24735) );
  XOR2X4 U12591 ( .A(n6855), .B(n9041), .Y(n24666) );
  AOI21X4 U12592 ( .A0(n9074), .A1(n9073), .B0(n9037), .Y(n6855) );
  XOR2X4 U12593 ( .A(n6856), .B(n5762), .Y(U1_U1_z1[15]) );
  NOR2X2 U12594 ( .A(n10768), .B(n10776), .Y(n8254) );
  NAND2X1 U12595 ( .A(n7053), .B(BOPD[14]), .Y(n7388) );
  NOR2X2 U12596 ( .A(n7058), .B(BOPD[41]), .Y(n10768) );
  NAND2BX1 U12597 ( .AN(n9080), .B(n5793), .Y(n9034) );
  OAI21XL U12598 ( .A0(n22848), .A1(n22855), .B0(n22849), .Y(n22839) );
  AOI21X1 U12599 ( .A0(n22771), .A1(n14130), .B0(n14135), .Y(n6857) );
  OAI21X4 U12600 ( .A0(n24699), .A1(n7728), .B0(n24694), .Y(n7763) );
  OR2X2 U12601 ( .A(n5814), .B(n24696), .Y(n6859) );
  AOI21X4 U12602 ( .A0(n10761), .A1(n6861), .B0(n6860), .Y(n6878) );
  OAI21X4 U12603 ( .A0(n8256), .A1(n10789), .B0(n8255), .Y(n6860) );
  NOR2X2 U12604 ( .A(n8256), .B(n10790), .Y(n6861) );
  XOR2X4 U12605 ( .A(n6862), .B(n10138), .Y(U0_U0_z1[9]) );
  AOI21X4 U12606 ( .A0(n10140), .A1(n10116), .B0(n10115), .Y(n6863) );
  NAND2X2 U12607 ( .A(n10141), .B(n10116), .Y(n6864) );
  AOI21X4 U12608 ( .A0(n10153), .A1(n10110), .B0(n10109), .Y(n10139) );
  AOI21X4 U12609 ( .A0(n10664), .A1(n6866), .B0(n6865), .Y(n10644) );
  OAI21X2 U12610 ( .A0(n10665), .A1(n10687), .B0(n10666), .Y(n6865) );
  NAND2X1 U12611 ( .A(n8135), .B(BOPB[29]), .Y(n10666) );
  NOR2X2 U12612 ( .A(n10665), .B(n10686), .Y(n6866) );
  NOR2X2 U12613 ( .A(n7051), .B(BOPB[28]), .Y(n10686) );
  OAI21X4 U12614 ( .A0(n10681), .A1(n10684), .B0(n10682), .Y(n10664) );
  NAND2X2 U12615 ( .A(n8166), .B(BOPB[27]), .Y(n10682) );
  NOR2X2 U12616 ( .A(n8193), .B(BOPB[26]), .Y(n10684) );
  NOR2X2 U12617 ( .A(n8166), .B(BOPB[27]), .Y(n10681) );
  NOR2X4 U12618 ( .A(n8043), .B(W0[23]), .Y(n10114) );
  XOR2X2 U12619 ( .A(n6867), .B(n10653), .Y(U1_U0_z0[6]) );
  NOR2X1 U12620 ( .A(n19580), .B(n19562), .Y(n6868) );
  NAND2X1 U12621 ( .A(n19560), .B(n19589), .Y(n19580) );
  NAND2BX1 U12622 ( .AN(n19248), .B(n14852), .Y(n19560) );
  NOR2BX2 U12623 ( .AN(n7878), .B(n6870), .Y(n6869) );
  NOR2X1 U12624 ( .A(n19597), .B(n19556), .Y(n6870) );
  AOI21X2 U12625 ( .A0(n6873), .A1(n13045), .B0(n6871), .Y(n6872) );
  OAI21XL U12626 ( .A0(n13044), .A1(n13043), .B0(n13042), .Y(n6871) );
  NOR2X2 U12627 ( .A(n13006), .B(n13007), .Y(n13044) );
  OAI21X4 U12628 ( .A0(n13047), .A1(n13046), .B0(n6872), .Y(n13603) );
  NAND2X2 U12629 ( .A(n6873), .B(n13040), .Y(n13046) );
  INVX1 U12630 ( .A(n19561), .Y(n6874) );
  OAI21X2 U12631 ( .A0(n24205), .A1(n24204), .B0(n24203), .Y(n24247) );
  NAND2X1 U12632 ( .A(n19553), .B(n20013), .Y(n19604) );
  XOR2X2 U12633 ( .A(n14800), .B(n6917), .Y(n20013) );
  NAND2X1 U12634 ( .A(n23483), .B(n23484), .Y(n23572) );
  NOR2X2 U12635 ( .A(n14658), .B(n14659), .Y(n14820) );
  NOR2X1 U12636 ( .A(n8071), .B(AOPD[31]), .Y(n11005) );
  AND2X2 U12637 ( .A(U2_U0_y2[21]), .B(U2_U0_y0[21]), .Y(n23524) );
  XOR2X1 U12638 ( .A(U2_U0_y2[21]), .B(U2_U0_y0[21]), .Y(n23482) );
  OAI21X1 U12639 ( .A0(n25373), .A1(n12382), .B0(n12381), .Y(n12383) );
  MXI2X1 U12640 ( .A(U1_pipe12[24]), .B(n19801), .S0(n19405), .Y(n4719) );
  XNOR2X1 U12641 ( .A(n19800), .B(n19799), .Y(n19801) );
  NOR2X1 U12642 ( .A(n24100), .B(n24099), .Y(n24156) );
  NOR2X2 U12643 ( .A(n10600), .B(n9555), .Y(n9557) );
  NAND2X1 U12644 ( .A(n10597), .B(n9557), .Y(n9559) );
  AOI21X1 U12645 ( .A0(n13130), .A1(n21992), .B0(n13129), .Y(n22320) );
  NAND2X1 U12646 ( .A(n13371), .B(n13370), .Y(n13372) );
  OAI21X1 U12647 ( .A0(n10336), .A1(n10291), .B0(n10290), .Y(n10294) );
  AOI21X1 U12648 ( .A0(n18495), .A1(n18494), .B0(n18493), .Y(n18862) );
  MXI2X1 U12649 ( .A(U0_pipe3[18]), .B(n24747), .S0(n25273), .Y(n4357) );
  XOR2X1 U12650 ( .A(n24746), .B(n25020), .Y(n24747) );
  NOR2X1 U12651 ( .A(n12602), .B(n12607), .Y(n12619) );
  AOI21X1 U12652 ( .A0(n7025), .A1(n20314), .B0(n20313), .Y(n20315) );
  OAI21X1 U12653 ( .A0(n10817), .A1(n10790), .B0(n10789), .Y(n10793) );
  XOR2X1 U12654 ( .A(n13300), .B(n13299), .Y(n24414) );
  AND2X2 U12655 ( .A(n11418), .B(BOPA[3]), .Y(n6937) );
  NOR2X2 U12656 ( .A(n8309), .B(BOPA[28]), .Y(n8310) );
  CLKINVX3 U12657 ( .A(n7297), .Y(n11585) );
  XNOR2X1 U12658 ( .A(n16666), .B(n16965), .Y(n16667) );
  OR2X2 U12659 ( .A(n8681), .B(n16654), .Y(n7402) );
  INVX1 U12660 ( .A(n16654), .Y(n16700) );
  XOR2X1 U12661 ( .A(n22301), .B(n22300), .Y(n22302) );
  NOR2X1 U12662 ( .A(n9769), .B(n9789), .Y(n9735) );
  NOR2X1 U12663 ( .A(W3[11]), .B(W3[27]), .Y(n9769) );
  AOI21X1 U12664 ( .A0(n9767), .A1(n9735), .B0(n9734), .Y(n9758) );
  OAI21X1 U12665 ( .A0(n9786), .A1(n9797), .B0(n9787), .Y(n9767) );
  NAND2X2 U12666 ( .A(n8028), .B(W2[17]), .Y(n7195) );
  NOR2X1 U12667 ( .A(n8025), .B(W0[27]), .Y(n10119) );
  MXI2X1 U12668 ( .A(U0_pipe13[24]), .B(n25297), .S0(n25318), .Y(n4668) );
  AOI21X1 U12669 ( .A0(n13455), .A1(n13454), .B0(n13453), .Y(n13456) );
  OAI21X1 U12670 ( .A0(n9742), .A1(n9804), .B0(n9743), .Y(n9755) );
  NOR2X1 U12671 ( .A(n8007), .B(W1[29]), .Y(n10205) );
  OAI21X2 U12672 ( .A0(n10198), .A1(n10233), .B0(n10197), .Y(n7360) );
  NAND2X1 U12673 ( .A(n7950), .B(W1[23]), .Y(n10197) );
  AOI21X1 U12674 ( .A0(n18816), .A1(n18709), .B0(n18708), .Y(n18766) );
  INVX1 U12675 ( .A(n18862), .Y(n18816) );
  INVX4 U12676 ( .A(n10414), .Y(n10477) );
  NAND2X1 U12677 ( .A(n16688), .B(n8574), .Y(n8609) );
  AOI21X1 U12678 ( .A0(n17610), .A1(n7969), .B0(n7968), .Y(n17603) );
  AOI21X4 U12679 ( .A0(n9870), .A1(n9815), .B0(n5923), .Y(n9862) );
  NOR2X2 U12680 ( .A(n9833), .B(n9837), .Y(n7374) );
  MXI2X1 U12681 ( .A(U1_pipe2[20]), .B(n19111), .S0(n5812), .Y(n5032) );
  XOR2X1 U12682 ( .A(n19110), .B(n19109), .Y(n19111) );
  OAI21XL U12683 ( .A0(n19153), .A1(n9684), .B0(n9683), .Y(n9685) );
  NOR2X1 U12684 ( .A(n9302), .B(n9303), .Y(n9353) );
  AOI21X1 U12685 ( .A0(n23084), .A1(n23087), .B0(n22910), .Y(n22911) );
  OAI21X1 U12686 ( .A0(n12539), .A1(n12538), .B0(n12537), .Y(n12540) );
  NAND2X2 U12687 ( .A(n7945), .B(W0[21]), .Y(n10111) );
  AOI21X1 U12688 ( .A0(n18859), .A1(n6935), .B0(n18858), .Y(n18860) );
  AOI21X1 U12689 ( .A0(n25207), .A1(n14392), .B0(n14391), .Y(n25155) );
  XOR2X1 U12690 ( .A(n14379), .B(n14378), .Y(n25216) );
  MXI2X1 U12691 ( .A(n7015), .B(n7340), .S0(n13392), .Y(n7233) );
  ADDHX2 U12692 ( .A(U0_U0_y0[22]), .B(U0_U0_y1[22]), .CO(n13260), .S(n13257)
         );
  AOI21X2 U12693 ( .A0(n13427), .A1(n13383), .B0(n13382), .Y(n13392) );
  NOR2X2 U12694 ( .A(W2[28]), .B(W2[12]), .Y(n9941) );
  OAI21X1 U12695 ( .A0(n9806), .A1(n9803), .B0(n9804), .Y(n9745) );
  NOR2X1 U12696 ( .A(W3[10]), .B(W3[26]), .Y(n9789) );
  MXI2X1 U12697 ( .A(U2_pipe3[14]), .B(n18414), .S0(n18987), .Y(n4227) );
  XOR2X1 U12698 ( .A(n18413), .B(n18412), .Y(n18414) );
  NOR2X1 U12699 ( .A(n17980), .B(n17979), .Y(n18044) );
  OAI21X1 U12700 ( .A0(n18359), .A1(n18358), .B0(n18357), .Y(n18406) );
  INVX1 U12701 ( .A(n18301), .Y(n18359) );
  OAI21X1 U12702 ( .A0(n10193), .A1(n10155), .B0(n10154), .Y(n10158) );
  NAND2X2 U12703 ( .A(n7974), .B(W2[26]), .Y(n10300) );
  OAI21X2 U12704 ( .A0(n7280), .A1(n7266), .B0(n7264), .Y(n7263) );
  NOR2X1 U12705 ( .A(n5814), .B(n21946), .Y(n22592) );
  OAI21X2 U12706 ( .A0(n9944), .A1(n9941), .B0(n9942), .Y(n9884) );
  AOI21X1 U12707 ( .A0(n25572), .A1(n25556), .B0(n25555), .Y(n25563) );
  OAI21X1 U12708 ( .A0(n25595), .A1(n25484), .B0(n25483), .Y(n25485) );
  NAND2X1 U12709 ( .A(n6980), .B(n5775), .Y(n25484) );
  XOR2X2 U12710 ( .A(U1_U0_y1[29]), .B(U1_U0_y0[29]), .Y(n9320) );
  MXI2X1 U12711 ( .A(U1_pipe2[22]), .B(n19097), .S0(n5805), .Y(n5034) );
  XNOR2X1 U12712 ( .A(n19096), .B(n19095), .Y(n19097) );
  NAND2X1 U12713 ( .A(n11302), .B(n8338), .Y(n8340) );
  OAI21X2 U12714 ( .A0(n11389), .A1(n11279), .B0(n11278), .Y(n11283) );
  ADDHX2 U12715 ( .A(U2_U0_y1[29]), .B(U2_U0_y0[29]), .CO(n26645), .S(n26607)
         );
  NAND2X1 U12716 ( .A(n21268), .B(n21267), .Y(n21305) );
  AOI21X4 U12717 ( .A0(n24691), .A1(n24701), .B0(n7257), .Y(n24699) );
  OAI21X2 U12718 ( .A0(n24702), .A1(n24690), .B0(n24689), .Y(n7257) );
  AOI21X2 U12719 ( .A0(n24711), .A1(n24686), .B0(n7966), .Y(n24702) );
  NOR2X1 U12720 ( .A(n9090), .B(n9084), .Y(n9163) );
  NAND2XL U12721 ( .A(n20005), .B(n14945), .Y(n20372) );
  NAND2BX2 U12722 ( .AN(n21187), .B(n7344), .Y(n21528) );
  NOR2X1 U12723 ( .A(n19764), .B(n19847), .Y(n19823) );
  OAI21X2 U12724 ( .A0(n7197), .A1(n10906), .B0(n10905), .Y(n10910) );
  INVX1 U12725 ( .A(n26908), .Y(n21573) );
  NAND2X2 U12726 ( .A(n7766), .B(n7765), .Y(n7764) );
  INVX1 U12727 ( .A(n10159), .Y(n10161) );
  AOI21X1 U12728 ( .A0(n6802), .A1(n22924), .B0(n22923), .Y(n23052) );
  OAI21XL U12729 ( .A0(n23068), .A1(n23074), .B0(n23069), .Y(n22923) );
  AND2X2 U12730 ( .A(n7064), .B(n19738), .Y(n16722) );
  AND2X2 U12731 ( .A(n7065), .B(n19738), .Y(n19892) );
  XOR2X2 U12732 ( .A(n8530), .B(n6925), .Y(n19738) );
  INVX1 U12733 ( .A(n22599), .Y(n22614) );
  OAI21X2 U12734 ( .A0(n10246), .A1(n10219), .B0(n10218), .Y(n10222) );
  NOR2X2 U12735 ( .A(n7952), .B(W1[26]), .Y(n10219) );
  NAND2X1 U12736 ( .A(n9705), .B(n19107), .Y(n9707) );
  AOI21X1 U12737 ( .A0(n9705), .A1(n19106), .B0(n9704), .Y(n9706) );
  OAI21X2 U12738 ( .A0(n10269), .A1(n10312), .B0(n10268), .Y(n7192) );
  NAND2X1 U12739 ( .A(n23032), .B(n23037), .Y(n22946) );
  AOI21X1 U12740 ( .A0(n23032), .A1(n22944), .B0(n22943), .Y(n22945) );
  OAI21X1 U12741 ( .A0(n10285), .A1(n10279), .B0(n10278), .Y(n10280) );
  NAND2X1 U12742 ( .A(n10288), .B(n10277), .Y(n10279) );
  NOR3X2 U12743 ( .A(n9829), .B(n7281), .C(n7266), .Y(n7265) );
  XNOR2X2 U12744 ( .A(U1_U0_y1[25]), .B(n7623), .Y(n9312) );
  AOI21X2 U12745 ( .A0(n10331), .A1(n10281), .B0(n10280), .Y(n10327) );
  XNOR2X2 U12746 ( .A(n10294), .B(n10293), .Y(U1_U2_z1[14]) );
  NOR2X2 U12747 ( .A(W0[13]), .B(W0[29]), .Y(n9820) );
  NAND2X2 U12748 ( .A(W0[9]), .B(W0[25]), .Y(n9811) );
  NAND2X2 U12749 ( .A(n10840), .B(n8250), .Y(n7324) );
  XOR2X1 U12750 ( .A(n10163), .B(n10162), .Y(U0_U0_z1[1]) );
  OAI21X2 U12751 ( .A0(n9439), .A1(n9445), .B0(n9440), .Y(n7695) );
  XNOR2X2 U12752 ( .A(n10158), .B(n10157), .Y(U0_U0_z1[3]) );
  INVX1 U12753 ( .A(n10156), .Y(n10157) );
  NOR2X2 U12754 ( .A(n8014), .B(W0[20]), .Y(n10146) );
  OAI21X4 U12755 ( .A0(n10112), .A1(n10147), .B0(n10111), .Y(n10140) );
  NOR2X4 U12756 ( .A(n7945), .B(W0[21]), .Y(n10112) );
  CLKINVX3 U12757 ( .A(n5924), .Y(n6881) );
  CLKINVX3 U12758 ( .A(n5924), .Y(n6882) );
  CLKINVX3 U12759 ( .A(n5924), .Y(n6886) );
  AND2X2 U12760 ( .A(n7390), .B(U2_B_i[15]), .Y(n11437) );
  INVXL U12761 ( .A(U2_B_r[15]), .Y(n7390) );
  NAND2X1 U12762 ( .A(n11438), .B(U2_B_r[14]), .Y(n11539) );
  XOR2X1 U12763 ( .A(n7987), .B(n6897), .Y(n7361) );
  XNOR2X2 U12764 ( .A(n11167), .B(n11166), .Y(U1_U1_z0[9]) );
  NAND2XL U12765 ( .A(n11165), .B(n11164), .Y(n11166) );
  OAI21XL U12766 ( .A0(n11172), .A1(n11168), .B0(n11169), .Y(n11167) );
  INVXL U12767 ( .A(n11163), .Y(n11165) );
  INVXL U12768 ( .A(n11150), .Y(n11152) );
  OAI21X1 U12769 ( .A0(n11141), .A1(n11140), .B0(n11139), .Y(n11145) );
  OAI21X2 U12770 ( .A0(n11141), .A1(n11133), .B0(n11132), .Y(n11138) );
  INVXL U12771 ( .A(n11134), .Y(n11136) );
  OAI21XL U12772 ( .A0(n11172), .A1(n11122), .B0(n11121), .Y(n11127) );
  INVXL U12773 ( .A(n11123), .Y(n11125) );
  NAND2XL U12774 ( .A(n11170), .B(n11169), .Y(n11171) );
  INVXL U12775 ( .A(n11168), .Y(n11170) );
  OAI21XL U12776 ( .A0(n7294), .A1(n11181), .B0(n11182), .Y(n11180) );
  OAI21XL U12777 ( .A0(n10643), .A1(n10610), .B0(n10609), .Y(n10615) );
  INVXL U12778 ( .A(n10611), .Y(n10613) );
  INVXL U12779 ( .A(n11337), .Y(n11338) );
  NAND2XL U12780 ( .A(n12435), .B(n12442), .Y(n12444) );
  INVXL U12781 ( .A(n14710), .Y(n7794) );
  INVXL U12782 ( .A(n10502), .Y(n10504) );
  NAND2XL U12783 ( .A(n10509), .B(n10508), .Y(n10510) );
  INVXL U12784 ( .A(n10507), .Y(n10509) );
  NOR2X2 U12785 ( .A(n11442), .B(n7780), .Y(n7779) );
  NOR2X1 U12786 ( .A(n11530), .B(n11443), .Y(n7780) );
  XOR2X2 U12787 ( .A(n11595), .B(n11594), .Y(U2_U0_z0[3]) );
  NAND2XL U12788 ( .A(n11593), .B(n11592), .Y(n11594) );
  NAND2X1 U12789 ( .A(n7760), .B(n11583), .Y(n11590) );
  XNOR2XL U12790 ( .A(n10839), .B(n10838), .Y(U1_U2_z0[4]) );
  OAI21XL U12791 ( .A0(n8289), .A1(n11104), .B0(n11105), .Y(n11103) );
  NAND2XL U12792 ( .A(n11199), .B(n11198), .Y(n11200) );
  INVXL U12793 ( .A(n11197), .Y(n11199) );
  NAND2X1 U12794 ( .A(n7935), .B(n10623), .Y(n7936) );
  INVXL U12795 ( .A(n10624), .Y(n10626) );
  XOR2X1 U12796 ( .A(n7941), .B(n10620), .Y(U1_U0_z0[12]) );
  NAND2XL U12797 ( .A(n10619), .B(n10618), .Y(n10620) );
  AOI21XL U12798 ( .A0(n7934), .A1(n10606), .B0(n10608), .Y(n7941) );
  NAND2XL U12799 ( .A(n10662), .B(n10661), .Y(n10663) );
  INVXL U12800 ( .A(n10686), .Y(n10688) );
  INVXL U12801 ( .A(n10960), .Y(n10962) );
  INVXL U12802 ( .A(n10980), .Y(n10981) );
  INVXL U12803 ( .A(n10989), .Y(n10991) );
  OAI21X2 U12804 ( .A0(n7197), .A1(n10914), .B0(n10913), .Y(n10919) );
  INVXL U12805 ( .A(n10915), .Y(n10917) );
  INVXL U12806 ( .A(n10868), .Y(n8332) );
  XNOR2X1 U12807 ( .A(n11372), .B(n11371), .Y(U0_U1_z0[4]) );
  NAND2XL U12808 ( .A(n11393), .B(n11392), .Y(n11394) );
  OAI21X1 U12809 ( .A0(n14410), .A1(n14417), .B0(n14411), .Y(n14395) );
  AOI21XL U12810 ( .A0(n13241), .A1(n13333), .B0(n13240), .Y(n13242) );
  NAND2XL U12811 ( .A(n8797), .B(n8876), .Y(n8799) );
  CMPR22X1 U12812 ( .A(U1_U2_y2[28]), .B(U1_U2_y0[28]), .CO(n13901), .S(n13898) );
  NOR2X2 U12813 ( .A(n14696), .B(n14692), .Y(n14703) );
  NOR2X1 U12814 ( .A(n13076), .B(n7882), .Y(n13564) );
  XOR2XL U12815 ( .A(n10528), .B(n10527), .Y(U0_U0_z0[1]) );
  INVXL U12816 ( .A(n10524), .Y(n10526) );
  XOR2XL U12817 ( .A(n11221), .B(n7293), .Y(U1_U1_z0[1]) );
  XOR2XL U12818 ( .A(n10685), .B(n10684), .Y(U1_U0_z0[1]) );
  NAND2XL U12819 ( .A(n10683), .B(n10682), .Y(n10685) );
  INVXL U12820 ( .A(n10681), .Y(n10683) );
  XOR2XL U12821 ( .A(n11400), .B(n11399), .Y(U0_U1_z0[1]) );
  OAI21X1 U12822 ( .A0(n7978), .A1(n8001), .B0(n7236), .Y(n7234) );
  NAND2XL U12823 ( .A(n9544), .B(n9543), .Y(n9545) );
  INVXL U12824 ( .A(n9542), .Y(n9544) );
  NAND2X1 U12825 ( .A(n13692), .B(n7073), .Y(n9503) );
  INVX1 U12826 ( .A(n13062), .Y(n7523) );
  INVX1 U12827 ( .A(n12906), .Y(n12873) );
  AOI21X1 U12828 ( .A0(n14702), .A1(n14703), .B0(n14701), .Y(n14768) );
  XOR2X2 U12829 ( .A(n14862), .B(n14861), .Y(n20029) );
  INVXL U12830 ( .A(n14858), .Y(n14860) );
  NAND2BX1 U12831 ( .AN(n19243), .B(n20041), .Y(n14855) );
  NAND2X1 U12832 ( .A(n13713), .B(n7074), .Y(n9716) );
  NAND2XL U12833 ( .A(n26050), .B(n26056), .Y(n26058) );
  NOR2XL U12834 ( .A(n26049), .B(n26053), .Y(n26056) );
  NAND2XL U12835 ( .A(n23373), .B(n23379), .Y(n23381) );
  AOI21XL U12836 ( .A0(n23379), .A1(n23378), .B0(n23377), .Y(n23380) );
  NOR2XL U12837 ( .A(n23372), .B(n23376), .Y(n23379) );
  AOI21XL U12838 ( .A0(n17814), .A1(n17813), .B0(n17812), .Y(n18011) );
  NOR2XL U12839 ( .A(n17811), .B(n17808), .Y(n17814) );
  NAND2XL U12840 ( .A(n28894), .B(U1_pipe11[1]), .Y(n17743) );
  NOR2XL U12841 ( .A(n28894), .B(U1_pipe11[1]), .Y(n17745) );
  NOR2XL U12842 ( .A(n9235), .B(n9234), .Y(n12349) );
  OAI21XL U12843 ( .A0(n25741), .A1(n25747), .B0(n25742), .Y(n12168) );
  AOI21XL U12844 ( .A0(n13548), .A1(n13547), .B0(n13546), .Y(n17373) );
  CLKINVX3 U12845 ( .A(n20050), .Y(n20016) );
  INVX1 U12846 ( .A(n14902), .Y(n19970) );
  XOR2X2 U12847 ( .A(n13639), .B(n6967), .Y(n14968) );
  NAND2XL U12848 ( .A(n19878), .B(n12300), .Y(n12307) );
  INVXL U12849 ( .A(n20179), .Y(n19377) );
  NAND2XL U12850 ( .A(n24251), .B(n24250), .Y(n24286) );
  NOR2X1 U12851 ( .A(n8066), .B(AOPB[33]), .Y(n10481) );
  NOR2X1 U12852 ( .A(n10490), .B(n10492), .Y(n10480) );
  NAND2X1 U12853 ( .A(n8069), .B(AOPB[32]), .Y(n10486) );
  INVXL U12854 ( .A(n12021), .Y(n12029) );
  NOR2XL U12855 ( .A(U0_U2_y2[7]), .B(U0_U2_y0[7]), .Y(n12021) );
  OR2XL U12856 ( .A(U0_U1_y2[3]), .B(U0_U1_y0[3]), .Y(n12414) );
  OR2XL U12857 ( .A(U0_U1_y1[3]), .B(U0_U1_y0[3]), .Y(n8759) );
  NOR2XL U12858 ( .A(U1_U2_y2[3]), .B(U1_U2_y0[3]), .Y(n13736) );
  NOR2XL U12859 ( .A(U1_U2_y2[7]), .B(U1_U2_y0[7]), .Y(n13745) );
  INVXL U12860 ( .A(n14588), .Y(n14592) );
  NOR2XL U12861 ( .A(U1_U1_y1[3]), .B(U1_U1_y0[3]), .Y(n14588) );
  XNOR2X2 U12862 ( .A(n10468), .B(n10467), .Y(U0_U0_z0[10]) );
  INVXL U12863 ( .A(n10462), .Y(n10463) );
  INVXL U12864 ( .A(n10441), .Y(n10443) );
  INVXL U12865 ( .A(n10409), .Y(n10411) );
  OAI21XL U12866 ( .A0(n10477), .A1(n10420), .B0(n10419), .Y(n10425) );
  NAND2XL U12867 ( .A(n10432), .B(n10431), .Y(n10433) );
  INVX1 U12868 ( .A(n11544), .Y(n7185) );
  INVXL U12869 ( .A(n10755), .Y(n9239) );
  INVXL U12870 ( .A(n10592), .Y(n10594) );
  INVXL U12871 ( .A(n11382), .Y(n11229) );
  INVXL U12872 ( .A(n11316), .Y(n11318) );
  XNOR2X2 U12873 ( .A(n9650), .B(n9649), .Y(U0_U1_z0[9]) );
  NAND2XL U12874 ( .A(n9648), .B(n9647), .Y(n9649) );
  INVXL U12875 ( .A(n9646), .Y(n9648) );
  OAI21X1 U12876 ( .A0(n11348), .A1(n11304), .B0(n11303), .Y(n11309) );
  INVXL U12877 ( .A(n11305), .Y(n11307) );
  INVXL U12878 ( .A(n11288), .Y(n11290) );
  NOR2XL U12879 ( .A(n10017), .B(n10058), .Y(n10043) );
  NAND2XL U12880 ( .A(W3[14]), .B(W3[30]), .Y(n9753) );
  INVX1 U12881 ( .A(n9956), .Y(n7394) );
  NOR2XL U12882 ( .A(n10123), .B(n10172), .Y(n10179) );
  INVX1 U12883 ( .A(n10185), .Y(n7579) );
  NAND2XL U12884 ( .A(n12039), .B(n12046), .Y(n12048) );
  OAI21X1 U12885 ( .A0(n9016), .A1(n9015), .B0(n9014), .Y(n7179) );
  NOR2X1 U12886 ( .A(n13468), .B(n13470), .Y(n7723) );
  NAND2X1 U12887 ( .A(n14672), .B(n14673), .Y(n14795) );
  INVXL U12888 ( .A(n14615), .Y(n14616) );
  NOR2XL U12889 ( .A(U1_U1_y1[10]), .B(U1_U1_y0[10]), .Y(n14615) );
  OAI21X2 U12890 ( .A0(n10522), .A1(n10399), .B0(n10398), .Y(n10403) );
  INVXL U12891 ( .A(n10376), .Y(n10378) );
  OR2X2 U12892 ( .A(n9638), .B(U2_B_r[12]), .Y(n11545) );
  INVXL U12893 ( .A(n10741), .Y(n10743) );
  OAI21X1 U12894 ( .A0(n6878), .A1(n10749), .B0(n10748), .Y(n10753) );
  INVXL U12895 ( .A(n10747), .Y(n10748) );
  XNOR2X2 U12896 ( .A(n10730), .B(n10729), .Y(U1_U2_z0[22]) );
  INVXL U12897 ( .A(n10785), .Y(n10787) );
  OAI21XL U12898 ( .A0(n10829), .A1(n10825), .B0(n10826), .Y(n10824) );
  INVXL U12899 ( .A(n10820), .Y(n10822) );
  NAND2XL U12900 ( .A(n10834), .B(n10833), .Y(n10835) );
  NAND2XL U12901 ( .A(n10863), .B(n10862), .Y(n10864) );
  INVXL U12902 ( .A(n11104), .Y(n11106) );
  OAI21XL U12903 ( .A0(n8289), .A1(n11063), .B0(n11062), .Y(n11068) );
  INVXL U12904 ( .A(n11064), .Y(n11066) );
  OAI21X1 U12905 ( .A0(n6712), .A1(n10573), .B0(n10572), .Y(n10578) );
  INVXL U12906 ( .A(n10574), .Y(n10576) );
  XNOR2X2 U12907 ( .A(n10638), .B(n10637), .Y(U1_U0_z0[9]) );
  NAND2XL U12908 ( .A(n10636), .B(n10635), .Y(n10637) );
  INVXL U12909 ( .A(n10634), .Y(n10636) );
  OAI21XL U12910 ( .A0(n10643), .A1(n10629), .B0(n10628), .Y(n10633) );
  INVXL U12911 ( .A(n10627), .Y(n10629) );
  XOR2X2 U12912 ( .A(n10643), .B(n10642), .Y(U1_U0_z0[8]) );
  NAND2XL U12913 ( .A(n10641), .B(n10640), .Y(n10642) );
  INVXL U12914 ( .A(n10639), .Y(n10641) );
  INVXL U12915 ( .A(n10587), .Y(n10589) );
  OAI21XL U12916 ( .A0(n6712), .A1(n10582), .B0(n10581), .Y(n10586) );
  INVXL U12917 ( .A(n10580), .Y(n10581) );
  OAI21X2 U12918 ( .A0(n6712), .A1(n10549), .B0(n7150), .Y(n7149) );
  INVXL U12919 ( .A(n10550), .Y(n10552) );
  NAND2XL U12920 ( .A(n10932), .B(n10931), .Y(n10933) );
  INVXL U12921 ( .A(n10930), .Y(n10932) );
  INVXL U12922 ( .A(n10926), .Y(n10928) );
  INVXL U12923 ( .A(n10900), .Y(n10902) );
  XNOR2X1 U12924 ( .A(n11013), .B(n11012), .Y(U0_U2_z0[4]) );
  NAND2XL U12925 ( .A(n11017), .B(n11016), .Y(n11018) );
  NAND2XL U12926 ( .A(n11039), .B(n11038), .Y(n11040) );
  INVXL U12927 ( .A(n11037), .Y(n11039) );
  OAI21X1 U12928 ( .A0(n11389), .A1(n11270), .B0(n11269), .Y(n11275) );
  INVXL U12929 ( .A(n11271), .Y(n11273) );
  OAI21X1 U12930 ( .A0(n11389), .A1(n11288), .B0(n11289), .Y(n11287) );
  INVXL U12931 ( .A(n11284), .Y(n11286) );
  INVXL U12932 ( .A(n11277), .Y(n11278) );
  INVXL U12933 ( .A(n11256), .Y(n11258) );
  OAI21X1 U12934 ( .A0(n11389), .A1(n8348), .B0(n8347), .Y(n8351) );
  INVXL U12935 ( .A(n11224), .Y(n8349) );
  NAND2XL U12936 ( .A(n9751), .B(n9740), .Y(n9757) );
  AOI21X1 U12937 ( .A0(n10089), .A1(n10043), .B0(n10042), .Y(n10106) );
  INVXL U12938 ( .A(n10039), .Y(n10040) );
  INVXL U12939 ( .A(n10052), .Y(n10053) );
  OAI21XL U12940 ( .A0(n10123), .A1(n10171), .B0(n10122), .Y(n10182) );
  XOR2X1 U12941 ( .A(n10169), .B(n10170), .Y(U0_U0_z1[6]) );
  INVXL U12942 ( .A(n10168), .Y(n10169) );
  INVXL U12943 ( .A(n10264), .Y(n10265) );
  INVX1 U12944 ( .A(n14330), .Y(n14226) );
  OAI21XL U12945 ( .A0(n12492), .A1(n12453), .B0(n12452), .Y(n12541) );
  AOI21XL U12946 ( .A0(n12451), .A1(n12493), .B0(n12450), .Y(n12452) );
  NAND2XL U12947 ( .A(n12451), .B(n12494), .Y(n12453) );
  NOR2X1 U12948 ( .A(n8972), .B(n8974), .Y(n8936) );
  NOR2XL U12949 ( .A(n8833), .B(n8830), .Y(n8930) );
  CMPR22X1 U12950 ( .A(U0_U1_y1[20]), .B(U0_U1_y0[20]), .CO(n8836), .S(n8812)
         );
  OAI21XL U12951 ( .A0(n8909), .A1(n8931), .B0(n8937), .Y(n8834) );
  CMPR22X1 U12952 ( .A(U1_U2_y2[33]), .B(U1_U2_y0[33]), .CO(n13931), .S(n13928) );
  CMPR22X1 U12953 ( .A(U1_U2_y2[32]), .B(U1_U2_y0[32]), .CO(n13929), .S(n13926) );
  NAND2BX1 U12954 ( .AN(n12936), .B(n7933), .Y(n7822) );
  NAND2X1 U12955 ( .A(n12988), .B(n12989), .Y(n13059) );
  OAI21XL U12956 ( .A0(n12873), .A1(n12901), .B0(n12905), .Y(n12790) );
  CMPR22X1 U12957 ( .A(U1_U2_y1[20]), .B(U1_U2_y0[20]), .CO(n12792), .S(n12766) );
  NOR2X1 U12958 ( .A(n12786), .B(n12789), .Y(n12900) );
  NAND2X1 U12959 ( .A(n13052), .B(n13053), .Y(n13072) );
  NOR2X2 U12960 ( .A(n13053), .B(n13052), .Y(n13074) );
  NAND2BX1 U12961 ( .AN(n13041), .B(n13048), .Y(n7901) );
  XNOR2X2 U12962 ( .A(n10369), .B(n10368), .Y(U0_U0_z0[23]) );
  OAI21X1 U12963 ( .A0(n10522), .A1(n10364), .B0(n10363), .Y(n10369) );
  NAND2XL U12964 ( .A(n11531), .B(n11530), .Y(n11532) );
  XOR2X2 U12965 ( .A(n11555), .B(n11554), .Y(U2_U0_z0[10]) );
  NAND2XL U12966 ( .A(n11553), .B(n11552), .Y(n11554) );
  NAND2XL U12967 ( .A(n10859), .B(n10858), .Y(n10860) );
  INVXL U12968 ( .A(n11055), .Y(n11057) );
  XNOR2X2 U12969 ( .A(n11048), .B(n11047), .Y(U1_U1_z0[25]) );
  OAI21XL U12970 ( .A0(n8289), .A1(n11045), .B0(n11044), .Y(n11048) );
  INVXL U12971 ( .A(n11211), .Y(n11046) );
  XOR2XL U12972 ( .A(n11036), .B(n11035), .Y(U0_U2_z0[1]) );
  NAND2XL U12973 ( .A(n11034), .B(n11033), .Y(n11036) );
  XOR2X1 U12974 ( .A(n9783), .B(n10062), .Y(U2_U0_z2[5]) );
  INVXL U12975 ( .A(n9797), .Y(n9785) );
  INVX1 U12976 ( .A(n11608), .Y(n29101) );
  XOR2X1 U12977 ( .A(n10086), .B(n10085), .Y(U2_U0_z1[2]) );
  INVXL U12978 ( .A(n10084), .Y(n10085) );
  XOR2X1 U12979 ( .A(n10050), .B(n10049), .Y(U2_U0_z1[1]) );
  INVXL U12980 ( .A(n10048), .Y(n10050) );
  NOR2XL U12981 ( .A(n26311), .B(n26315), .Y(n26318) );
  NOR2XL U12982 ( .A(n23848), .B(n23853), .Y(n23856) );
  NOR2XL U12983 ( .A(n23617), .B(n23621), .Y(n23624) );
  NOR2XL U12984 ( .A(n26543), .B(n26548), .Y(n26551) );
  NOR2XL U12985 ( .A(n18424), .B(n18429), .Y(n18432) );
  NOR2XL U12986 ( .A(n20965), .B(n20969), .Y(n20972) );
  NOR2XL U12987 ( .A(n21196), .B(n21201), .Y(n21204) );
  NOR2XL U12988 ( .A(n18259), .B(n18263), .Y(n18266) );
  NOR2XL U12989 ( .A(n18500), .B(n18505), .Y(n18508) );
  NOR2XL U12990 ( .A(n18209), .B(n18213), .Y(n18216) );
  NOR2XL U12991 ( .A(n18443), .B(n18448), .Y(n18451) );
  NOR2XL U12992 ( .A(n20978), .B(n20982), .Y(n20985) );
  NOR2XL U12993 ( .A(n21244), .B(n21249), .Y(n21252) );
  NOR2XL U12994 ( .A(n18196), .B(n18200), .Y(n18203) );
  NOR2XL U12995 ( .A(n18462), .B(n18467), .Y(n18470) );
  NOR2XL U12996 ( .A(n20919), .B(n20923), .Y(n20926) );
  NOR2XL U12997 ( .A(n21147), .B(n21152), .Y(n21155) );
  INVXL U12998 ( .A(n25800), .Y(n20469) );
  CMPR22X1 U12999 ( .A(U2_U0_y1[22]), .B(U2_U0_y0[22]), .CO(n26241), .S(n26189) );
  CMPR22X1 U13000 ( .A(U2_U0_y1[25]), .B(U2_U0_y0[25]), .CO(n26403), .S(n26356) );
  NOR2XL U13001 ( .A(n17752), .B(U2_U0_y0[13]), .Y(n16616) );
  NOR2XL U13002 ( .A(n16601), .B(n16610), .Y(n16613) );
  NOR2XL U13003 ( .A(U2_U0_y0[10]), .B(U2_U0_y2[10]), .Y(n16601) );
  NOR2XL U13004 ( .A(n16586), .B(n16593), .Y(n16596) );
  NOR2XL U13005 ( .A(n20468), .B(U2_U0_y0[13]), .Y(n19057) );
  NOR2XL U13006 ( .A(n19027), .B(n19034), .Y(n19037) );
  OAI21X1 U13007 ( .A0(n24659), .A1(n24753), .B0(n24658), .Y(n24729) );
  AOI21X1 U13008 ( .A0(n24758), .A1(n24657), .B0(n24656), .Y(n24658) );
  NOR2XL U13009 ( .A(n13394), .B(n24519), .Y(n13397) );
  OAI21X1 U13010 ( .A0(n22320), .A1(n7428), .B0(n7427), .Y(n7426) );
  INVXL U13011 ( .A(n25243), .Y(n21751) );
  NAND2XL U13012 ( .A(n12556), .B(n12555), .Y(n12557) );
  INVX1 U13013 ( .A(n12541), .Y(n12515) );
  NOR2XL U13014 ( .A(n13296), .B(n13295), .Y(n13494) );
  NAND2XL U13015 ( .A(n13296), .B(n13295), .Y(n13495) );
  INVXL U13016 ( .A(n13483), .Y(n13294) );
  NOR2X1 U13017 ( .A(n13244), .B(n13245), .Y(n13353) );
  INVXL U13018 ( .A(n12356), .Y(n12283) );
  AND2X2 U13019 ( .A(n14564), .B(n24640), .Y(n7964) );
  NAND2X1 U13020 ( .A(n8811), .B(n8810), .Y(n8832) );
  INVX1 U13021 ( .A(n8834), .Y(n8820) );
  INVXL U13022 ( .A(n14473), .Y(n14475) );
  INVXL U13023 ( .A(n12945), .Y(n7816) );
  NOR2XL U13024 ( .A(n19738), .B(U1_A_r_d0[10]), .Y(n19740) );
  NOR2XL U13025 ( .A(n19738), .B(U1_A_i_d0[10]), .Y(n8659) );
  INVX1 U13026 ( .A(n19976), .Y(n14783) );
  INVXL U13027 ( .A(n8478), .Y(n8481) );
  INVXL U13028 ( .A(n8482), .Y(n8490) );
  INVXL U13029 ( .A(n12936), .Y(n12915) );
  NAND2XL U13030 ( .A(n9355), .B(n9354), .Y(n9356) );
  AOI21XL U13031 ( .A0(n9362), .A1(n7431), .B0(n7714), .Y(n7713) );
  OAI21X1 U13032 ( .A0(n7748), .A1(n7719), .B0(n7717), .Y(n7716) );
  NAND2X1 U13033 ( .A(n13076), .B(n7882), .Y(n13567) );
  OAI21X2 U13034 ( .A0(n29106), .A1(n28751), .B0(n7302), .Y(U2_B_i[0]) );
  AOI21XL U13035 ( .A0(n26678), .A1(n26630), .B0(n26677), .Y(n26734) );
  INVXL U13036 ( .A(n26676), .Y(n26677) );
  NAND2XL U13037 ( .A(n26675), .B(n26630), .Y(n26731) );
  NOR2XL U13038 ( .A(n26682), .B(n26681), .Y(n26733) );
  AOI21XL U13039 ( .A0(n26498), .A1(n26497), .B0(n26496), .Y(n26797) );
  NOR2XL U13040 ( .A(n26486), .B(n26494), .Y(n26497) );
  NAND2XL U13041 ( .A(n26485), .B(n26492), .Y(n26494) );
  AOI21XL U13042 ( .A0(n25867), .A1(n25866), .B0(n25865), .Y(n26059) );
  NOR2XL U13043 ( .A(n25864), .B(n25861), .Y(n25867) );
  NOR2XL U13044 ( .A(n26395), .B(n26394), .Y(n26445) );
  NOR2XL U13045 ( .A(n26321), .B(n26320), .Y(n26442) );
  NOR2XL U13046 ( .A(n26225), .B(n26228), .Y(n26312) );
  NAND2XL U13047 ( .A(n26127), .B(n26133), .Y(n26135) );
  AOI21XL U13048 ( .A0(n26133), .A1(n26132), .B0(n26131), .Y(n26134) );
  NOR2XL U13049 ( .A(n26126), .B(n26130), .Y(n26133) );
  AOI21XL U13050 ( .A0(n23824), .A1(n23823), .B0(n23822), .Y(n24123) );
  NOR2XL U13051 ( .A(n23812), .B(n23820), .Y(n23823) );
  NAND2XL U13052 ( .A(n23811), .B(n23818), .Y(n23820) );
  AOI21XL U13053 ( .A0(n23189), .A1(n23188), .B0(n23187), .Y(n23421) );
  NOR2XL U13054 ( .A(n23186), .B(n23183), .Y(n23189) );
  AOI21XL U13055 ( .A0(n26585), .A1(n26584), .B0(n26583), .Y(n26785) );
  NOR2XL U13056 ( .A(n26573), .B(n26581), .Y(n26584) );
  NAND2XL U13057 ( .A(n26572), .B(n26579), .Y(n26581) );
  AOI21XL U13058 ( .A0(n23843), .A1(n23842), .B0(n23841), .Y(n24136) );
  NOR2XL U13059 ( .A(n23831), .B(n23839), .Y(n23842) );
  NAND2XL U13060 ( .A(n23830), .B(n23837), .Y(n23839) );
  AOI21XL U13061 ( .A0(n23200), .A1(n23199), .B0(n23198), .Y(n23398) );
  NOR2XL U13062 ( .A(n23197), .B(n23194), .Y(n23200) );
  AOI21XL U13063 ( .A0(n23892), .A1(n23891), .B0(n23890), .Y(n24111) );
  NOR2XL U13064 ( .A(n23880), .B(n23888), .Y(n23891) );
  NAND2XL U13065 ( .A(n23879), .B(n23886), .Y(n23888) );
  NOR2XL U13066 ( .A(n26525), .B(n26533), .Y(n26536) );
  NAND2XL U13067 ( .A(n26524), .B(n26531), .Y(n26533) );
  NOR2XL U13068 ( .A(n23465), .B(n23464), .Y(n23491) );
  AOI21XL U13069 ( .A0(n23218), .A1(n23217), .B0(n23216), .Y(n23382) );
  NOR2XL U13070 ( .A(n23215), .B(n23212), .Y(n23218) );
  AOI21XL U13071 ( .A0(n21230), .A1(n21229), .B0(n21228), .Y(n21447) );
  NOR2XL U13072 ( .A(n21218), .B(n21226), .Y(n21229) );
  NAND2XL U13073 ( .A(n21217), .B(n21224), .Y(n21226) );
  NAND2XL U13074 ( .A(n17986), .B(n17992), .Y(n17994) );
  AOI21XL U13075 ( .A0(n17992), .A1(n17991), .B0(n17990), .Y(n17993) );
  NOR2XL U13076 ( .A(n17985), .B(n17989), .Y(n17992) );
  NOR2XL U13077 ( .A(n18100), .B(n18103), .Y(n18232) );
  AOI21XL U13078 ( .A0(n18238), .A1(n18237), .B0(n18236), .Y(n18435) );
  NAND2XL U13079 ( .A(n18232), .B(n18238), .Y(n18426) );
  NOR2XL U13080 ( .A(n18241), .B(n18240), .Y(n18319) );
  NOR2XL U13081 ( .A(n18276), .B(n18275), .Y(n18322) );
  NOR2XL U13082 ( .A(n18319), .B(n18322), .Y(n18425) );
  NAND2XL U13083 ( .A(n20781), .B(n20787), .Y(n20789) );
  AOI21XL U13084 ( .A0(n20787), .A1(n20786), .B0(n20785), .Y(n20788) );
  NOR2XL U13085 ( .A(n20780), .B(n20784), .Y(n20787) );
  NOR2XL U13086 ( .A(n20879), .B(n20882), .Y(n20966) );
  NOR2XL U13087 ( .A(n20975), .B(n20974), .Y(n21076) );
  NOR2XL U13088 ( .A(n21029), .B(n21028), .Y(n21079) );
  NOR2XL U13089 ( .A(n21076), .B(n21079), .Y(n21197) );
  NAND2XL U13090 ( .A(n18071), .B(n18077), .Y(n18079) );
  AOI21XL U13091 ( .A0(n18077), .A1(n18076), .B0(n18075), .Y(n18078) );
  NOR2XL U13092 ( .A(n18070), .B(n18074), .Y(n18077) );
  NOR2XL U13093 ( .A(n18166), .B(n18169), .Y(n18260) );
  NOR2XL U13094 ( .A(n18269), .B(n18268), .Y(n18366) );
  NOR2XL U13095 ( .A(n18314), .B(n18313), .Y(n18369) );
  NOR2XL U13096 ( .A(n18366), .B(n18369), .Y(n18501) );
  NAND2XL U13097 ( .A(n18002), .B(n18008), .Y(n18010) );
  AOI21XL U13098 ( .A0(n18008), .A1(n18007), .B0(n18006), .Y(n18009) );
  NOR2XL U13099 ( .A(n18001), .B(n18005), .Y(n18008) );
  NOR2XL U13100 ( .A(n18110), .B(n18113), .Y(n18210) );
  NOR2XL U13101 ( .A(n18338), .B(n18337), .Y(n18443) );
  NOR2XL U13102 ( .A(n18390), .B(n18389), .Y(n18448) );
  NAND2XL U13103 ( .A(n20759), .B(n20765), .Y(n20767) );
  AOI21XL U13104 ( .A0(n20765), .A1(n20764), .B0(n20763), .Y(n20766) );
  NOR2XL U13105 ( .A(n20758), .B(n20762), .Y(n20765) );
  NOR2XL U13106 ( .A(n20889), .B(n20892), .Y(n20979) );
  NOR2XL U13107 ( .A(n20988), .B(n20987), .Y(n21087) );
  NOR2XL U13108 ( .A(n21038), .B(n21037), .Y(n21090) );
  NOR2XL U13109 ( .A(n21087), .B(n21090), .Y(n21245) );
  NOR2XL U13110 ( .A(n17782), .B(n17781), .Y(n17829) );
  NOR2XL U13111 ( .A(n18059), .B(n18058), .Y(n18129) );
  NAND2XL U13112 ( .A(n18025), .B(n18031), .Y(n18033) );
  AOI21XL U13113 ( .A0(n18031), .A1(n18030), .B0(n18029), .Y(n18032) );
  NOR2XL U13114 ( .A(n18024), .B(n18028), .Y(n18031) );
  NOR2XL U13115 ( .A(n18133), .B(n18132), .Y(n18196) );
  NOR2XL U13116 ( .A(n18126), .B(n18129), .Y(n18197) );
  NOR2XL U13117 ( .A(n20735), .B(n20734), .Y(n20800) );
  NOR2XL U13118 ( .A(n20657), .B(n20660), .Y(n20797) );
  NAND2XL U13119 ( .A(n20711), .B(n20717), .Y(n20719) );
  AOI21XL U13120 ( .A0(n20717), .A1(n20716), .B0(n20715), .Y(n20718) );
  NOR2XL U13121 ( .A(n20710), .B(n20714), .Y(n20717) );
  NOR2XL U13122 ( .A(n20826), .B(n20829), .Y(n20920) );
  NOR2XL U13123 ( .A(n20929), .B(n20928), .Y(n21043) );
  NOR2XL U13124 ( .A(n20995), .B(n20994), .Y(n21046) );
  NOR2XL U13125 ( .A(n21043), .B(n21046), .Y(n21148) );
  NOR2X1 U13126 ( .A(n26146), .B(n26142), .Y(n26149) );
  NOR2X1 U13127 ( .A(n26648), .B(n26647), .Y(n26701) );
  INVXL U13128 ( .A(n23167), .Y(n23170) );
  NOR2X1 U13129 ( .A(n20814), .B(n20815), .Y(n20851) );
  NOR2XL U13130 ( .A(n18591), .B(n18594), .Y(n18701) );
  INVXL U13131 ( .A(n25838), .Y(n25841) );
  INVXL U13132 ( .A(n25009), .Y(n25010) );
  NOR2XL U13133 ( .A(n25050), .B(n9010), .Y(n9012) );
  NAND2X1 U13134 ( .A(n24781), .B(n9004), .Y(n9010) );
  NAND2XL U13135 ( .A(n8914), .B(n8913), .Y(n8915) );
  INVXL U13136 ( .A(n8912), .Y(n8914) );
  NAND2X1 U13137 ( .A(n22200), .B(n22162), .Y(n22164) );
  NAND2XL U13138 ( .A(n7565), .B(n24615), .Y(n24797) );
  NAND2XL U13139 ( .A(n22452), .B(U2_A_r_d[23]), .Y(n24435) );
  AOI21XL U13140 ( .A0(n24501), .A1(n24451), .B0(n24450), .Y(n24465) );
  AND2X1 U13141 ( .A(n14056), .B(n7067), .Y(n24559) );
  AOI21XL U13142 ( .A0(n25503), .A1(n25502), .B0(n25501), .Y(n25554) );
  INVXL U13143 ( .A(n13187), .Y(n13184) );
  NAND2XL U13144 ( .A(n14518), .B(n22897), .Y(n14519) );
  NOR2XL U13145 ( .A(n14518), .B(n22897), .Y(n14520) );
  NAND2XL U13146 ( .A(n25140), .B(U2_A_i_d[23]), .Y(n22170) );
  NAND2XL U13147 ( .A(n21739), .B(U2_A_i_d[2]), .Y(n21740) );
  NAND2XL U13148 ( .A(n21739), .B(U2_A_r_d[2]), .Y(n14336) );
  INVXL U13149 ( .A(n12349), .Y(n9236) );
  NAND2XL U13150 ( .A(n9206), .B(n9219), .Y(n9207) );
  INVXL U13151 ( .A(n9220), .Y(n9206) );
  INVX1 U13152 ( .A(n14025), .Y(n14067) );
  NOR2X1 U13153 ( .A(n25725), .B(n12173), .Y(n12175) );
  NAND2X1 U13154 ( .A(n25728), .B(n25733), .Y(n12173) );
  NOR2X1 U13155 ( .A(n24615), .B(n13114), .Y(n25741) );
  NAND2XL U13156 ( .A(n12116), .B(n12120), .Y(n12117) );
  INVXL U13157 ( .A(n12121), .Y(n12116) );
  INVXL U13158 ( .A(n9080), .Y(n9082) );
  XOR2X2 U13159 ( .A(n12605), .B(n6963), .Y(n22935) );
  INVXL U13160 ( .A(n12602), .Y(n12604) );
  INVXL U13161 ( .A(n12581), .Y(n12569) );
  XOR2X1 U13162 ( .A(n8897), .B(n8854), .Y(n24590) );
  XOR2XL U13163 ( .A(n12515), .B(n12491), .Y(n22892) );
  NAND2XL U13164 ( .A(n12490), .B(n12489), .Y(n12491) );
  INVXL U13165 ( .A(n12488), .Y(n12490) );
  NAND2XL U13166 ( .A(n12504), .B(n12503), .Y(n12505) );
  AOI21XL U13167 ( .A0(n12501), .A1(n12500), .B0(n12499), .Y(n12506) );
  INVXL U13168 ( .A(n12502), .Y(n12504) );
  INVXL U13169 ( .A(n22727), .Y(n22891) );
  NAND2XL U13170 ( .A(n8871), .B(n8870), .Y(n8872) );
  NAND2XL U13171 ( .A(n22452), .B(U2_A_i_d[23]), .Y(n22477) );
  NOR2X1 U13172 ( .A(n22440), .B(n22433), .Y(n22443) );
  INVXL U13173 ( .A(n9225), .Y(n9226) );
  INVXL U13174 ( .A(n9119), .Y(n9121) );
  NAND2XL U13175 ( .A(n8857), .B(n8856), .Y(n8858) );
  INVXL U13176 ( .A(n8855), .Y(n8857) );
  NAND2XL U13177 ( .A(n8886), .B(n8885), .Y(n8887) );
  INVXL U13178 ( .A(n8884), .Y(n8886) );
  OR2X2 U13179 ( .A(n25199), .B(U2_A_r_d[14]), .Y(n25493) );
  OR2X2 U13180 ( .A(n20029), .B(n20028), .Y(n20332) );
  NOR2XL U13181 ( .A(n17374), .B(n13551), .Y(n13553) );
  NAND2XL U13182 ( .A(n7795), .B(n14710), .Y(n14711) );
  INVXL U13183 ( .A(n13808), .Y(n13810) );
  NAND2BX1 U13184 ( .AN(n19996), .B(n14835), .Y(n20308) );
  NAND2BX1 U13185 ( .AN(n20047), .B(n14852), .Y(n20324) );
  NAND2XL U13186 ( .A(n9655), .B(U1_A_i_d0[2]), .Y(n9409) );
  NOR2XL U13187 ( .A(n9655), .B(U1_A_i_d0[2]), .Y(n9410) );
  INVXL U13188 ( .A(n16932), .Y(n17446) );
  INVXL U13189 ( .A(n12813), .Y(n12815) );
  NAND2XL U13190 ( .A(n12912), .B(n12947), .Y(n12913) );
  NAND2XL U13191 ( .A(n17671), .B(n17676), .Y(n12973) );
  NAND2BX1 U13192 ( .AN(n7915), .B(n13069), .Y(n17341) );
  NOR2XL U13193 ( .A(n17621), .B(n14509), .Y(n17609) );
  NAND2XL U13194 ( .A(n19714), .B(U1_A_r_d0[2]), .Y(n19715) );
  NOR2XL U13195 ( .A(n19714), .B(U1_A_r_d0[2]), .Y(n19716) );
  NOR2XL U13196 ( .A(n14951), .B(n19994), .Y(n13912) );
  NOR2X1 U13197 ( .A(n13905), .B(n7464), .Y(n7463) );
  NAND2XL U13198 ( .A(n19714), .B(U1_A_i_d0[2]), .Y(n8645) );
  NOR2XL U13199 ( .A(n19714), .B(U1_A_i_d0[2]), .Y(n8646) );
  AOI21X1 U13200 ( .A0(n16702), .A1(n8667), .B0(n8666), .Y(n16654) );
  INVXL U13201 ( .A(n12865), .Y(n12856) );
  INVXL U13202 ( .A(n14904), .Y(n19961) );
  NAND2X1 U13203 ( .A(n14958), .B(n14949), .Y(n16811) );
  NAND2XL U13204 ( .A(n12332), .B(U1_A_r_d0[24]), .Y(n19798) );
  NAND2XL U13205 ( .A(n9655), .B(U1_A_r_d0[2]), .Y(n9656) );
  NOR2XL U13206 ( .A(n9655), .B(U1_A_r_d0[2]), .Y(n9657) );
  NAND2XL U13207 ( .A(n14745), .B(n19369), .Y(n14746) );
  AOI21XL U13208 ( .A0(n8174), .A1(n8611), .B0(n8610), .Y(n16960) );
  NAND2XL U13209 ( .A(n12838), .B(n12837), .Y(n12839) );
  AOI21XL U13210 ( .A0(n12835), .A1(n12834), .B0(n12833), .Y(n12840) );
  INVXL U13211 ( .A(n12836), .Y(n12838) );
  INVXL U13212 ( .A(n12920), .Y(n12784) );
  INVXL U13213 ( .A(n13863), .Y(n13799) );
  OAI21XL U13214 ( .A0(n19172), .A1(n19462), .B0(n19173), .Y(n13684) );
  OAI21XL U13215 ( .A0(n19411), .A1(n13706), .B0(n13705), .Y(n13707) );
  NAND2X1 U13216 ( .A(n19408), .B(n13708), .Y(n7686) );
  NAND2XL U13217 ( .A(n12853), .B(n12852), .Y(n12854) );
  NAND2XL U13218 ( .A(n14728), .B(n14727), .Y(n14729) );
  AOI21XL U13219 ( .A0(n14725), .A1(n14724), .B0(n14723), .Y(n14730) );
  NAND2XL U13220 ( .A(n14704), .B(n14766), .Y(n14705) );
  NAND2XL U13221 ( .A(n13022), .B(n13021), .Y(n13023) );
  INVXL U13222 ( .A(n13039), .Y(n13013) );
  INVXL U13223 ( .A(n14812), .Y(n14814) );
  NAND2X1 U13224 ( .A(n7915), .B(n20011), .Y(n19550) );
  NOR2XL U13225 ( .A(n28703), .B(n11959), .Y(n11975) );
  NOR2XL U13226 ( .A(n28704), .B(n11641), .Y(n11973) );
  NAND2XL U13227 ( .A(n14897), .B(n29008), .Y(n12337) );
  NAND2BX1 U13228 ( .AN(n9605), .B(n7750), .Y(n7749) );
  NAND2X1 U13229 ( .A(n7313), .B(n7311), .Y(n7319) );
  INVXL U13230 ( .A(n18283), .Y(n18336) );
  AOI21XL U13231 ( .A0(n21590), .A1(n21547), .B0(n21589), .Y(n21648) );
  INVXL U13232 ( .A(n21588), .Y(n21589) );
  NAND2XL U13233 ( .A(n18036), .B(n18035), .Y(n18128) );
  NOR2XL U13234 ( .A(n18036), .B(n18035), .Y(n18126) );
  NAND2XL U13235 ( .A(n18059), .B(n18058), .Y(n18127) );
  INVXL U13236 ( .A(n18476), .Y(n18204) );
  NAND2X1 U13237 ( .A(n26608), .B(n26609), .Y(n26700) );
  OAI21X1 U13238 ( .A0(n26701), .A1(n26700), .B0(n26699), .Y(n26756) );
  NAND2XL U13239 ( .A(n27035), .B(n27034), .Y(n27036) );
  NAND2XL U13240 ( .A(n24163), .B(n24162), .Y(n24200) );
  NAND2XL U13241 ( .A(n24375), .B(n24374), .Y(n24376) );
  INVXL U13242 ( .A(n21693), .Y(n7415) );
  INVXL U13243 ( .A(n18765), .Y(n18806) );
  NAND2X2 U13244 ( .A(n22180), .B(n22177), .Y(n7709) );
  INVXL U13245 ( .A(n24477), .Y(n24480) );
  NAND2BX2 U13246 ( .AN(n9584), .B(n7621), .Y(n17230) );
  OAI21XL U13247 ( .A0(n17233), .A1(n9583), .B0(n9582), .Y(n9584) );
  NOR2XL U13248 ( .A(n17234), .B(n9583), .Y(n9585) );
  NAND2X1 U13249 ( .A(n14959), .B(n19553), .Y(n17334) );
  INVX1 U13250 ( .A(n17304), .Y(n17320) );
  NAND2X1 U13251 ( .A(n20051), .B(n20050), .Y(n20344) );
  NOR2XL U13252 ( .A(n19231), .B(U1_A_i_d0[0]), .Y(n17592) );
  NAND2X1 U13253 ( .A(n9460), .B(n17526), .Y(n7629) );
  NOR2X1 U13254 ( .A(n17528), .B(n9458), .Y(n9460) );
  NOR2XL U13255 ( .A(n17446), .B(n19507), .Y(n17739) );
  NOR2XL U13256 ( .A(n16780), .B(U1_A_r_d0[0]), .Y(n19947) );
  NOR2XL U13257 ( .A(n20180), .B(n16932), .Y(n16929) );
  NAND2X1 U13258 ( .A(n7434), .B(n14951), .Y(n16848) );
  NOR2X1 U13259 ( .A(n12323), .B(n20211), .Y(n12325) );
  OAI21XL U13260 ( .A0(n20195), .A1(n19805), .B0(n19806), .Y(n12330) );
  NOR2XL U13261 ( .A(n19231), .B(U1_A_r_d0[0]), .Y(n19228) );
  NOR2XL U13262 ( .A(n19377), .B(n19507), .Y(n19374) );
  NAND2X1 U13263 ( .A(n19301), .B(n7849), .Y(n7848) );
  NOR2X1 U13264 ( .A(n7846), .B(n7845), .Y(n7844) );
  NOR2XL U13265 ( .A(n19303), .B(n14792), .Y(n7849) );
  OR2X2 U13266 ( .A(n14826), .B(n19542), .Y(n19293) );
  NOR2XL U13267 ( .A(n16996), .B(n8559), .Y(n8561) );
  INVX1 U13268 ( .A(n19408), .Y(n7711) );
  INVX1 U13269 ( .A(n19409), .Y(n7712) );
  NAND2XL U13270 ( .A(n5922), .B(n11946), .Y(n11637) );
  INVX1 U13271 ( .A(n15024), .Y(n11984) );
  NOR2X1 U13272 ( .A(n8128), .B(BOPD[31]), .Y(n10832) );
  NAND2X1 U13273 ( .A(n8117), .B(BOPC[35]), .Y(n11164) );
  INVXL U13274 ( .A(n11192), .Y(n11186) );
  NOR2X2 U13275 ( .A(n8190), .B(BOPB[36]), .Y(n10621) );
  NAND2X1 U13276 ( .A(n8059), .B(AOPC[35]), .Y(n9647) );
  OAI21X2 U13277 ( .A0(n9974), .A1(n9989), .B0(n9975), .Y(n9966) );
  NAND2X2 U13278 ( .A(W1[5]), .B(W1[21]), .Y(n9975) );
  NAND2XL U13279 ( .A(n8101), .B(AOPB[46]), .Y(n10383) );
  INVXL U13280 ( .A(n10469), .Y(n10471) );
  INVXL U13281 ( .A(n10474), .Y(n10476) );
  AOI21X1 U13282 ( .A0(n7185), .A1(n6989), .B0(n11431), .Y(n11432) );
  OAI21X1 U13283 ( .A0(n10832), .A1(n10836), .B0(n10833), .Y(n10818) );
  NAND2X1 U13284 ( .A(n8125), .B(BOPD[32]), .Y(n10826) );
  NOR2X1 U13285 ( .A(n8125), .B(BOPD[32]), .Y(n10825) );
  NAND2X1 U13286 ( .A(n8134), .B(BOPD[30]), .Y(n10836) );
  NOR2BX2 U13287 ( .AN(n10842), .B(n7323), .Y(n7322) );
  NOR2X2 U13288 ( .A(n10841), .B(n10862), .Y(n7323) );
  INVXL U13289 ( .A(n11069), .Y(n11082) );
  INVX1 U13290 ( .A(n10564), .Y(n10556) );
  NAND2XL U13291 ( .A(n8163), .B(BOPB[46]), .Y(n10566) );
  INVXL U13292 ( .A(n11023), .Y(n10873) );
  NAND2XL U13293 ( .A(n8100), .B(AOPD[46]), .Y(n10907) );
  NOR2X1 U13294 ( .A(n8097), .B(AOPD[47]), .Y(n10868) );
  NAND2XL U13295 ( .A(n8099), .B(AOPC[46]), .Y(n11263) );
  INVXL U13296 ( .A(n11297), .Y(n11299) );
  NOR2X1 U13297 ( .A(n8096), .B(AOPC[47]), .Y(n11224) );
  INVXL U13298 ( .A(n11357), .Y(n11359) );
  NAND2XL U13299 ( .A(n11418), .B(BOPA[11]), .Y(n8245) );
  XOR2X1 U13300 ( .A(n8244), .B(n28747), .Y(n7226) );
  NOR2X1 U13301 ( .A(W3[25]), .B(W3[9]), .Y(n9786) );
  OAI21X1 U13302 ( .A0(n8301), .A1(n29106), .B0(n8300), .Y(U2_B_i[1]) );
  NAND2XL U13303 ( .A(n8018), .B(W3[27]), .Y(n10024) );
  INVXL U13304 ( .A(n10179), .Y(n10125) );
  INVXL U13305 ( .A(n10251), .Y(n10206) );
  NOR2X2 U13306 ( .A(n7972), .B(W1[28]), .Y(n10214) );
  INVXL U13307 ( .A(n9952), .Y(n9954) );
  INVX1 U13308 ( .A(n10211), .Y(n7584) );
  AND2XL U13309 ( .A(U0_U0_y2[8]), .B(U0_U0_y0[8]), .Y(n14163) );
  AND2XL U13310 ( .A(U0_U0_y2[10]), .B(U0_U0_y0[10]), .Y(n14166) );
  NAND2XL U13311 ( .A(n14164), .B(n14167), .Y(n14177) );
  NAND2XL U13312 ( .A(n14183), .B(n14186), .Y(n14188) );
  OR2XL U13313 ( .A(U0_U0_y2[2]), .B(U0_U0_y0[2]), .Y(n14183) );
  AOI21XL U13314 ( .A0(n14182), .A1(n14181), .B0(n14180), .Y(n14189) );
  OR2XL U13315 ( .A(U0_U0_y2[1]), .B(U0_U0_y0[1]), .Y(n14182) );
  AND2XL U13316 ( .A(U0_U0_y2[1]), .B(U0_U0_y0[1]), .Y(n14180) );
  AND2XL U13317 ( .A(U0_U0_y2[2]), .B(U0_U0_y0[2]), .Y(n14185) );
  AOI21XL U13318 ( .A0(n14196), .A1(n14195), .B0(n14194), .Y(n14202) );
  AND2XL U13319 ( .A(U0_U0_y2[4]), .B(U0_U0_y0[4]), .Y(n14195) );
  AOI21XL U13320 ( .A0(n14199), .A1(n14198), .B0(n14197), .Y(n14200) );
  AND2XL U13321 ( .A(U0_U0_y2[7]), .B(U0_U0_y0[7]), .Y(n14197) );
  NAND2XL U13322 ( .A(n14192), .B(n14199), .Y(n14201) );
  INVXL U13323 ( .A(n14191), .Y(n14192) );
  NOR2XL U13324 ( .A(U0_U0_y2[6]), .B(U0_U0_y0[6]), .Y(n14191) );
  NAND2XL U13325 ( .A(n14190), .B(n14196), .Y(n14193) );
  AND2XL U13326 ( .A(U0_U2_y1[9]), .B(U0_U2_y0[9]), .Y(n8723) );
  AND2XL U13327 ( .A(U0_U2_y1[8]), .B(U0_U2_y0[8]), .Y(n8724) );
  AND2XL U13328 ( .A(U0_U2_y1[10]), .B(U0_U2_y0[10]), .Y(n8727) );
  NAND2XL U13329 ( .A(n8721), .B(n8728), .Y(n8730) );
  AND2XL U13330 ( .A(U0_U2_y1[1]), .B(U0_U2_y0[1]), .Y(n7995) );
  AND2XL U13331 ( .A(U0_U2_y1[3]), .B(U0_U2_y0[3]), .Y(n7993) );
  AND2XL U13332 ( .A(U0_U2_y1[5]), .B(U0_U2_y0[5]), .Y(n7943) );
  AND2XL U13333 ( .A(U0_U2_y1[7]), .B(U0_U2_y0[7]), .Y(n7944) );
  AND2XL U13334 ( .A(U0_U2_y1[6]), .B(U0_U2_y0[6]), .Y(n8711) );
  INVXL U13335 ( .A(n8702), .Y(n8704) );
  NOR2XL U13336 ( .A(U0_U2_y1[4]), .B(U0_U2_y0[4]), .Y(n8702) );
  NOR2X2 U13337 ( .A(n13264), .B(n13263), .Y(n13384) );
  NAND2XL U13338 ( .A(n13226), .B(n13231), .Y(n13233) );
  INVXL U13339 ( .A(n13224), .Y(n13226) );
  NOR2XL U13340 ( .A(U0_U0_y1[10]), .B(U0_U0_y0[10]), .Y(n13224) );
  AND2XL U13341 ( .A(U0_U0_y1[10]), .B(U0_U0_y0[10]), .Y(n7977) );
  INVXL U13342 ( .A(n13225), .Y(n13231) );
  NOR2XL U13343 ( .A(U0_U0_y1[11]), .B(U0_U0_y0[11]), .Y(n13225) );
  AND2XL U13344 ( .A(U0_U0_y1[11]), .B(U0_U0_y0[11]), .Y(n13230) );
  INVXL U13345 ( .A(n13223), .Y(n13229) );
  NOR2XL U13346 ( .A(U0_U0_y1[9]), .B(U0_U0_y0[9]), .Y(n13223) );
  AND2XL U13347 ( .A(U0_U1_y1[10]), .B(U0_U1_y0[10]), .Y(n8787) );
  AND2XL U13348 ( .A(U0_U1_y1[11]), .B(U0_U1_y0[11]), .Y(n8786) );
  AND2XL U13349 ( .A(U0_U1_y1[9]), .B(U0_U1_y0[9]), .Y(n8783) );
  INVXL U13350 ( .A(n8779), .Y(n8785) );
  NOR2XL U13351 ( .A(U0_U1_y1[9]), .B(U0_U1_y0[9]), .Y(n8779) );
  NAND2XL U13352 ( .A(n8781), .B(n5779), .Y(n8789) );
  AND2XL U13353 ( .A(U0_U1_y1[5]), .B(U0_U1_y0[5]), .Y(n8766) );
  AND2XL U13354 ( .A(U0_U1_y1[4]), .B(U0_U1_y0[4]), .Y(n8767) );
  AND2XL U13355 ( .A(U0_U1_y1[6]), .B(U0_U1_y0[6]), .Y(n8770) );
  AND2XL U13356 ( .A(U0_U1_y1[3]), .B(U0_U1_y0[3]), .Y(n8757) );
  AND2XL U13357 ( .A(U0_U1_y1[1]), .B(U0_U1_y0[1]), .Y(n8753) );
  OR2XL U13358 ( .A(U0_U1_y1[2]), .B(U0_U1_y0[2]), .Y(n8756) );
  NAND2XL U13359 ( .A(n8763), .B(n8768), .Y(n8765) );
  OR2XL U13360 ( .A(U0_U1_y1[4]), .B(U0_U1_y0[4]), .Y(n8763) );
  NAND2XL U13361 ( .A(n8764), .B(n8771), .Y(n8773) );
  CLKINVX3 U13362 ( .A(n7595), .Y(n7593) );
  INVX1 U13363 ( .A(n14394), .Y(n7594) );
  OAI21XL U13364 ( .A0(n14462), .A1(n14465), .B0(n14466), .Y(n14259) );
  AOI21XL U13365 ( .A0(n9243), .A1(n9242), .B0(n9241), .Y(n9251) );
  AND2XL U13366 ( .A(U1_U0_y1[1]), .B(U1_U0_y0[1]), .Y(n9241) );
  OR2XL U13367 ( .A(U1_U0_y1[1]), .B(U1_U0_y0[1]), .Y(n9243) );
  AND2XL U13368 ( .A(U1_U0_y1[0]), .B(U1_U0_y0[0]), .Y(n9242) );
  AND2XL U13369 ( .A(U1_U0_y1[3]), .B(U1_U0_y0[3]), .Y(n9246) );
  AND2XL U13370 ( .A(U1_U0_y1[2]), .B(U1_U0_y0[2]), .Y(n9247) );
  INVXL U13371 ( .A(n9244), .Y(n9245) );
  NOR2XL U13372 ( .A(U1_U0_y1[2]), .B(U1_U0_y0[2]), .Y(n9244) );
  AOI21XL U13373 ( .A0(n9259), .A1(n9258), .B0(n9257), .Y(n9265) );
  AND2XL U13374 ( .A(U1_U0_y1[4]), .B(U1_U0_y0[4]), .Y(n9258) );
  AOI21XL U13375 ( .A0(n9262), .A1(n9261), .B0(n9260), .Y(n9263) );
  AND2XL U13376 ( .A(U1_U0_y1[7]), .B(U1_U0_y0[7]), .Y(n9260) );
  NAND2XL U13377 ( .A(n9255), .B(n9262), .Y(n9264) );
  INVXL U13378 ( .A(n9254), .Y(n9255) );
  NOR2XL U13379 ( .A(U1_U0_y1[6]), .B(U1_U0_y0[6]), .Y(n9254) );
  NAND2XL U13380 ( .A(n9253), .B(n9259), .Y(n9256) );
  INVXL U13381 ( .A(n9252), .Y(n9253) );
  NOR2XL U13382 ( .A(U1_U0_y1[4]), .B(U1_U0_y0[4]), .Y(n9252) );
  AND2XL U13383 ( .A(U1_U0_y1[10]), .B(U1_U0_y0[10]), .Y(n9280) );
  AND2XL U13384 ( .A(U1_U0_y1[11]), .B(U1_U0_y0[11]), .Y(n9279) );
  INVXL U13385 ( .A(n9273), .Y(n9281) );
  NOR2XL U13386 ( .A(U1_U0_y1[11]), .B(U1_U0_y0[11]), .Y(n9273) );
  AND2XL U13387 ( .A(U1_U0_y1[9]), .B(U1_U0_y0[9]), .Y(n9276) );
  NAND2XL U13388 ( .A(n9274), .B(n9281), .Y(n9283) );
  INVXL U13389 ( .A(n9272), .Y(n9274) );
  NOR2XL U13390 ( .A(U1_U0_y1[10]), .B(U1_U0_y0[10]), .Y(n9272) );
  AND2XL U13391 ( .A(U1_U0_y2[1]), .B(U1_U0_y0[1]), .Y(n8360) );
  OR2XL U13392 ( .A(U1_U0_y2[1]), .B(U1_U0_y0[1]), .Y(n8362) );
  AND2XL U13393 ( .A(U1_U0_y2[3]), .B(U1_U0_y0[3]), .Y(n8364) );
  AND2XL U13394 ( .A(U1_U0_y2[2]), .B(U1_U0_y0[2]), .Y(n8365) );
  OR2XL U13395 ( .A(U1_U0_y2[2]), .B(U1_U0_y0[2]), .Y(n8363) );
  AND2XL U13396 ( .A(U1_U0_y2[7]), .B(U1_U0_y0[7]), .Y(n8376) );
  AND2XL U13397 ( .A(U1_U0_y2[6]), .B(U1_U0_y0[6]), .Y(n8377) );
  AOI21XL U13398 ( .A0(n8375), .A1(n8140), .B0(n8374), .Y(n8381) );
  AND2XL U13399 ( .A(U1_U0_y2[4]), .B(U1_U0_y0[4]), .Y(n8140) );
  NAND2XL U13400 ( .A(n8372), .B(n8378), .Y(n8380) );
  NAND2XL U13401 ( .A(n8371), .B(n8375), .Y(n8373) );
  INVXL U13402 ( .A(n8370), .Y(n8371) );
  NOR2XL U13403 ( .A(U1_U0_y2[4]), .B(U1_U0_y0[4]), .Y(n8370) );
  AND2XL U13404 ( .A(U1_U0_y2[10]), .B(U1_U0_y0[10]), .Y(n8393) );
  AND2XL U13405 ( .A(U1_U0_y2[11]), .B(U1_U0_y0[11]), .Y(n8392) );
  AND2XL U13406 ( .A(U1_U0_y2[8]), .B(U1_U0_y0[8]), .Y(n8390) );
  NAND2XL U13407 ( .A(n8387), .B(n8394), .Y(n8396) );
  AND2XL U13408 ( .A(U1_U2_y2[3]), .B(U1_U2_y0[3]), .Y(n13738) );
  AND2XL U13409 ( .A(U1_U2_y2[2]), .B(U1_U2_y0[2]), .Y(n8143) );
  AND2XL U13410 ( .A(U1_U2_y2[5]), .B(U1_U2_y0[5]), .Y(n13748) );
  AND2XL U13411 ( .A(U1_U2_y2[4]), .B(U1_U2_y0[4]), .Y(n13749) );
  AND2XL U13412 ( .A(U1_U2_y2[7]), .B(U1_U2_y0[7]), .Y(n13750) );
  AND2XL U13413 ( .A(U1_U2_y2[6]), .B(U1_U2_y0[6]), .Y(n13751) );
  NAND2XL U13414 ( .A(n13744), .B(n13743), .Y(n13747) );
  OR2XL U13415 ( .A(U1_U2_y2[4]), .B(U1_U2_y0[4]), .Y(n13744) );
  NAND2XL U13416 ( .A(n13763), .B(n13762), .Y(n13769) );
  AND2XL U13417 ( .A(U1_U2_y2[8]), .B(U1_U2_y0[8]), .Y(n13766) );
  AND2XL U13418 ( .A(U1_U2_y2[9]), .B(U1_U2_y0[9]), .Y(n13765) );
  AND2XL U13419 ( .A(U1_U2_y2[10]), .B(U1_U2_y0[10]), .Y(n7957) );
  CMPR22X1 U13420 ( .A(U1_U0_y1[21]), .B(U1_U0_y0[21]), .CO(n9307), .S(n9304)
         );
  NOR2X1 U13421 ( .A(n9497), .B(n9492), .Y(n9482) );
  AOI21X2 U13422 ( .A0(n7330), .A1(n9463), .B0(n7328), .Y(n7327) );
  AOI21XL U13423 ( .A0(n12726), .A1(n12725), .B0(n12724), .Y(n12727) );
  OR2XL U13424 ( .A(U1_U2_y1[6]), .B(U1_U2_y0[6]), .Y(n12719) );
  NAND2XL U13425 ( .A(n12718), .B(n12723), .Y(n12720) );
  OR2XL U13426 ( .A(U1_U2_y1[4]), .B(U1_U2_y0[4]), .Y(n12718) );
  AND2XL U13427 ( .A(U1_U2_y1[8]), .B(U1_U2_y0[8]), .Y(n12738) );
  AND2XL U13428 ( .A(U1_U2_y1[9]), .B(U1_U2_y0[9]), .Y(n12737) );
  AND2XL U13429 ( .A(U1_U2_y1[10]), .B(U1_U2_y0[10]), .Y(n12741) );
  AND2X2 U13430 ( .A(U1_U1_y0[15]), .B(U1_U1_y1[15]), .Y(n14637) );
  AOI21X1 U13431 ( .A0(n12763), .A1(n12808), .B0(n7173), .Y(n12905) );
  NAND2XL U13432 ( .A(AOPB[25]), .B(n8073), .Y(n10514) );
  INVXL U13433 ( .A(U2_B_r[25]), .Y(n11459) );
  NAND2X1 U13434 ( .A(n9638), .B(U2_B_r[12]), .Y(n11544) );
  INVXL U13435 ( .A(n10850), .Y(n10701) );
  NOR2XL U13436 ( .A(n8151), .B(BOPC[50]), .Y(n11207) );
  OAI21XL U13437 ( .A0(n10868), .A1(n10907), .B0(n10867), .Y(n10895) );
  NAND2XL U13438 ( .A(n10896), .B(n10870), .Y(n10872) );
  NAND2XL U13439 ( .A(n11252), .B(n11226), .Y(n11228) );
  INVXL U13440 ( .A(n11383), .Y(n11232) );
  OAI21XL U13441 ( .A0(n11419), .A1(n11418), .B0(n11417), .Y(U2_B_i[20]) );
  NAND2XL U13442 ( .A(n11427), .B(BOPA[20]), .Y(n11417) );
  XOR2X1 U13443 ( .A(n11416), .B(n28708), .Y(n11419) );
  INVXL U13444 ( .A(n9753), .Y(n9754) );
  NOR2XL U13445 ( .A(n9742), .B(n9803), .Y(n9751) );
  OAI21X1 U13446 ( .A0(n28711), .A1(n11430), .B0(n11403), .Y(U2_B_r[18]) );
  NAND2XL U13447 ( .A(BOPA[18]), .B(n11428), .Y(n11403) );
  NAND2XL U13448 ( .A(n8016), .B(W3[29]), .Y(n10030) );
  INVXL U13449 ( .A(n10091), .Y(n10033) );
  OAI21X2 U13450 ( .A0(n7273), .A1(n10172), .B0(n10171), .Y(n10174) );
  AOI21X2 U13451 ( .A0(n10331), .A1(n10287), .B0(n10286), .Y(n10336) );
  INVXL U13452 ( .A(n10284), .Y(n10287) );
  INVXL U13453 ( .A(n10285), .Y(n10286) );
  NOR2XL U13454 ( .A(n12040), .B(n12048), .Y(n12104) );
  NAND2XL U13455 ( .A(n12038), .B(n12043), .Y(n12040) );
  AOI21XL U13456 ( .A0(n12043), .A1(n12042), .B0(n12041), .Y(n12049) );
  AOI21XL U13457 ( .A0(n12046), .A1(n12045), .B0(n12044), .Y(n12047) );
  AND2XL U13458 ( .A(U0_U2_y2[8]), .B(U0_U2_y0[8]), .Y(n12042) );
  AOI21XL U13459 ( .A0(n12035), .A1(n12034), .B0(n12033), .Y(n12102) );
  NOR2XL U13460 ( .A(n12023), .B(n12031), .Y(n12034) );
  CMPR22X1 U13461 ( .A(U0_U1_y2[19]), .B(U0_U1_y0[19]), .CO(n12467), .S(n12464) );
  NOR2XL U13462 ( .A(n12436), .B(n12444), .Y(n12494) );
  NAND2XL U13463 ( .A(n12434), .B(n12439), .Y(n12436) );
  AOI21XL U13464 ( .A0(n12442), .A1(n12441), .B0(n12440), .Y(n12443) );
  AOI21XL U13465 ( .A0(n12439), .A1(n12438), .B0(n12437), .Y(n12445) );
  AND2XL U13466 ( .A(U0_U1_y2[11]), .B(U0_U1_y0[11]), .Y(n12440) );
  NOR2XL U13467 ( .A(n12420), .B(n12428), .Y(n12431) );
  CMPR22X1 U13468 ( .A(U0_U2_y1[14]), .B(U0_U2_y0[14]), .CO(n8739), .S(n8735)
         );
  AOI2BB1X2 U13469 ( .A0N(n13467), .A1N(n13470), .B0(n7722), .Y(n7169) );
  OAI21X2 U13470 ( .A0(n7724), .A1(n13429), .B0(n7723), .Y(n7168) );
  INVXL U13471 ( .A(n13471), .Y(n7722) );
  INVXL U13472 ( .A(n13384), .Y(n13386) );
  NAND2X1 U13473 ( .A(U0_U0_y1[19]), .B(U0_U0_y0[19]), .Y(n7604) );
  NOR2X1 U13474 ( .A(n13354), .B(n13353), .Y(n13317) );
  INVXL U13475 ( .A(n14470), .Y(n14263) );
  INVXL U13476 ( .A(n25162), .Y(n21784) );
  NAND2XL U13477 ( .A(n25162), .B(n8077), .Y(n14455) );
  INVXL U13478 ( .A(n13567), .Y(n13086) );
  NAND2BX1 U13479 ( .AN(n13074), .B(n13071), .Y(n7880) );
  NOR2X1 U13480 ( .A(n13569), .B(n13086), .Y(n7911) );
  NOR2BX1 U13481 ( .AN(U1_U2_y1[33]), .B(n7905), .Y(n13089) );
  NOR2XL U13482 ( .A(n13976), .B(n13963), .Y(n7474) );
  CMPR22X1 U13483 ( .A(U1_U0_y2[20]), .B(U1_U0_y0[20]), .CO(n8418), .S(n8415)
         );
  CMPR22X1 U13484 ( .A(U1_U1_y2[25]), .B(U1_U1_y0[25]), .CO(n12943), .S(n12940) );
  OAI21X1 U13485 ( .A0(n12939), .A1(n12938), .B0(n12937), .Y(n12980) );
  INVX1 U13486 ( .A(n7822), .Y(n12975) );
  CMPR22X1 U13487 ( .A(U1_U1_y2[31]), .B(U1_U1_y0[31]), .CO(n13067), .S(n13064) );
  CMPR22X1 U13488 ( .A(U1_U1_y2[33]), .B(U1_U1_y0[33]), .CO(n13093), .S(n13083) );
  NAND2X1 U13489 ( .A(n13927), .B(n13926), .Y(n13935) );
  INVXL U13490 ( .A(n14763), .Y(n14759) );
  NAND2X1 U13491 ( .A(n14652), .B(n14653), .Y(n14761) );
  AOI21X1 U13492 ( .A0(n14793), .A1(n14674), .B0(n7806), .Y(n14839) );
  CMPR22X1 U13493 ( .A(U1_U0_y2[17]), .B(U1_U0_y0[17]), .CO(n8412), .S(n8409)
         );
  INVXL U13494 ( .A(n8489), .Y(n8483) );
  INVXL U13495 ( .A(n8531), .Y(n8526) );
  NOR2X2 U13496 ( .A(n8417), .B(n8418), .Y(n8534) );
  NAND2X1 U13497 ( .A(n8444), .B(n8445), .Y(n8590) );
  AOI21XL U13498 ( .A0(n12678), .A1(n12677), .B0(n12676), .Y(n12826) );
  NAND2XL U13499 ( .A(n12680), .B(n12681), .Y(n12683) );
  AND2XL U13500 ( .A(U1_U1_y2[11]), .B(U1_U1_y0[11]), .Y(n12685) );
  NAND2X1 U13501 ( .A(n13776), .B(n13775), .Y(n13835) );
  CMPR22X1 U13502 ( .A(U1_U1_y2[19]), .B(U1_U1_y0[19]), .CO(n12705), .S(n12702) );
  NOR2X1 U13503 ( .A(n12780), .B(n12777), .Y(n12890) );
  OAI21X2 U13504 ( .A0(n12780), .A1(n12779), .B0(n12778), .Y(n12893) );
  CMPR22X1 U13505 ( .A(U1_U1_y2[20]), .B(U1_U1_y0[20]), .CO(n12783), .S(n12704) );
  NAND2X1 U13506 ( .A(n12892), .B(n6709), .Y(n12923) );
  NAND2X1 U13507 ( .A(n9306), .B(n9307), .Y(n9434) );
  NOR2X2 U13508 ( .A(n7636), .B(n9486), .Y(n9332) );
  NAND2X1 U13509 ( .A(n9332), .B(n9482), .Y(n9519) );
  XOR2X1 U13510 ( .A(U1_U1_y0[15]), .B(U1_U1_y1[15]), .Y(n14634) );
  NOR2XL U13511 ( .A(n14600), .B(n14608), .Y(n14611) );
  NOR2XL U13512 ( .A(n14617), .B(n14625), .Y(n14718) );
  NAND2XL U13513 ( .A(n14614), .B(n14620), .Y(n14617) );
  AND2XL U13514 ( .A(U1_U1_y1[8]), .B(U1_U1_y0[8]), .Y(n14619) );
  CMPR22X1 U13515 ( .A(U1_U1_y1[18]), .B(U1_U1_y0[18]), .CO(n14643), .S(n14640) );
  NAND2X1 U13516 ( .A(n7451), .B(n14690), .Y(n7450) );
  NAND2XL U13517 ( .A(n7310), .B(n7309), .Y(n7798) );
  CMPR22X1 U13518 ( .A(U1_U1_y1[20]), .B(U1_U1_y0[20]), .CO(n14647), .S(n14644) );
  CMPR22X1 U13519 ( .A(U1_U2_y1[21]), .B(U1_U2_y0[21]), .CO(n12903), .S(n12791) );
  OAI21X1 U13520 ( .A0(n12873), .A1(n12901), .B0(n12905), .Y(n7202) );
  NAND2X1 U13521 ( .A(n12903), .B(n12902), .Y(n12931) );
  NAND2X1 U13522 ( .A(n7894), .B(n7220), .Y(n7439) );
  NOR2X1 U13523 ( .A(n9294), .B(n9295), .Y(n9370) );
  NOR2X2 U13524 ( .A(n9296), .B(n9297), .Y(n9372) );
  INVXL U13525 ( .A(n9376), .Y(n9371) );
  NAND2X1 U13526 ( .A(n6989), .B(n9642), .Y(n9643) );
  INVXL U13527 ( .A(n11431), .Y(n9642) );
  NAND2XL U13528 ( .A(BOPA[17]), .B(n11428), .Y(n11407) );
  INVXL U13529 ( .A(n10104), .Y(n10105) );
  NOR2BX2 U13530 ( .AN(n10183), .B(n7363), .Y(n7362) );
  NAND2BX1 U13531 ( .AN(n9694), .B(n7069), .Y(n9507) );
  NOR2X1 U13532 ( .A(n9340), .B(n9339), .Y(n9528) );
  NAND2XL U13533 ( .A(n9343), .B(n9342), .Y(n9533) );
  NAND2BXL U13534 ( .AN(n9529), .B(n9341), .Y(n7664) );
  NOR2XL U13535 ( .A(n26484), .B(n26489), .Y(n26492) );
  NOR2XL U13536 ( .A(n26256), .B(n26260), .Y(n26263) );
  NOR2XL U13537 ( .A(n23810), .B(n23815), .Y(n23818) );
  NOR2XL U13538 ( .A(n26571), .B(n26576), .Y(n26579) );
  NOR2XL U13539 ( .A(n26333), .B(n26337), .Y(n26340) );
  NOR2XL U13540 ( .A(n23829), .B(n23834), .Y(n23837) );
  NOR2XL U13541 ( .A(n23878), .B(n23883), .Y(n23886) );
  NOR2XL U13542 ( .A(n23641), .B(n23645), .Y(n23648) );
  NOR2XL U13543 ( .A(n26523), .B(n26528), .Y(n26531) );
  NOR2XL U13544 ( .A(n26298), .B(n26302), .Y(n26305) );
  NOR2XL U13545 ( .A(n21216), .B(n21221), .Y(n21224) );
  AOI21XL U13546 ( .A0(n18470), .A1(n18469), .B0(n18468), .Y(n18471) );
  NOR2XL U13547 ( .A(n21000), .B(n21004), .Y(n21007) );
  NOR2XL U13548 ( .A(U2_U0_y0[11]), .B(U2_U0_y2[11]), .Y(n16610) );
  NOR2XL U13549 ( .A(U2_U0_y0[9]), .B(U2_U0_y2[9]), .Y(n16607) );
  NOR2XL U13550 ( .A(U2_U0_y0[7]), .B(U2_U0_y2[7]), .Y(n16593) );
  NOR2XL U13551 ( .A(U2_U0_y0[7]), .B(U2_U0_y1[7]), .Y(n19034) );
  AND2XL U13552 ( .A(n24539), .B(n24541), .Y(n6981) );
  NOR2XL U13553 ( .A(n14572), .B(n22958), .Y(n14574) );
  AND2XL U13554 ( .A(n21751), .B(U2_A_i_d[7]), .Y(n21752) );
  INVXL U13555 ( .A(n14359), .Y(n14290) );
  XNOR2X1 U13556 ( .A(n14281), .B(n14280), .Y(n25251) );
  NAND2XL U13557 ( .A(n14279), .B(n14278), .Y(n14280) );
  CLKINVX3 U13558 ( .A(n14100), .Y(n14048) );
  NOR2XL U13559 ( .A(n22535), .B(n22533), .Y(n14034) );
  NAND2XL U13560 ( .A(n14412), .B(n14411), .Y(n14413) );
  OAI21XL U13561 ( .A0(n14420), .A1(n14416), .B0(n14417), .Y(n14414) );
  NOR2XL U13562 ( .A(n9450), .B(U1_A_i_d0[10]), .Y(n9452) );
  NOR2X2 U13563 ( .A(n13088), .B(n13089), .Y(n13568) );
  NAND2XL U13564 ( .A(n13088), .B(n13089), .Y(n13566) );
  INVXL U13565 ( .A(n12296), .Y(n19727) );
  INVX1 U13566 ( .A(n12290), .Y(n19714) );
  AND2XL U13567 ( .A(n19727), .B(U1_A_i_d0[7]), .Y(n8653) );
  OR2X2 U13568 ( .A(n19745), .B(U1_A_i_d0[12]), .Y(n8663) );
  NAND2XL U13569 ( .A(n8456), .B(n8455), .Y(n8632) );
  INVXL U13570 ( .A(n14911), .Y(n19957) );
  NOR2XL U13571 ( .A(n14937), .B(n16871), .Y(n14939) );
  NAND2X1 U13572 ( .A(n13065), .B(n13064), .Y(n13080) );
  NOR2X1 U13573 ( .A(n13064), .B(n13065), .Y(n13078) );
  NAND2XL U13574 ( .A(n13972), .B(n13971), .Y(n13975) );
  NAND2XL U13575 ( .A(n13985), .B(n13984), .Y(n13989) );
  NAND2X1 U13576 ( .A(n13699), .B(n7071), .Y(n7679) );
  INVXL U13577 ( .A(n8635), .Y(n8637) );
  NAND2X1 U13578 ( .A(n12703), .B(n12702), .Y(n12779) );
  NAND2X1 U13579 ( .A(n12704), .B(n12705), .Y(n12778) );
  NAND2X1 U13580 ( .A(n19134), .B(n19138), .Y(n13697) );
  NAND2X1 U13581 ( .A(n14634), .B(n14635), .Y(n14738) );
  NAND2X1 U13582 ( .A(n14642), .B(n14643), .Y(n14697) );
  AOI21X1 U13583 ( .A0(n7879), .A1(n6947), .B0(n19555), .Y(n7878) );
  NAND2X1 U13584 ( .A(n9294), .B(n9295), .Y(n9376) );
  INVXL U13585 ( .A(n9366), .Y(n9369) );
  INVXL U13586 ( .A(n9370), .Y(n9377) );
  OAI21XL U13587 ( .A0(n20045), .A1(n20018), .B0(n20017), .Y(n20038) );
  NOR2XL U13588 ( .A(n19251), .B(n14854), .Y(n19239) );
  INVXL U13589 ( .A(n24677), .Y(n24688) );
  NOR2X1 U13590 ( .A(n20033), .B(n20032), .Y(n20330) );
  NOR2X1 U13591 ( .A(n13709), .B(n7072), .Y(n7671) );
  NOR2XL U13592 ( .A(n19092), .B(n9714), .Y(n19081) );
  INVXL U13593 ( .A(n13713), .Y(n9537) );
  NOR2X1 U13594 ( .A(n19074), .B(n9719), .Y(n7678) );
  NOR2XL U13595 ( .A(n26380), .B(n26383), .Y(n26485) );
  NOR2XL U13596 ( .A(n26328), .B(n26327), .Y(n26383) );
  NOR2XL U13597 ( .A(n26266), .B(n26265), .Y(n26380) );
  NOR2XL U13598 ( .A(n26166), .B(n26169), .Y(n26257) );
  NOR2XL U13599 ( .A(n26105), .B(n26104), .Y(n26169) );
  NOR2XL U13600 ( .A(n26005), .B(n26004), .Y(n26053) );
  NOR2XL U13601 ( .A(n25957), .B(n25960), .Y(n26050) );
  NOR2XL U13602 ( .A(n25869), .B(n25868), .Y(n25957) );
  NOR2XL U13603 ( .A(n25909), .B(n25908), .Y(n25960) );
  NOR2XL U13604 ( .A(n25816), .B(n25815), .Y(n25864) );
  NOR2XL U13605 ( .A(n26161), .B(n26160), .Y(n26228) );
  NOR2XL U13606 ( .A(n26044), .B(n26043), .Y(n26130) );
  NOR2XL U13607 ( .A(n25993), .B(n25996), .Y(n26127) );
  NOR2XL U13608 ( .A(n25881), .B(n25880), .Y(n25928) );
  AOI21XL U13609 ( .A0(n24003), .A1(n23973), .B0(n24002), .Y(n24083) );
  INVXL U13610 ( .A(n24001), .Y(n24002) );
  NAND2XL U13611 ( .A(n24000), .B(n23973), .Y(n24080) );
  NOR2XL U13612 ( .A(n24007), .B(n24006), .Y(n24082) );
  NOR2XL U13613 ( .A(n23728), .B(n23731), .Y(n23811) );
  AOI21XL U13614 ( .A0(n23589), .A1(n23588), .B0(n23587), .Y(n23821) );
  NAND2XL U13615 ( .A(n23583), .B(n23589), .Y(n23812) );
  NOR2XL U13616 ( .A(n23658), .B(n23657), .Y(n23731) );
  NOR2XL U13617 ( .A(n23592), .B(n23591), .Y(n23728) );
  NOR2XL U13618 ( .A(n23514), .B(n23517), .Y(n23583) );
  NOR2XL U13619 ( .A(n23437), .B(n23436), .Y(n23517) );
  NAND2XL U13620 ( .A(n23412), .B(n23418), .Y(n23420) );
  AOI21XL U13621 ( .A0(n23418), .A1(n23417), .B0(n23416), .Y(n23419) );
  NOR2XL U13622 ( .A(n23411), .B(n23415), .Y(n23418) );
  NOR2XL U13623 ( .A(n23355), .B(n23354), .Y(n23415) );
  NOR2XL U13624 ( .A(n23309), .B(n23312), .Y(n23412) );
  NOR2XL U13625 ( .A(n23235), .B(n23234), .Y(n23312) );
  NOR2XL U13626 ( .A(n23191), .B(n23190), .Y(n23309) );
  NOR2XL U13627 ( .A(n23139), .B(n23138), .Y(n23186) );
  NAND2XL U13628 ( .A(n28890), .B(U0_pipe11[1]), .Y(n23124) );
  NOR2XL U13629 ( .A(n28890), .B(U0_pipe11[1]), .Y(n23126) );
  NAND2XL U13630 ( .A(n26586), .B(n26620), .Y(n26742) );
  AOI21XL U13631 ( .A0(n26620), .A1(n26666), .B0(n26665), .Y(n26745) );
  INVXL U13632 ( .A(n26664), .Y(n26665) );
  NOR2XL U13633 ( .A(n26670), .B(n26669), .Y(n26744) );
  NOR2XL U13634 ( .A(n26422), .B(n26425), .Y(n26572) );
  NOR2XL U13635 ( .A(n26375), .B(n26374), .Y(n26425) );
  NOR2XL U13636 ( .A(n26343), .B(n26342), .Y(n26422) );
  NOR2XL U13637 ( .A(n26196), .B(n26199), .Y(n26334) );
  NOR2XL U13638 ( .A(n26183), .B(n26182), .Y(n26199) );
  NAND2XL U13639 ( .A(n26089), .B(n26095), .Y(n26097) );
  AOI21XL U13640 ( .A0(n26095), .A1(n26094), .B0(n26093), .Y(n26096) );
  NOR2XL U13641 ( .A(n26088), .B(n26092), .Y(n26095) );
  NOR2XL U13642 ( .A(n26074), .B(n26073), .Y(n26092) );
  NOR2XL U13643 ( .A(n26020), .B(n26023), .Y(n26089) );
  NOR2XL U13644 ( .A(n25856), .B(n25855), .Y(n25898) );
  AOI21XL U13645 ( .A0(n24015), .A1(n23963), .B0(n24014), .Y(n24072) );
  INVXL U13646 ( .A(n24013), .Y(n24014) );
  NAND2XL U13647 ( .A(n24012), .B(n23963), .Y(n24069) );
  NOR2XL U13648 ( .A(n24019), .B(n24018), .Y(n24071) );
  NOR2XL U13649 ( .A(n23717), .B(n23720), .Y(n23830) );
  AOI21XL U13650 ( .A0(n23602), .A1(n23601), .B0(n23600), .Y(n23840) );
  NAND2XL U13651 ( .A(n23596), .B(n23602), .Y(n23831) );
  NOR2XL U13652 ( .A(n23667), .B(n23666), .Y(n23720) );
  NOR2XL U13653 ( .A(n23605), .B(n23604), .Y(n23717) );
  NOR2XL U13654 ( .A(n23498), .B(n23501), .Y(n23596) );
  NOR2XL U13655 ( .A(n23443), .B(n23442), .Y(n23501) );
  NAND2XL U13656 ( .A(n23389), .B(n23395), .Y(n23397) );
  AOI21XL U13657 ( .A0(n23395), .A1(n23394), .B0(n23393), .Y(n23396) );
  NOR2XL U13658 ( .A(n23388), .B(n23392), .Y(n23395) );
  NOR2XL U13659 ( .A(n23338), .B(n23337), .Y(n23392) );
  NOR2XL U13660 ( .A(n23291), .B(n23294), .Y(n23389) );
  NOR2XL U13661 ( .A(n23244), .B(n23243), .Y(n23294) );
  NOR2XL U13662 ( .A(n23202), .B(n23201), .Y(n23291) );
  NOR2XL U13663 ( .A(n23146), .B(n23145), .Y(n23197) );
  NAND2XL U13664 ( .A(n28889), .B(U0_pipe5[1]), .Y(n22425) );
  NOR2XL U13665 ( .A(n28889), .B(U0_pipe5[1]), .Y(n22427) );
  NAND2XL U13666 ( .A(n28888), .B(U0_pipe1[1]), .Y(n25115) );
  NOR2XL U13667 ( .A(n28888), .B(U0_pipe1[1]), .Y(n25117) );
  NAND2XL U13668 ( .A(n23893), .B(n23943), .Y(n24047) );
  AOI21XL U13669 ( .A0(n23943), .A1(n23991), .B0(n23990), .Y(n24050) );
  INVXL U13670 ( .A(n23989), .Y(n23990) );
  NOR2XL U13671 ( .A(n23995), .B(n23994), .Y(n24049) );
  NOR2XL U13672 ( .A(n23750), .B(n23753), .Y(n23879) );
  NOR2XL U13673 ( .A(n23701), .B(n23700), .Y(n23753) );
  NOR2XL U13674 ( .A(n23651), .B(n23650), .Y(n23750) );
  NOR2XL U13675 ( .A(n23550), .B(n23553), .Y(n23642) );
  NOR2XL U13676 ( .A(n23509), .B(n23508), .Y(n23553) );
  NAND2XL U13677 ( .A(n23449), .B(n23455), .Y(n23457) );
  AOI21XL U13678 ( .A0(n23455), .A1(n23454), .B0(n23453), .Y(n23456) );
  NOR2XL U13679 ( .A(n23448), .B(n23452), .Y(n23455) );
  NOR2XL U13680 ( .A(n23406), .B(n23405), .Y(n23452) );
  NOR2XL U13681 ( .A(n23343), .B(n23346), .Y(n23449) );
  NOR2XL U13682 ( .A(n23207), .B(n23206), .Y(n23252) );
  NAND2XL U13683 ( .A(n26538), .B(n26613), .Y(n26709) );
  AOI21XL U13684 ( .A0(n26613), .A1(n26655), .B0(n26654), .Y(n26712) );
  INVXL U13685 ( .A(n26653), .Y(n26654) );
  NOR2XL U13686 ( .A(n26659), .B(n26658), .Y(n26711) );
  NOR2XL U13687 ( .A(n26411), .B(n26414), .Y(n26524) );
  NOR2XL U13688 ( .A(n26366), .B(n26365), .Y(n26414) );
  NOR2XL U13689 ( .A(n26308), .B(n26307), .Y(n26411) );
  NOR2XL U13690 ( .A(n26215), .B(n26218), .Y(n26299) );
  NOR2XL U13691 ( .A(n26177), .B(n26176), .Y(n26218) );
  NAND2XL U13692 ( .A(n26111), .B(n26117), .Y(n26119) );
  AOI21XL U13693 ( .A0(n26117), .A1(n26116), .B0(n26115), .Y(n26118) );
  NOR2XL U13694 ( .A(n26110), .B(n26114), .Y(n26117) );
  NOR2XL U13695 ( .A(n26067), .B(n26066), .Y(n26114) );
  NOR2XL U13696 ( .A(n26010), .B(n26013), .Y(n26111) );
  NOR2XL U13697 ( .A(n25874), .B(n25873), .Y(n25917) );
  AOI21XL U13698 ( .A0(n24027), .A1(n23953), .B0(n24026), .Y(n24061) );
  INVXL U13699 ( .A(n24025), .Y(n24026) );
  NAND2XL U13700 ( .A(n24024), .B(n23953), .Y(n24058) );
  NOR2XL U13701 ( .A(n24031), .B(n24030), .Y(n24060) );
  AOI21XL U13702 ( .A0(n23862), .A1(n23861), .B0(n23860), .Y(n24148) );
  NOR2XL U13703 ( .A(n23850), .B(n23858), .Y(n23861) );
  NAND2XL U13704 ( .A(n23849), .B(n23856), .Y(n23858) );
  NOR2XL U13705 ( .A(n23864), .B(n23863), .Y(n23949) );
  NOR2XL U13706 ( .A(n23706), .B(n23709), .Y(n23849) );
  NOR2XL U13707 ( .A(n23676), .B(n23675), .Y(n23709) );
  NOR2XL U13708 ( .A(n23627), .B(n23626), .Y(n23706) );
  NOR2XL U13709 ( .A(n23536), .B(n23535), .Y(n23621) );
  NOR2XL U13710 ( .A(n23495), .B(n23494), .Y(n23617) );
  NOR2XL U13711 ( .A(n23331), .B(n23330), .Y(n23376) );
  NOR2XL U13712 ( .A(n23281), .B(n23284), .Y(n23373) );
  NOR2XL U13713 ( .A(n23263), .B(n23262), .Y(n23284) );
  NOR2XL U13714 ( .A(n23220), .B(n23219), .Y(n23281) );
  NOR2XL U13715 ( .A(n23161), .B(n23160), .Y(n23215) );
  NAND2XL U13716 ( .A(n28891), .B(U0_pipe7[1]), .Y(n22101) );
  NOR2XL U13717 ( .A(n28891), .B(U0_pipe7[1]), .Y(n22103) );
  AOI21XL U13718 ( .A0(n26637), .A1(n26689), .B0(n26688), .Y(n26723) );
  INVXL U13719 ( .A(n26687), .Y(n26688) );
  NAND2XL U13720 ( .A(n26558), .B(n26637), .Y(n26720) );
  NOR2XL U13721 ( .A(n26693), .B(n26692), .Y(n26722) );
  AOI21XL U13722 ( .A0(n26557), .A1(n26556), .B0(n26555), .Y(n26809) );
  NOR2XL U13723 ( .A(n26545), .B(n26553), .Y(n26556) );
  NAND2XL U13724 ( .A(n26544), .B(n26551), .Y(n26553) );
  NOR2XL U13725 ( .A(n26442), .B(n26445), .Y(n26544) );
  NOR2XL U13726 ( .A(n21107), .B(n21110), .Y(n21217) );
  INVXL U13727 ( .A(n21326), .Y(n21327) );
  NAND2XL U13728 ( .A(n21231), .B(n21298), .Y(n21380) );
  NOR2XL U13729 ( .A(n21332), .B(n21331), .Y(n21382) );
  NOR2XL U13730 ( .A(n17760), .B(n17759), .Y(n17800) );
  NAND2XL U13731 ( .A(n28895), .B(U1_pipe7[1]), .Y(n16933) );
  NOR2XL U13732 ( .A(n28895), .B(U1_pipe7[1]), .Y(n16935) );
  NOR2XL U13733 ( .A(n17947), .B(n17946), .Y(n17989) );
  NOR2XL U13734 ( .A(n17923), .B(n17926), .Y(n17986) );
  NOR2XL U13735 ( .A(n18087), .B(n18086), .Y(n18103) );
  AOI21XL U13736 ( .A0(n18616), .A1(n18585), .B0(n18615), .Y(n18692) );
  INVXL U13737 ( .A(n18614), .Y(n18615) );
  NAND2XL U13738 ( .A(n18613), .B(n18585), .Y(n18689) );
  NOR2XL U13739 ( .A(n18620), .B(n18619), .Y(n18691) );
  AOI21XL U13740 ( .A0(n18438), .A1(n18437), .B0(n18436), .Y(n18759) );
  NOR2XL U13741 ( .A(n18426), .B(n18434), .Y(n18437) );
  NAND2XL U13742 ( .A(n18425), .B(n18432), .Y(n18434) );
  NOR2XL U13743 ( .A(n20535), .B(n20534), .Y(n20582) );
  NOR2XL U13744 ( .A(n20728), .B(n20727), .Y(n20784) );
  NOR2XL U13745 ( .A(n20674), .B(n20677), .Y(n20781) );
  NOR2XL U13746 ( .A(n20837), .B(n20836), .Y(n20882) );
  NOR2XL U13747 ( .A(n20886), .B(n20885), .Y(n20965) );
  NOR2XL U13748 ( .A(n20936), .B(n20935), .Y(n20969) );
  AOI21XL U13749 ( .A0(n21274), .A1(n21317), .B0(n21316), .Y(n21372) );
  INVXL U13750 ( .A(n21315), .Y(n21316) );
  NAND2XL U13751 ( .A(n21211), .B(n21274), .Y(n21369) );
  NOR2XL U13752 ( .A(n21321), .B(n21320), .Y(n21371) );
  AOI21XL U13753 ( .A0(n21210), .A1(n21209), .B0(n21208), .Y(n21435) );
  NOR2XL U13754 ( .A(n21198), .B(n21206), .Y(n21209) );
  NAND2XL U13755 ( .A(n21197), .B(n21204), .Y(n21206) );
  NOR2XL U13756 ( .A(n17821), .B(n17820), .Y(n17869) );
  NOR2XL U13757 ( .A(n18019), .B(n18018), .Y(n18074) );
  NOR2XL U13758 ( .A(n17959), .B(n17962), .Y(n18071) );
  NOR2XL U13759 ( .A(n18121), .B(n18120), .Y(n18169) );
  NOR2XL U13760 ( .A(n18173), .B(n18172), .Y(n18259) );
  NOR2XL U13761 ( .A(n18226), .B(n18225), .Y(n18263) );
  AOI21XL U13762 ( .A0(n18555), .A1(n18604), .B0(n18603), .Y(n18659) );
  INVXL U13763 ( .A(n18602), .Y(n18603) );
  NAND2XL U13764 ( .A(n18515), .B(n18555), .Y(n18656) );
  NOR2XL U13765 ( .A(n18608), .B(n18607), .Y(n18658) );
  AOI21XL U13766 ( .A0(n18514), .A1(n18513), .B0(n18512), .Y(n18722) );
  NOR2XL U13767 ( .A(n18502), .B(n18510), .Y(n18513) );
  NAND2XL U13768 ( .A(n18501), .B(n18508), .Y(n18510) );
  NOR2XL U13769 ( .A(n17767), .B(n17766), .Y(n17811) );
  NAND2XL U13770 ( .A(n28893), .B(U1_pipe5[1]), .Y(n17167) );
  NOR2XL U13771 ( .A(n28893), .B(U1_pipe5[1]), .Y(n17169) );
  NOR2XL U13772 ( .A(n17816), .B(n17815), .Y(n17905) );
  NOR2XL U13773 ( .A(n17861), .B(n17860), .Y(n17908) );
  NOR2XL U13774 ( .A(n17954), .B(n17953), .Y(n18005) );
  NOR2XL U13775 ( .A(n17905), .B(n17908), .Y(n18002) );
  NOR2XL U13776 ( .A(n18065), .B(n18064), .Y(n18113) );
  NOR2XL U13777 ( .A(n18117), .B(n18116), .Y(n18209) );
  NOR2XL U13778 ( .A(n18161), .B(n18160), .Y(n18213) );
  AOI21XL U13779 ( .A0(n18628), .A1(n18575), .B0(n18627), .Y(n18681) );
  INVXL U13780 ( .A(n18626), .Y(n18627) );
  NAND2XL U13781 ( .A(n18625), .B(n18575), .Y(n18678) );
  NOR2XL U13782 ( .A(n18632), .B(n18631), .Y(n18680) );
  AOI21XL U13783 ( .A0(n18457), .A1(n18456), .B0(n18455), .Y(n18747) );
  NOR2XL U13784 ( .A(n18445), .B(n18453), .Y(n18456) );
  NAND2XL U13785 ( .A(n18444), .B(n18451), .Y(n18453) );
  NOR2XL U13786 ( .A(n20542), .B(n20541), .Y(n20563) );
  NOR2XL U13787 ( .A(n20705), .B(n20704), .Y(n20762) );
  NOR2XL U13788 ( .A(n20684), .B(n20687), .Y(n20759) );
  NOR2XL U13789 ( .A(n20843), .B(n20842), .Y(n20892) );
  NOR2XL U13790 ( .A(n20896), .B(n20895), .Y(n20978) );
  NOR2XL U13791 ( .A(n20945), .B(n20944), .Y(n20982) );
  AOI21XL U13792 ( .A0(n21281), .A1(n21351), .B0(n21350), .Y(n21405) );
  INVXL U13793 ( .A(n21349), .Y(n21350) );
  NAND2XL U13794 ( .A(n21259), .B(n21281), .Y(n21402) );
  NOR2XL U13795 ( .A(n21355), .B(n21354), .Y(n21404) );
  AOI21XL U13796 ( .A0(n21258), .A1(n21257), .B0(n21256), .Y(n21471) );
  NOR2XL U13797 ( .A(n21246), .B(n21254), .Y(n21257) );
  NAND2XL U13798 ( .A(n21245), .B(n21252), .Y(n21254) );
  AOI21XL U13799 ( .A0(n17832), .A1(n17831), .B0(n17830), .Y(n18034) );
  NOR2XL U13800 ( .A(n17829), .B(n17826), .Y(n17832) );
  NOR2XL U13801 ( .A(n17971), .B(n17970), .Y(n18028) );
  NOR2XL U13802 ( .A(n17895), .B(n17898), .Y(n18025) );
  AOI21XL U13803 ( .A0(n18203), .A1(n18202), .B0(n18201), .Y(n18473) );
  NAND2XL U13804 ( .A(n18197), .B(n18203), .Y(n18464) );
  NOR2XL U13805 ( .A(n18206), .B(n18205), .Y(n18341) );
  NOR2XL U13806 ( .A(n18294), .B(n18293), .Y(n18344) );
  NOR2XL U13807 ( .A(n18349), .B(n18348), .Y(n18462) );
  NOR2XL U13808 ( .A(n18381), .B(n18380), .Y(n18467) );
  NOR2XL U13809 ( .A(n18341), .B(n18344), .Y(n18463) );
  NOR2XL U13810 ( .A(n18539), .B(n18538), .Y(n18564) );
  NOR2XL U13811 ( .A(n20517), .B(n20516), .Y(n20593) );
  NOR2XL U13812 ( .A(n20821), .B(n20820), .Y(n20863) );
  NAND2XL U13813 ( .A(n20797), .B(n20803), .Y(n20805) );
  AOI21XL U13814 ( .A0(n20803), .A1(n20802), .B0(n20801), .Y(n20804) );
  NOR2XL U13815 ( .A(n20796), .B(n20800), .Y(n20803) );
  NOR2XL U13816 ( .A(n20867), .B(n20866), .Y(n21000) );
  NOR2XL U13817 ( .A(n20914), .B(n20913), .Y(n21004) );
  NOR2XL U13818 ( .A(n20860), .B(n20863), .Y(n21001) );
  NOR2XL U13819 ( .A(n21010), .B(n21009), .Y(n21107) );
  NOR2XL U13820 ( .A(n21058), .B(n21057), .Y(n21110) );
  NOR2XL U13821 ( .A(n20484), .B(n20483), .Y(n20525) );
  NAND2XL U13822 ( .A(n28892), .B(U1_pipe1[1]), .Y(n19702) );
  NOR2XL U13823 ( .A(n28892), .B(U1_pipe1[1]), .Y(n19704) );
  NOR2XL U13824 ( .A(n20669), .B(n20668), .Y(n20714) );
  NOR2XL U13825 ( .A(n20619), .B(n20622), .Y(n20711) );
  NOR2XL U13826 ( .A(n20775), .B(n20774), .Y(n20829) );
  NOR2XL U13827 ( .A(n20833), .B(n20832), .Y(n20919) );
  NOR2XL U13828 ( .A(n20874), .B(n20873), .Y(n20923) );
  AOI21XL U13829 ( .A0(n21340), .A1(n21291), .B0(n21339), .Y(n21394) );
  INVXL U13830 ( .A(n21338), .Y(n21339) );
  NAND2XL U13831 ( .A(n21337), .B(n21291), .Y(n21391) );
  NOR2XL U13832 ( .A(n21344), .B(n21343), .Y(n21393) );
  AOI21XL U13833 ( .A0(n21161), .A1(n21160), .B0(n21159), .Y(n21459) );
  NOR2XL U13834 ( .A(n21149), .B(n21157), .Y(n21160) );
  NAND2XL U13835 ( .A(n21148), .B(n21155), .Y(n21157) );
  NOR2X1 U13836 ( .A(n26083), .B(n26082), .Y(n26146) );
  NOR2XL U13837 ( .A(n23227), .B(n23226), .Y(n23271) );
  CMPR32X1 U13838 ( .A(n23982), .B(n23981), .C(U2_A_i_d[16]), .CO(n23983), .S(
        n23939) );
  INVXL U13839 ( .A(n25847), .Y(n20507) );
  INVX1 U13840 ( .A(n26188), .Y(n20854) );
  INVX1 U13841 ( .A(n26355), .Y(n21016) );
  CLKINVX2 U13842 ( .A(n26866), .Y(n21529) );
  ADDFX2 U13843 ( .A(n21616), .B(n21615), .CI(U2_A_r_d[22]), .CO(n21617), .S(
        n21577) );
  INVXL U13844 ( .A(n26948), .Y(n21615) );
  INVXL U13845 ( .A(n23176), .Y(n17789) );
  INVX1 U13846 ( .A(n23365), .Y(n17977) );
  INVXL U13847 ( .A(n23577), .Y(n18189) );
  ADDFX2 U13848 ( .A(n18254), .B(n18253), .CI(U2_A_i_d[10]), .CO(n18255), .S(
        n18191) );
  INVX1 U13849 ( .A(n23690), .Y(n18302) );
  INVX1 U13850 ( .A(n24041), .Y(n18651) );
  INVXL U13851 ( .A(n24332), .Y(n18944) );
  INVXL U13852 ( .A(n24331), .Y(n18943) );
  NOR2XL U13853 ( .A(n24606), .B(n24583), .Y(n25079) );
  AOI21XL U13854 ( .A0(n13510), .A1(n13509), .B0(n13508), .Y(n24920) );
  NOR2XL U13855 ( .A(n14030), .B(U2_A_r_d[8]), .Y(n24930) );
  NOR2XL U13856 ( .A(n14024), .B(U2_A_r_d[5]), .Y(n24951) );
  OR2X2 U13857 ( .A(n24619), .B(n24633), .Y(n24781) );
  INVXL U13858 ( .A(n8900), .Y(n8902) );
  NOR2XL U13859 ( .A(n24440), .B(n7720), .Y(n24430) );
  INVXL U13860 ( .A(n24891), .Y(n24473) );
  NAND2XL U13861 ( .A(n14073), .B(U2_A_r_d[12]), .Y(n24508) );
  NOR2XL U13862 ( .A(n14073), .B(U2_A_r_d[12]), .Y(n13506) );
  NAND2XL U13863 ( .A(n14074), .B(U2_A_r_d[11]), .Y(n24513) );
  NOR2XL U13864 ( .A(n24565), .B(n24559), .Y(n13361) );
  NOR2X1 U13865 ( .A(n9144), .B(n25008), .Y(n9146) );
  INVXL U13866 ( .A(n14465), .Y(n14467) );
  INVXL U13867 ( .A(n14403), .Y(n14405) );
  NAND2XL U13868 ( .A(n14319), .B(n14318), .Y(n14320) );
  NOR2XL U13869 ( .A(n12282), .B(n12281), .Y(n12356) );
  NAND2XL U13870 ( .A(n12282), .B(n12281), .Y(n12355) );
  INVX1 U13871 ( .A(n13103), .Y(n14522) );
  NAND2XL U13872 ( .A(n22897), .B(n13101), .Y(n22092) );
  NOR2X1 U13873 ( .A(n25226), .B(U2_A_i_d[10]), .Y(n22110) );
  INVXL U13874 ( .A(n13150), .Y(n13144) );
  NAND2X1 U13875 ( .A(n22918), .B(n14533), .Y(n22034) );
  AOI21XL U13876 ( .A0(n13117), .A1(n13116), .B0(n13115), .Y(n22362) );
  NOR2X1 U13877 ( .A(n22965), .B(n24687), .Y(n7755) );
  INVX1 U13878 ( .A(n7346), .Y(n22942) );
  NOR2XL U13879 ( .A(n22920), .B(n24621), .Y(n23065) );
  INVXL U13880 ( .A(n13470), .Y(n13472) );
  AOI21XL U13881 ( .A0(n14081), .A1(n14080), .B0(n14079), .Y(n22808) );
  INVX1 U13882 ( .A(n14024), .Y(n14065) );
  XNOR2X1 U13883 ( .A(n9174), .B(n9173), .Y(n24674) );
  NAND2XL U13884 ( .A(n9172), .B(n9177), .Y(n9173) );
  OAI21XL U13885 ( .A0(n9169), .A1(n9175), .B0(n9179), .Y(n9174) );
  INVXL U13886 ( .A(n9178), .Y(n9172) );
  NAND2BX1 U13887 ( .AN(n13167), .B(n24681), .Y(n25311) );
  INVXL U13888 ( .A(n12210), .Y(n12189) );
  INVXL U13889 ( .A(n12205), .Y(n12191) );
  INVXL U13890 ( .A(n12199), .Y(n12201) );
  INVXL U13891 ( .A(n12179), .Y(n12163) );
  INVXL U13892 ( .A(n12149), .Y(n12085) );
  NOR2XL U13893 ( .A(n24583), .B(n13106), .Y(n25762) );
  NAND2XL U13894 ( .A(n12099), .B(n12098), .Y(n12100) );
  NAND2XL U13895 ( .A(n12113), .B(n12112), .Y(n12114) );
  AOI21XL U13896 ( .A0(n12110), .A1(n12109), .B0(n12108), .Y(n12115) );
  NAND2X1 U13897 ( .A(n22594), .B(n7734), .Y(n7210) );
  INVXL U13898 ( .A(n22596), .Y(n7734) );
  INVXL U13899 ( .A(n9113), .Y(n9103) );
  INVXL U13900 ( .A(n12618), .Y(n12594) );
  NAND2X1 U13901 ( .A(n6997), .B(n12572), .Y(n12578) );
  INVXL U13902 ( .A(n12607), .Y(n12609) );
  NAND2XL U13903 ( .A(n9133), .B(n9132), .Y(n9134) );
  INVXL U13904 ( .A(n9131), .Y(n9133) );
  XNOR2X1 U13905 ( .A(n5821), .B(n8964), .Y(n24623) );
  NAND2XL U13906 ( .A(n8828), .B(n8965), .Y(n8829) );
  NAND2XL U13907 ( .A(n24602), .B(n22889), .Y(n22709) );
  OAI21XL U13908 ( .A0(n12510), .A1(n22725), .B0(n12509), .Y(n22707) );
  INVXL U13909 ( .A(n22723), .Y(n12508) );
  INVXL U13910 ( .A(n22718), .Y(n22724) );
  NAND2XL U13911 ( .A(n13496), .B(n13495), .Y(n13497) );
  INVXL U13912 ( .A(n13494), .Y(n13496) );
  INVXL U13913 ( .A(n13421), .Y(n13423) );
  NAND2XL U13914 ( .A(n14031), .B(U2_A_i_d[10]), .Y(n22536) );
  INVXL U13915 ( .A(n13374), .Y(n13315) );
  NOR2XL U13916 ( .A(n14024), .B(U2_A_i_d[5]), .Y(n22556) );
  INVXL U13917 ( .A(n13323), .Y(n13325) );
  NAND2XL U13918 ( .A(n13356), .B(n13355), .Y(n13357) );
  NAND2XL U13919 ( .A(n13344), .B(n13343), .Y(n13345) );
  AOI21XL U13920 ( .A0(n13341), .A1(n13340), .B0(n13339), .Y(n13346) );
  INVXL U13921 ( .A(n13342), .Y(n13344) );
  INVXL U13922 ( .A(n9106), .Y(n9097) );
  XOR2X1 U13923 ( .A(n9001), .B(n9000), .Y(n24620) );
  NAND2XL U13924 ( .A(n8999), .B(n9045), .Y(n9000) );
  INVX1 U13925 ( .A(n14533), .Y(n12378) );
  NAND2XL U13926 ( .A(n8837), .B(n8971), .Y(n8838) );
  INVXL U13927 ( .A(n8972), .Y(n8837) );
  INVX1 U13928 ( .A(n13108), .Y(n14527) );
  INVX1 U13929 ( .A(n13107), .Y(n14526) );
  XNOR2X1 U13930 ( .A(n8816), .B(n8815), .Y(n24582) );
  NAND2XL U13931 ( .A(n8814), .B(n8831), .Y(n8815) );
  INVX1 U13932 ( .A(n13106), .Y(n14525) );
  NAND2XL U13933 ( .A(n8922), .B(n8921), .Y(n8923) );
  INVXL U13934 ( .A(n13102), .Y(n14521) );
  NOR2XL U13935 ( .A(n19968), .B(n19967), .Y(n20145) );
  NOR2XL U13936 ( .A(n19966), .B(n19965), .Y(n20143) );
  NOR2X1 U13937 ( .A(n7893), .B(n14798), .Y(n7892) );
  NOR2XL U13938 ( .A(n13674), .B(U1_A_i_d0[5]), .Y(n17266) );
  OAI21XL U13939 ( .A0(n17278), .A1(n17284), .B0(n17279), .Y(n9572) );
  NOR2XL U13940 ( .A(n13681), .B(U1_A_i_d0[8]), .Y(n17242) );
  AOI21XL U13941 ( .A0(n9580), .A1(n9579), .B0(n9578), .Y(n17233) );
  NAND2X1 U13942 ( .A(n13728), .B(n17199), .Y(n9596) );
  XNOR2X1 U13943 ( .A(n12870), .B(n12869), .Y(n14912) );
  INVXL U13944 ( .A(n12802), .Y(n12804) );
  OAI21XL U13945 ( .A0(n13539), .A1(n17443), .B0(n13538), .Y(n17423) );
  NOR2XL U13946 ( .A(n19518), .B(n14921), .Y(n17410) );
  OAI21XL U13947 ( .A0(n20443), .A1(n20441), .B0(n20444), .Y(n14868) );
  NAND2XL U13948 ( .A(n19567), .B(n20026), .Y(n20337) );
  NAND2XL U13949 ( .A(n13669), .B(U1_A_i_d0[2]), .Y(n17289) );
  NAND2XL U13950 ( .A(n13676), .B(U1_A_i_d0[7]), .Y(n17262) );
  NAND2X1 U13951 ( .A(n9694), .B(n7069), .Y(n17217) );
  XNOR2X1 U13952 ( .A(n12878), .B(n12877), .Y(n19369) );
  NAND2XL U13953 ( .A(n12876), .B(n12875), .Y(n12877) );
  NOR2XL U13954 ( .A(n12884), .B(n19518), .Y(n17706) );
  OAI21XL U13955 ( .A0(n6931), .A1(n7923), .B0(n7921), .Y(n7920) );
  NAND2X1 U13956 ( .A(n7919), .B(n7924), .Y(n7918) );
  INVX1 U13957 ( .A(n19248), .Y(n7171) );
  AOI21XL U13958 ( .A0(n19743), .A1(n19742), .B0(n19741), .Y(n19873) );
  NAND2XL U13959 ( .A(n9391), .B(n9390), .Y(n9392) );
  AOI21XL U13960 ( .A0(n9388), .A1(n9387), .B0(n9386), .Y(n9393) );
  INVXL U13961 ( .A(n9389), .Y(n9391) );
  INVXL U13962 ( .A(n13890), .Y(n13878) );
  AND2X2 U13963 ( .A(n6051), .B(n7721), .Y(n13917) );
  INVXL U13964 ( .A(n13918), .Y(n13906) );
  XOR2X2 U13965 ( .A(n7512), .B(n6994), .Y(n14962) );
  INVXL U13966 ( .A(n8464), .Y(n8466) );
  NAND2XL U13967 ( .A(n7217), .B(n8656), .Y(n16704) );
  AOI21XL U13968 ( .A0(n16700), .A1(n16656), .B0(n16655), .Y(n16668) );
  INVX1 U13969 ( .A(n14901), .Y(n19966) );
  INVX1 U13970 ( .A(n14900), .Y(n19968) );
  NOR2X1 U13971 ( .A(n14922), .B(n19968), .Y(n16898) );
  INVXL U13972 ( .A(n13056), .Y(n13010) );
  NOR2X1 U13973 ( .A(n14962), .B(n20016), .Y(n16800) );
  INVXL U13974 ( .A(n16782), .Y(n7939) );
  NAND2XL U13975 ( .A(n12290), .B(U1_A_r_d0[2]), .Y(n19941) );
  OR2X2 U13976 ( .A(n19734), .B(U1_A_r_d0[12]), .Y(n19878) );
  NAND2X1 U13977 ( .A(n7542), .B(U1_A_r_d0[18]), .Y(n19838) );
  NAND2BXL U13978 ( .AN(n8675), .B(U1_A_r_d0[20]), .Y(n19828) );
  NAND2X1 U13979 ( .A(n19829), .B(n19833), .Y(n12323) );
  NOR2X1 U13980 ( .A(n19237), .B(n20033), .Y(n19564) );
  NAND2XL U13981 ( .A(n13669), .B(U1_A_r_d0[2]), .Y(n19222) );
  NOR2X1 U13982 ( .A(n19154), .B(n9684), .Y(n9686) );
  NAND2XL U13983 ( .A(n6953), .B(n19156), .Y(n9684) );
  AOI21XL U13984 ( .A0(n19150), .A1(n19103), .B0(n19102), .Y(n19116) );
  INVX1 U13985 ( .A(n19967), .Y(n7357) );
  NOR2X1 U13986 ( .A(n7357), .B(n19519), .Y(n19344) );
  NOR2XL U13987 ( .A(n14754), .B(n19518), .Y(n19342) );
  NAND2XL U13988 ( .A(n14790), .B(n14773), .Y(n19303) );
  INVXL U13989 ( .A(n14817), .Y(n14819) );
  NAND2X1 U13990 ( .A(n14834), .B(n19268), .Y(n19257) );
  NOR2X1 U13991 ( .A(n14832), .B(n19276), .Y(n7204) );
  NAND2XL U13992 ( .A(n8505), .B(n8504), .Y(n8506) );
  INVXL U13993 ( .A(n8503), .Y(n8505) );
  NAND2XL U13994 ( .A(n12290), .B(U1_A_i_d0[2]), .Y(n16771) );
  NAND2XL U13995 ( .A(n8490), .B(n8489), .Y(n8491) );
  INVXL U13996 ( .A(n8601), .Y(n8603) );
  NAND2X1 U13997 ( .A(n7542), .B(U1_A_i_d0[18]), .Y(n16670) );
  INVXL U13998 ( .A(n8592), .Y(n8593) );
  NAND2XL U13999 ( .A(n7301), .B(U1_A_i_d0[20]), .Y(n16661) );
  NAND2XL U14000 ( .A(n12332), .B(U1_A_i_d0[24]), .Y(n16636) );
  NAND2XL U14001 ( .A(n13828), .B(n13827), .Y(n13829) );
  AOI21XL U14002 ( .A0(n13825), .A1(n13822), .B0(n13824), .Y(n13830) );
  INVXL U14003 ( .A(n13826), .Y(n13828) );
  NAND2XL U14004 ( .A(n12819), .B(n12818), .Y(n12820) );
  NAND2XL U14005 ( .A(n12915), .B(n12938), .Y(n12916) );
  NOR2XL U14006 ( .A(n13674), .B(U1_A_r_d0[5]), .Y(n19203) );
  NOR2X1 U14007 ( .A(n13675), .B(U1_A_r_d0[6]), .Y(n19197) );
  NAND2X1 U14008 ( .A(n9694), .B(n7070), .Y(n19134) );
  NAND2XL U14009 ( .A(n13710), .B(U1_A_r_d0[22]), .Y(n19093) );
  NOR2X1 U14010 ( .A(n19519), .B(n19967), .Y(n19673) );
  NOR2XL U14011 ( .A(n19518), .B(n19965), .Y(n19671) );
  XOR2X1 U14012 ( .A(n12929), .B(n12794), .Y(n19520) );
  INVXL U14013 ( .A(n12928), .Y(n12793) );
  AOI21XL U14014 ( .A0(n19684), .A1(n19517), .B0(n19516), .Y(n19664) );
  INVXL U14015 ( .A(n14779), .Y(n14781) );
  NAND2XL U14016 ( .A(n12960), .B(n12995), .Y(n12961) );
  INVXL U14017 ( .A(n12992), .Y(n12960) );
  NAND2XL U14018 ( .A(n12954), .B(n12994), .Y(n12955) );
  INVX1 U14019 ( .A(n19281), .Y(n19548) );
  INVXL U14020 ( .A(n14798), .Y(n14799) );
  NAND3X1 U14021 ( .A(n7500), .B(n7499), .C(n13075), .Y(n7498) );
  INVXL U14022 ( .A(n13569), .Y(n13075) );
  NAND2XL U14023 ( .A(n19552), .B(n19538), .Y(n19596) );
  NOR2X1 U14024 ( .A(n19551), .B(n7791), .Y(n19597) );
  NOR2X1 U14025 ( .A(n7792), .B(n19609), .Y(n7791) );
  XOR2X2 U14026 ( .A(n7190), .B(n13576), .Y(n19557) );
  NAND2XL U14027 ( .A(n9377), .B(n9376), .Y(n9378) );
  NAND3X1 U14028 ( .A(n5922), .B(n28675), .C(n28707), .Y(n14981) );
  NAND2XL U14029 ( .A(CQ0[9]), .B(n27814), .Y(n27851) );
  NAND2XL U14030 ( .A(CQ0[7]), .B(n27814), .Y(n27843) );
  NAND2XL U14031 ( .A(CQ0[6]), .B(n27814), .Y(n27839) );
  NAND2XL U14032 ( .A(CQ0[5]), .B(n27814), .Y(n27835) );
  NAND2XL U14033 ( .A(CQ0[51]), .B(n27814), .Y(n28051) );
  INVXL U14034 ( .A(n28051), .Y(n28053) );
  NAND2XL U14035 ( .A(n27814), .B(n28051), .Y(n28052) );
  NAND2XL U14036 ( .A(CQ0[50]), .B(n27814), .Y(n28045) );
  INVXL U14037 ( .A(n28045), .Y(n28047) );
  NAND2XL U14038 ( .A(n28921), .B(n28045), .Y(n28046) );
  NAND2XL U14039 ( .A(CQ0[4]), .B(n27814), .Y(n27831) );
  NAND2XL U14040 ( .A(n27814), .B(n28040), .Y(n28041) );
  NAND2XL U14041 ( .A(CQ0[48]), .B(n27814), .Y(n28035) );
  INVXL U14042 ( .A(n28035), .Y(n28037) );
  NAND2XL U14043 ( .A(n27814), .B(n28035), .Y(n28036) );
  NAND2XL U14044 ( .A(CQ0[46]), .B(n27814), .Y(n28025) );
  INVXL U14045 ( .A(n28025), .Y(n28027) );
  NAND2XL U14046 ( .A(n28921), .B(n28025), .Y(n28026) );
  INVXL U14047 ( .A(n28020), .Y(n28022) );
  NAND2XL U14048 ( .A(n27814), .B(n28020), .Y(n28021) );
  NAND2XL U14049 ( .A(CQ0[45]), .B(n27814), .Y(n28020) );
  NAND2XL U14050 ( .A(CQ0[44]), .B(n27814), .Y(n28015) );
  INVXL U14051 ( .A(n28015), .Y(n28017) );
  NAND2XL U14052 ( .A(n28921), .B(n28015), .Y(n28016) );
  NAND2XL U14053 ( .A(CQ0[43]), .B(n27814), .Y(n28010) );
  INVXL U14054 ( .A(n28010), .Y(n28012) );
  NAND2XL U14055 ( .A(n28921), .B(n28010), .Y(n28011) );
  INVXL U14056 ( .A(n28000), .Y(n28002) );
  NAND2XL U14057 ( .A(n28921), .B(n28000), .Y(n28001) );
  NAND2XL U14058 ( .A(CQ0[41]), .B(n27814), .Y(n28000) );
  NAND2XL U14059 ( .A(CQ0[40]), .B(n27814), .Y(n27995) );
  INVXL U14060 ( .A(n27995), .Y(n27997) );
  NAND2XL U14061 ( .A(n28921), .B(n27995), .Y(n27996) );
  NAND2XL U14062 ( .A(CQ0[3]), .B(n27814), .Y(n27827) );
  NAND2XL U14063 ( .A(CQ0[39]), .B(n27814), .Y(n27990) );
  INVXL U14064 ( .A(n27990), .Y(n27992) );
  NAND2XL U14065 ( .A(n27814), .B(n27990), .Y(n27991) );
  NAND2XL U14066 ( .A(CQ0[36]), .B(n27814), .Y(n27975) );
  NAND2XL U14067 ( .A(CQ0[35]), .B(n27814), .Y(n27971) );
  NAND2XL U14068 ( .A(CQ0[34]), .B(n27814), .Y(n27967) );
  NAND2XL U14069 ( .A(CQ0[32]), .B(n27814), .Y(n27958) );
  NAND2XL U14070 ( .A(CQ0[31]), .B(n27814), .Y(n27954) );
  NAND2XL U14071 ( .A(CQ0[30]), .B(n27814), .Y(n27950) );
  NAND2XL U14072 ( .A(CQ0[2]), .B(n27814), .Y(n27823) );
  NAND2XL U14073 ( .A(CQ0[29]), .B(n27814), .Y(n27946) );
  NAND2XL U14074 ( .A(CQ0[27]), .B(n27814), .Y(n27938) );
  NAND2XL U14075 ( .A(CQ0[25]), .B(n27814), .Y(n27929) );
  INVXL U14076 ( .A(n27929), .Y(n27931) );
  NAND2XL U14077 ( .A(n28921), .B(n27929), .Y(n27930) );
  NAND2XL U14078 ( .A(CQ0[24]), .B(n27814), .Y(n27924) );
  INVXL U14079 ( .A(n27924), .Y(n27926) );
  NAND2XL U14080 ( .A(n28921), .B(n27924), .Y(n27925) );
  NAND2XL U14081 ( .A(n27814), .B(n27919), .Y(n27920) );
  INVXL U14082 ( .A(n27914), .Y(n27916) );
  NAND2XL U14083 ( .A(n28921), .B(n27914), .Y(n27915) );
  NAND2XL U14084 ( .A(CQ0[22]), .B(n27814), .Y(n27914) );
  NAND2XL U14085 ( .A(CQ0[21]), .B(n27814), .Y(n27909) );
  INVXL U14086 ( .A(n27909), .Y(n27911) );
  NAND2XL U14087 ( .A(n28921), .B(n27909), .Y(n27910) );
  NAND2XL U14088 ( .A(n27814), .B(n27904), .Y(n27905) );
  NAND2XL U14089 ( .A(CQ0[1]), .B(n27814), .Y(n27819) );
  NAND2XL U14090 ( .A(CQ0[19]), .B(n27814), .Y(n27899) );
  INVXL U14091 ( .A(n27899), .Y(n27901) );
  NAND2XL U14092 ( .A(n27814), .B(n27899), .Y(n27900) );
  NAND2XL U14093 ( .A(CQ0[18]), .B(n27814), .Y(n27894) );
  INVXL U14094 ( .A(n27894), .Y(n27896) );
  NAND2XL U14095 ( .A(n28921), .B(n27894), .Y(n27895) );
  NAND2XL U14096 ( .A(CQ0[17]), .B(n27814), .Y(n27889) );
  INVXL U14097 ( .A(n27889), .Y(n27891) );
  NAND2XL U14098 ( .A(n28921), .B(n27889), .Y(n27890) );
  NAND2XL U14099 ( .A(CQ0[16]), .B(n27814), .Y(n27884) );
  INVXL U14100 ( .A(n27884), .Y(n27886) );
  NAND2XL U14101 ( .A(n27814), .B(n27884), .Y(n27885) );
  NAND2XL U14102 ( .A(CQ0[14]), .B(n27814), .Y(n27874) );
  INVXL U14103 ( .A(n27874), .Y(n27876) );
  NAND2XL U14104 ( .A(n27814), .B(n27874), .Y(n27875) );
  NAND2XL U14105 ( .A(CQ0[12]), .B(n27814), .Y(n27864) );
  INVXL U14106 ( .A(n27864), .Y(n27866) );
  NAND2XL U14107 ( .A(n28921), .B(n27864), .Y(n27865) );
  NAND2XL U14108 ( .A(CQ0[11]), .B(n27814), .Y(n27859) );
  INVXL U14109 ( .A(n27859), .Y(n27861) );
  NAND2XL U14110 ( .A(n28921), .B(n27859), .Y(n27860) );
  NAND2XL U14111 ( .A(CQ0[10]), .B(n27814), .Y(n27855) );
  NAND2XL U14112 ( .A(CQ0[0]), .B(n27814), .Y(n27815) );
  NAND2BX1 U14113 ( .AN(n11613), .B(n11633), .Y(n11625) );
  INVXL U14114 ( .A(n11911), .Y(n28640) );
  XNOR2X1 U14115 ( .A(n8194), .B(BOPC[26]), .Y(U1_U1_z0[0]) );
  XNOR2X1 U14116 ( .A(n8206), .B(AOPC[26]), .Y(U0_U1_z0[0]) );
  AOI22XL U14117 ( .A0(B4_q[35]), .A1(n7126), .B0(B7_q[35]), .B1(n7127), .Y(
        n15009) );
  AOI22XL U14118 ( .A0(B7_q[37]), .A1(n7127), .B0(B6_q[37]), .B1(n16570), .Y(
        n15326) );
  AOI22XL U14119 ( .A0(B4_q[42]), .A1(n7126), .B0(B6_q[42]), .B1(n16570), .Y(
        n15288) );
  AOI22XL U14120 ( .A0(B7_q[16]), .A1(n16325), .B0(B5_q[16]), .B1(n16344), .Y(
        n15707) );
  AOI22XL U14121 ( .A0(B7_q[16]), .A1(n15982), .B0(B6_q[16]), .B1(n15958), .Y(
        n15913) );
  AOI22XL U14122 ( .A0(B7_q[15]), .A1(n16158), .B0(B4_q[15]), .B1(n15557), .Y(
        n15520) );
  AOI22XL U14123 ( .A0(B6_q[19]), .A1(n5926), .B0(B7_q[19]), .B1(n16325), .Y(
        n15695) );
  AOI22XL U14124 ( .A0(B4_q[11]), .A1(n15557), .B0(B6_q[11]), .B1(n16143), .Y(
        n15535) );
  INVXL U14125 ( .A(B6_q[13]), .Y(n15721) );
  AOI22XL U14126 ( .A0(B6_q[29]), .A1(n15958), .B0(B5_q[29]), .B1(n15963), .Y(
        n15861) );
  AOI22XL U14127 ( .A0(B6_q[5]), .A1(n16293), .B0(B7_q[5]), .B1(n16325), .Y(
        n15752) );
  INVXL U14128 ( .A(B3_q[35]), .Y(n16226) );
  INVXL U14129 ( .A(B2_q[26]), .Y(n15127) );
  INVXL U14130 ( .A(B3_q[37]), .Y(n16034) );
  AOI22XL U14131 ( .A0(B6_q[29]), .A1(n5926), .B0(B5_q[29]), .B1(n16344), .Y(
        n15658) );
  INVXL U14132 ( .A(B7_q[43]), .Y(n15610) );
  AOI22XL U14133 ( .A0(B6_q[37]), .A1(n16293), .B0(B7_q[37]), .B1(n16325), .Y(
        n15629) );
  AOI22XL U14134 ( .A0(B5_q[27]), .A1(n16344), .B0(B7_q[27]), .B1(n16325), .Y(
        n15666) );
  AOI22XL U14135 ( .A0(B6_q[27]), .A1(n15958), .B0(B5_q[27]), .B1(n15963), .Y(
        n15869) );
  AOI22XL U14136 ( .A0(B2_q[27]), .A1(n15958), .B0(B0_q[27]), .B1(n5925), .Y(
        n15121) );
  AOI22XL U14137 ( .A0(B3_q[32]), .A1(n5930), .B0(B0_q[32]), .B1(n5925), .Y(
        n15104) );
  AOI22XL U14138 ( .A0(B3_q[32]), .A1(n16158), .B0(B2_q[32]), .B1(n15431), .Y(
        n16050) );
  INVXL U14139 ( .A(B7_q[32]), .Y(n15851) );
  INVXL U14140 ( .A(B4_q[0]), .Y(n15387) );
  INVXL U14141 ( .A(n19240), .Y(n19241) );
  XOR2X1 U14142 ( .A(n7808), .B(n14689), .Y(n19567) );
  INVXL U14143 ( .A(n25299), .Y(n25300) );
  INVXL U14144 ( .A(n25298), .Y(n25301) );
  INVXL U14145 ( .A(n20037), .Y(n20040) );
  NAND2XL U14146 ( .A(n19239), .B(n14855), .Y(n19236) );
  INVXL U14147 ( .A(n20329), .Y(n7896) );
  INVXL U14148 ( .A(n14107), .Y(n7214) );
  INVXL U14149 ( .A(n22602), .Y(n22604) );
  OR2X2 U14150 ( .A(n19259), .B(n14960), .Y(n17330) );
  NAND2XL U14151 ( .A(n24735), .B(n24734), .Y(n25012) );
  INVX1 U14152 ( .A(n20330), .Y(n7337) );
  NAND2XL U14153 ( .A(n19553), .B(n14835), .Y(n19262) );
  AOI22XL U14154 ( .A0(B7_q[35]), .A1(n16325), .B0(B5_q[35]), .B1(n16344), .Y(
        n15637) );
  AOI22XL U14155 ( .A0(B6_q[37]), .A1(n16143), .B0(B4_q[37]), .B1(n15557), .Y(
        n15440) );
  AOI22XL U14156 ( .A0(B5_q[38]), .A1(n16344), .B0(B7_q[38]), .B1(n16325), .Y(
        n15625) );
  AOI22XL U14157 ( .A0(B4_q[44]), .A1(n15687), .B0(B6_q[44]), .B1(n5926), .Y(
        n15604) );
  AOI22XL U14158 ( .A0(B1_q[31]), .A1(n16344), .B0(B3_q[31]), .B1(n16325), .Y(
        n16238) );
  AOI22XL U14159 ( .A0(B3_q[31]), .A1(n16158), .B0(B2_q[31]), .B1(n16161), .Y(
        n16054) );
  INVXL U14160 ( .A(B3_q[33]), .Y(n16048) );
  AOI22XL U14161 ( .A0(B1_q[31]), .A1(n15963), .B0(B2_q[31]), .B1(n15958), .Y(
        n15108) );
  INVXL U14162 ( .A(B7_q[36]), .Y(n15446) );
  INVXL U14163 ( .A(B3_q[38]), .Y(n16215) );
  AOI22XL U14164 ( .A0(B7_q[5]), .A1(n7127), .B0(B6_q[5]), .B1(n16570), .Y(
        n15361) );
  AOI22XL U14165 ( .A0(B7_q[6]), .A1(n7127), .B0(B6_q[6]), .B1(n16570), .Y(
        n15354) );
  INVXL U14166 ( .A(B4_q[7]), .Y(n15352) );
  AOI22XL U14167 ( .A0(B4_q[2]), .A1(n7126), .B0(B7_q[2]), .B1(n7127), .Y(
        n15378) );
  NOR2XL U14168 ( .A(n7315), .B(n17176), .Y(n7318) );
  NOR2XL U14169 ( .A(n7654), .B(n9548), .Y(n7651) );
  INVXL U14170 ( .A(B4_q[47]), .Y(n15252) );
  INVXL U14171 ( .A(B4_q[45]), .Y(n15268) );
  AOI22XL U14172 ( .A0(B4_q[46]), .A1(n7126), .B0(B6_q[46]), .B1(n16570), .Y(
        n15258) );
  INVXL U14173 ( .A(B3_q[0]), .Y(n16168) );
  INVXL U14174 ( .A(B0_q[0]), .Y(n16573) );
  INVXL U14175 ( .A(B3_q[10]), .Y(n15185) );
  INVXL U14176 ( .A(B2_q[12]), .Y(n15177) );
  INVXL U14177 ( .A(B3_q[13]), .Y(n15173) );
  INVXL U14178 ( .A(B0_q[14]), .Y(n16515) );
  AOI22XL U14179 ( .A0(B2_q[15]), .A1(n15958), .B0(B3_q[15]), .B1(n5930), .Y(
        n15166) );
  INVXL U14180 ( .A(B2_q[15]), .Y(n16299) );
  INVXL U14181 ( .A(B1_q[15]), .Y(n16111) );
  INVXL U14182 ( .A(B3_q[16]), .Y(n16107) );
  INVXL U14183 ( .A(B1_q[16]), .Y(n16508) );
  AOI22XL U14184 ( .A0(B2_q[17]), .A1(n15958), .B0(B3_q[17]), .B1(n5930), .Y(
        n15157) );
  AOI22XL U14185 ( .A0(B3_q[17]), .A1(n16325), .B0(B0_q[17]), .B1(n15687), .Y(
        n16289) );
  AOI22XL U14186 ( .A0(B2_q[17]), .A1(n16161), .B0(B0_q[17]), .B1(n15557), .Y(
        n16101) );
  INVXL U14187 ( .A(B0_q[18]), .Y(n16499) );
  AOI22XL U14188 ( .A0(B3_q[1]), .A1(n5930), .B0(B2_q[1]), .B1(n15214), .Y(
        n15215) );
  AOI22XL U14189 ( .A0(B0_q[1]), .A1(n15687), .B0(B2_q[1]), .B1(n16354), .Y(
        n16350) );
  AOI22XL U14190 ( .A0(B3_q[1]), .A1(n16158), .B0(B0_q[1]), .B1(n5933), .Y(
        n16159) );
  AOI22XL U14191 ( .A0(B3_q[20]), .A1(n5930), .B0(B2_q[20]), .B1(n15958), .Y(
        n15147) );
  AOI22XL U14192 ( .A0(B3_q[20]), .A1(n16325), .B0(B1_q[20]), .B1(n16344), .Y(
        n16278) );
  AOI22XL U14193 ( .A0(B2_q[20]), .A1(n16161), .B0(B1_q[20]), .B1(n16165), .Y(
        n16091) );
  INVXL U14194 ( .A(B0_q[20]), .Y(n16490) );
  INVXL U14195 ( .A(B3_q[21]), .Y(n15145) );
  INVXL U14196 ( .A(B3_q[22]), .Y(n16086) );
  INVXL U14197 ( .A(B1_q[22]), .Y(n16481) );
  INVXL U14198 ( .A(B3_q[23]), .Y(n15138) );
  INVXL U14199 ( .A(B3_q[25]), .Y(n16263) );
  INVXL U14200 ( .A(B3_q[26]), .Y(n16259) );
  INVXL U14201 ( .A(B0_q[26]), .Y(n16464) );
  AOI22XL U14202 ( .A0(B1_q[27]), .A1(n16344), .B0(B3_q[27]), .B1(n16325), .Y(
        n16253) );
  AOI22XL U14203 ( .A0(B3_q[27]), .A1(n16158), .B0(B2_q[27]), .B1(n15431), .Y(
        n16068) );
  INVXL U14204 ( .A(B1_q[27]), .Y(n16459) );
  INVXL U14205 ( .A(B0_q[28]), .Y(n16455) );
  INVXL U14206 ( .A(B2_q[29]), .Y(n16063) );
  INVXL U14207 ( .A(B2_q[2]), .Y(n15212) );
  INVXL U14208 ( .A(B3_q[2]), .Y(n16347) );
  INVXL U14209 ( .A(B0_q[2]), .Y(n16562) );
  INVXL U14210 ( .A(B0_q[31]), .Y(n16443) );
  AOI22XL U14211 ( .A0(B2_q[32]), .A1(n5926), .B0(B0_q[32]), .B1(n15687), .Y(
        n16234) );
  AOI22XL U14212 ( .A0(B2_q[36]), .A1(n15958), .B0(B3_q[36]), .B1(n5930), .Y(
        n15091) );
  AOI22XL U14213 ( .A0(B2_q[36]), .A1(n5926), .B0(B1_q[36]), .B1(n16344), .Y(
        n16220) );
  AOI22XL U14214 ( .A0(B3_q[36]), .A1(n16158), .B0(B1_q[36]), .B1(n16165), .Y(
        n16036) );
  INVXL U14215 ( .A(B0_q[36]), .Y(n16423) );
  INVXL U14216 ( .A(B2_q[3]), .Y(n15208) );
  INVXL U14217 ( .A(B0_q[41]), .Y(n16402) );
  AOI22XL U14218 ( .A0(B2_q[43]), .A1(n15958), .B0(B1_q[43]), .B1(n15963), .Y(
        n15069) );
  AOI22XL U14219 ( .A0(B2_q[43]), .A1(n16354), .B0(B3_q[43]), .B1(n16325), .Y(
        n16196) );
  AOI22XL U14220 ( .A0(B3_q[43]), .A1(n16158), .B0(B1_q[43]), .B1(n16165), .Y(
        n16013) );
  INVXL U14221 ( .A(B0_q[43]), .Y(n16394) );
  INVXL U14222 ( .A(B3_q[45]), .Y(n16191) );
  INVXL U14223 ( .A(B0_q[45]), .Y(n16386) );
  AOI22XL U14224 ( .A0(B2_q[46]), .A1(n15958), .B0(B3_q[46]), .B1(n5930), .Y(
        n15059) );
  AOI22XL U14225 ( .A0(B0_q[46]), .A1(n15687), .B0(B3_q[46]), .B1(n16325), .Y(
        n16185) );
  AOI22XL U14226 ( .A0(B0_q[46]), .A1(n15557), .B0(B2_q[46]), .B1(n16143), .Y(
        n16003) );
  INVXL U14227 ( .A(B3_q[48]), .Y(n15054) );
  INVXL U14228 ( .A(B3_q[49]), .Y(n15995) );
  INVXL U14229 ( .A(B3_q[4]), .Y(n16338) );
  INVXL U14230 ( .A(B2_q[4]), .Y(n16149) );
  INVXL U14231 ( .A(B0_q[4]), .Y(n16554) );
  INVXL U14232 ( .A(B3_q[50]), .Y(n15047) );
  INVXL U14233 ( .A(B2_q[51]), .Y(n15043) );
  INVXL U14234 ( .A(B2_q[6]), .Y(n16331) );
  INVXL U14235 ( .A(B1_q[6]), .Y(n16141) );
  INVXL U14236 ( .A(B0_q[8]), .Y(n16539) );
  INVXL U14237 ( .A(B3_q[9]), .Y(n15189) );
  INVXL U14238 ( .A(B1_q[9]), .Y(n16319) );
  INVXL U14239 ( .A(B0_q[9]), .Y(n16535) );
  NAND2XL U14240 ( .A(n25869), .B(n25868), .Y(n25959) );
  AOI21XL U14241 ( .A0(n27015), .A1(n26973), .B0(n27014), .Y(n27059) );
  INVXL U14242 ( .A(n27013), .Y(n27014) );
  NOR2XL U14243 ( .A(n27017), .B(n27016), .Y(n27058) );
  NAND2XL U14244 ( .A(n27017), .B(n27016), .Y(n27057) );
  NAND2XL U14245 ( .A(n26800), .B(n26799), .Y(n26843) );
  NAND2XL U14246 ( .A(n26791), .B(n26736), .Y(n26796) );
  AOI21XL U14247 ( .A0(n26794), .A1(n26736), .B0(n26793), .Y(n26795) );
  INVXL U14248 ( .A(n26792), .Y(n26793) );
  NOR2XL U14249 ( .A(n26731), .B(n26733), .Y(n26791) );
  NAND2XL U14250 ( .A(n26738), .B(n26737), .Y(n26792) );
  NAND2XL U14251 ( .A(n26682), .B(n26681), .Y(n26732) );
  NAND2XL U14252 ( .A(n26105), .B(n26104), .Y(n26167) );
  INVXL U14253 ( .A(n26169), .Y(n26106) );
  NOR2XL U14254 ( .A(n26061), .B(n26060), .Y(n26166) );
  INVXL U14255 ( .A(n26498), .Y(n26264) );
  NAND2XL U14256 ( .A(n26061), .B(n26060), .Y(n26168) );
  NAND2XL U14257 ( .A(n26005), .B(n26004), .Y(n26051) );
  INVXL U14258 ( .A(n26053), .Y(n26006) );
  NOR2XL U14259 ( .A(n25963), .B(n25962), .Y(n26049) );
  AOI21XL U14260 ( .A0(n25961), .A1(n26050), .B0(n26055), .Y(n26003) );
  NAND2XL U14261 ( .A(n25963), .B(n25962), .Y(n26052) );
  INVXL U14262 ( .A(n25957), .Y(n25907) );
  INVXL U14263 ( .A(n25959), .Y(n25906) );
  NAND2XL U14264 ( .A(n25909), .B(n25908), .Y(n25958) );
  INVXL U14265 ( .A(n25960), .Y(n25910) );
  INVXL U14266 ( .A(n26059), .Y(n25961) );
  NAND2XL U14267 ( .A(n25816), .B(n25815), .Y(n25862) );
  INVXL U14268 ( .A(n25864), .Y(n25817) );
  NAND2XL U14269 ( .A(n26395), .B(n26394), .Y(n26443) );
  NAND2XL U14270 ( .A(n26321), .B(n26320), .Y(n26444) );
  INVXL U14271 ( .A(n26393), .Y(n26448) );
  NAND2XL U14272 ( .A(n26161), .B(n26160), .Y(n26226) );
  INVXL U14273 ( .A(n26228), .Y(n26162) );
  NOR2XL U14274 ( .A(n26138), .B(n26137), .Y(n26225) );
  INVXL U14275 ( .A(n26557), .Y(n26319) );
  NAND2XL U14276 ( .A(n26138), .B(n26137), .Y(n26227) );
  NAND2XL U14277 ( .A(n26044), .B(n26043), .Y(n26128) );
  INVXL U14278 ( .A(n26130), .Y(n26045) );
  NOR2XL U14279 ( .A(n25999), .B(n25998), .Y(n26126) );
  AOI21XL U14280 ( .A0(n25997), .A1(n26127), .B0(n26132), .Y(n26042) );
  NAND2XL U14281 ( .A(n25999), .B(n25998), .Y(n26129) );
  NAND2XL U14282 ( .A(n25881), .B(n25880), .Y(n25926) );
  INVXL U14283 ( .A(n25928), .Y(n25882) );
  NOR2XL U14284 ( .A(n25810), .B(n25809), .Y(n25925) );
  INVXL U14285 ( .A(n25930), .Y(n25879) );
  NAND2XL U14286 ( .A(n25810), .B(n25809), .Y(n25927) );
  AOI21XL U14287 ( .A0(n24857), .A1(n24856), .B0(n24855), .Y(n25808) );
  OR2XL U14288 ( .A(U0_pipe3[1]), .B(U0_pipe2[1]), .Y(n24857) );
  AND2XL U14289 ( .A(U0_pipe3[1]), .B(U0_pipe2[1]), .Y(n24855) );
  OR2XL U14290 ( .A(n28905), .B(U0_pipe2[0]), .Y(n24856) );
  NOR2XL U14291 ( .A(n24853), .B(n28897), .Y(n25807) );
  NAND2XL U14292 ( .A(n24853), .B(n28897), .Y(n25806) );
  AOI21XL U14293 ( .A0(n24348), .A1(n24306), .B0(n24347), .Y(n24404) );
  INVXL U14294 ( .A(n24346), .Y(n24347) );
  NOR2XL U14295 ( .A(n24350), .B(n24349), .Y(n24403) );
  NAND2XL U14296 ( .A(n24350), .B(n24349), .Y(n24402) );
  AOI21XL U14297 ( .A0(n24193), .A1(n24124), .B0(n24192), .Y(n24238) );
  INVXL U14298 ( .A(n24191), .Y(n24192) );
  NOR2XL U14299 ( .A(n24080), .B(n24082), .Y(n24117) );
  NAND2XL U14300 ( .A(n24087), .B(n24086), .Y(n24118) );
  NAND2XL U14301 ( .A(n24007), .B(n24006), .Y(n24081) );
  INVXL U14302 ( .A(n23730), .Y(n23654) );
  NAND2XL U14303 ( .A(n23658), .B(n23657), .Y(n23729) );
  INVXL U14304 ( .A(n23731), .Y(n23659) );
  NAND2XL U14305 ( .A(n23592), .B(n23591), .Y(n23730) );
  INVXL U14306 ( .A(n23728), .Y(n23655) );
  NAND2XL U14307 ( .A(n23437), .B(n23436), .Y(n23515) );
  INVXL U14308 ( .A(n23517), .Y(n23438) );
  NOR2XL U14309 ( .A(n23423), .B(n23422), .Y(n23514) );
  INVXL U14310 ( .A(n23824), .Y(n23590) );
  NAND2XL U14311 ( .A(n23423), .B(n23422), .Y(n23516) );
  NAND2XL U14312 ( .A(n23355), .B(n23354), .Y(n23413) );
  INVXL U14313 ( .A(n23415), .Y(n23356) );
  NOR2XL U14314 ( .A(n23315), .B(n23314), .Y(n23411) );
  AOI21XL U14315 ( .A0(n23313), .A1(n23412), .B0(n23417), .Y(n23353) );
  NAND2XL U14316 ( .A(n23315), .B(n23314), .Y(n23414) );
  INVXL U14317 ( .A(n23311), .Y(n23232) );
  NAND2XL U14318 ( .A(n23235), .B(n23234), .Y(n23310) );
  INVXL U14319 ( .A(n23312), .Y(n23236) );
  NAND2XL U14320 ( .A(n23191), .B(n23190), .Y(n23311) );
  INVXL U14321 ( .A(n23421), .Y(n23313) );
  INVXL U14322 ( .A(n23309), .Y(n23233) );
  NAND2XL U14323 ( .A(n23139), .B(n23138), .Y(n23184) );
  INVXL U14324 ( .A(n23186), .Y(n23140) );
  NOR2XL U14325 ( .A(n23127), .B(U0_pipe10[1]), .Y(n23183) );
  INVXL U14326 ( .A(n23188), .Y(n23137) );
  NAND2XL U14327 ( .A(n23127), .B(U0_pipe10[1]), .Y(n23185) );
  AOI21XL U14328 ( .A0(n27023), .A1(n26981), .B0(n27022), .Y(n27066) );
  INVXL U14329 ( .A(n27021), .Y(n27022) );
  NOR2XL U14330 ( .A(n27025), .B(n27024), .Y(n27065) );
  NAND2XL U14331 ( .A(n27025), .B(n27024), .Y(n27064) );
  INVXL U14332 ( .A(n26922), .Y(n26923) );
  NOR2XL U14333 ( .A(n26926), .B(n26925), .Y(n26979) );
  NAND2XL U14334 ( .A(n26926), .B(n26925), .Y(n26978) );
  AOI21XL U14335 ( .A0(n26837), .A1(n26786), .B0(n26836), .Y(n26882) );
  INVXL U14336 ( .A(n26835), .Y(n26836) );
  NAND2XL U14337 ( .A(n26183), .B(n26182), .Y(n26197) );
  INVXL U14338 ( .A(n26199), .Y(n26184) );
  NOR2XL U14339 ( .A(n26100), .B(n26099), .Y(n26196) );
  INVXL U14340 ( .A(n26585), .Y(n26341) );
  NAND2XL U14341 ( .A(n26100), .B(n26099), .Y(n26198) );
  NAND2XL U14342 ( .A(n26074), .B(n26073), .Y(n26090) );
  INVXL U14343 ( .A(n26092), .Y(n26075) );
  NOR2XL U14344 ( .A(n26026), .B(n26025), .Y(n26088) );
  AOI21XL U14345 ( .A0(n26024), .A1(n26089), .B0(n26094), .Y(n26072) );
  NAND2XL U14346 ( .A(n26026), .B(n26025), .Y(n26091) );
  NAND2XL U14347 ( .A(n25856), .B(n25855), .Y(n25896) );
  INVXL U14348 ( .A(n25898), .Y(n25857) );
  NOR2XL U14349 ( .A(n25833), .B(n25832), .Y(n25895) );
  INVXL U14350 ( .A(n25900), .Y(n25854) );
  NAND2XL U14351 ( .A(n25833), .B(n25832), .Y(n25897) );
  AOI21XL U14352 ( .A0(n24356), .A1(n24314), .B0(n24355), .Y(n24397) );
  INVXL U14353 ( .A(n24354), .Y(n24355) );
  NOR2XL U14354 ( .A(n24358), .B(n24357), .Y(n24396) );
  NAND2XL U14355 ( .A(n24358), .B(n24357), .Y(n24395) );
  AOI21XL U14356 ( .A0(n24185), .A1(n24137), .B0(n24184), .Y(n24230) );
  INVXL U14357 ( .A(n24183), .Y(n24184) );
  NOR2XL U14358 ( .A(n24069), .B(n24071), .Y(n24130) );
  NAND2XL U14359 ( .A(n24076), .B(n24075), .Y(n24131) );
  NAND2XL U14360 ( .A(n24019), .B(n24018), .Y(n24070) );
  INVXL U14361 ( .A(n23719), .Y(n23663) );
  NAND2XL U14362 ( .A(n23667), .B(n23666), .Y(n23718) );
  INVXL U14363 ( .A(n23720), .Y(n23668) );
  NAND2XL U14364 ( .A(n23605), .B(n23604), .Y(n23719) );
  INVXL U14365 ( .A(n23717), .Y(n23664) );
  NAND2XL U14366 ( .A(n23443), .B(n23442), .Y(n23499) );
  INVXL U14367 ( .A(n23501), .Y(n23444) );
  NOR2XL U14368 ( .A(n23400), .B(n23399), .Y(n23498) );
  INVXL U14369 ( .A(n23843), .Y(n23603) );
  NAND2XL U14370 ( .A(n23400), .B(n23399), .Y(n23500) );
  NAND2XL U14371 ( .A(n23338), .B(n23337), .Y(n23390) );
  INVXL U14372 ( .A(n23392), .Y(n23339) );
  NOR2XL U14373 ( .A(n23297), .B(n23296), .Y(n23388) );
  AOI21XL U14374 ( .A0(n23295), .A1(n23389), .B0(n23394), .Y(n23336) );
  NAND2XL U14375 ( .A(n23297), .B(n23296), .Y(n23391) );
  INVXL U14376 ( .A(n23293), .Y(n23241) );
  NAND2XL U14377 ( .A(n23244), .B(n23243), .Y(n23292) );
  INVXL U14378 ( .A(n23294), .Y(n23245) );
  NAND2XL U14379 ( .A(n23202), .B(n23201), .Y(n23293) );
  INVXL U14380 ( .A(n23398), .Y(n23295) );
  INVXL U14381 ( .A(n23291), .Y(n23242) );
  NAND2XL U14382 ( .A(n23146), .B(n23145), .Y(n23195) );
  INVXL U14383 ( .A(n23197), .Y(n23147) );
  NOR2XL U14384 ( .A(n22428), .B(U0_pipe4[1]), .Y(n23194) );
  INVXL U14385 ( .A(n23199), .Y(n23144) );
  NAND2XL U14386 ( .A(n22428), .B(U0_pipe4[1]), .Y(n23196) );
  NOR2XL U14387 ( .A(n25118), .B(U0_pipe0[1]), .Y(n25861) );
  INVXL U14388 ( .A(n25866), .Y(n25814) );
  NAND2XL U14389 ( .A(n25118), .B(U0_pipe0[1]), .Y(n25863) );
  AOI21XL U14390 ( .A0(n24340), .A1(n24298), .B0(n24339), .Y(n24383) );
  INVXL U14391 ( .A(n24338), .Y(n24339) );
  NOR2XL U14392 ( .A(n24342), .B(n24341), .Y(n24382) );
  NAND2XL U14393 ( .A(n24342), .B(n24341), .Y(n24381) );
  AOI21XL U14394 ( .A0(n24169), .A1(n24112), .B0(n24168), .Y(n24214) );
  INVXL U14395 ( .A(n24167), .Y(n24168) );
  INVXL U14396 ( .A(n23942), .Y(n23991) );
  NAND2XL U14397 ( .A(n23945), .B(n23944), .Y(n23989) );
  NAND2XL U14398 ( .A(n23895), .B(n23894), .Y(n23942) );
  NAND2XL U14399 ( .A(n23509), .B(n23508), .Y(n23551) );
  INVXL U14400 ( .A(n23553), .Y(n23510) );
  NOR2XL U14401 ( .A(n23460), .B(n23459), .Y(n23550) );
  NAND2XL U14402 ( .A(n23460), .B(n23459), .Y(n23552) );
  NAND2XL U14403 ( .A(n23406), .B(n23405), .Y(n23450) );
  INVXL U14404 ( .A(n23452), .Y(n23407) );
  NOR2XL U14405 ( .A(n23349), .B(n23348), .Y(n23448) );
  AOI21XL U14406 ( .A0(n23347), .A1(n23449), .B0(n23454), .Y(n23404) );
  NAND2XL U14407 ( .A(n23349), .B(n23348), .Y(n23451) );
  NAND2XL U14408 ( .A(n23207), .B(n23206), .Y(n23250) );
  INVXL U14409 ( .A(n23252), .Y(n23208) );
  NOR2XL U14410 ( .A(n23155), .B(n23154), .Y(n23249) );
  INVXL U14411 ( .A(n23254), .Y(n23205) );
  NAND2XL U14412 ( .A(n23155), .B(n23154), .Y(n23251) );
  AOI21XL U14413 ( .A0(n22732), .A1(n22731), .B0(n22730), .Y(n23153) );
  OR2XL U14414 ( .A(U0_pipe15[1]), .B(U0_pipe14[1]), .Y(n22732) );
  AND2XL U14415 ( .A(U0_pipe15[1]), .B(U0_pipe14[1]), .Y(n22730) );
  OR2XL U14416 ( .A(n28907), .B(U0_pipe14[0]), .Y(n22731) );
  NOR2XL U14417 ( .A(n22728), .B(n28899), .Y(n23152) );
  NAND2XL U14418 ( .A(n22728), .B(n28899), .Y(n23151) );
  AOI21XL U14419 ( .A0(n26999), .A1(n26957), .B0(n26998), .Y(n27045) );
  INVXL U14420 ( .A(n26997), .Y(n26998) );
  NOR2XL U14421 ( .A(n27001), .B(n27000), .Y(n27044) );
  NAND2XL U14422 ( .A(n27001), .B(n27000), .Y(n27043) );
  INVXL U14423 ( .A(n26827), .Y(n26828) );
  INVXL U14424 ( .A(n26364), .Y(n26417) );
  NAND2XL U14425 ( .A(n26308), .B(n26307), .Y(n26413) );
  INVXL U14426 ( .A(n26411), .Y(n26363) );
  NAND2XL U14427 ( .A(n26177), .B(n26176), .Y(n26216) );
  INVXL U14428 ( .A(n26218), .Y(n26178) );
  NOR2XL U14429 ( .A(n26122), .B(n26121), .Y(n26215) );
  INVXL U14430 ( .A(n26537), .Y(n26306) );
  NAND2XL U14431 ( .A(n26122), .B(n26121), .Y(n26217) );
  NAND2XL U14432 ( .A(n26067), .B(n26066), .Y(n26112) );
  INVXL U14433 ( .A(n26114), .Y(n26068) );
  NOR2XL U14434 ( .A(n26016), .B(n26015), .Y(n26110) );
  NAND2XL U14435 ( .A(n26016), .B(n26015), .Y(n26113) );
  NAND2XL U14436 ( .A(n25874), .B(n25873), .Y(n25915) );
  INVXL U14437 ( .A(n25917), .Y(n25875) );
  NOR2XL U14438 ( .A(n25825), .B(n25824), .Y(n25914) );
  INVXL U14439 ( .A(n25919), .Y(n25872) );
  NAND2XL U14440 ( .A(n25825), .B(n25824), .Y(n25916) );
  AOI21XL U14441 ( .A0(n25454), .A1(n25453), .B0(n25452), .Y(n25823) );
  OR2XL U14442 ( .A(U0_pipe13[1]), .B(U0_pipe12[1]), .Y(n25454) );
  AND2XL U14443 ( .A(U0_pipe13[1]), .B(U0_pipe12[1]), .Y(n25452) );
  OR2XL U14444 ( .A(n28906), .B(U0_pipe12[0]), .Y(n25453) );
  NOR2XL U14445 ( .A(n25450), .B(n28898), .Y(n25822) );
  NAND2XL U14446 ( .A(n25450), .B(n28898), .Y(n25821) );
  INVXL U14447 ( .A(n24362), .Y(n24363) );
  NOR2XL U14448 ( .A(n24366), .B(n24365), .Y(n24389) );
  NAND2XL U14449 ( .A(n24366), .B(n24365), .Y(n24388) );
  AOI21XL U14450 ( .A0(n24177), .A1(n24149), .B0(n24176), .Y(n24222) );
  INVXL U14451 ( .A(n24175), .Y(n24176) );
  NAND2XL U14452 ( .A(n23864), .B(n23863), .Y(n23951) );
  INVXL U14453 ( .A(n23949), .Y(n23899) );
  INVXL U14454 ( .A(n23620), .Y(n23532) );
  NAND2XL U14455 ( .A(n23536), .B(n23535), .Y(n23619) );
  INVXL U14456 ( .A(n23621), .Y(n23537) );
  NAND2XL U14457 ( .A(n23495), .B(n23494), .Y(n23620) );
  INVXL U14458 ( .A(n23618), .Y(n23493) );
  INVXL U14459 ( .A(n23623), .Y(n23492) );
  INVXL U14460 ( .A(n23617), .Y(n23533) );
  NAND2XL U14461 ( .A(n23465), .B(n23464), .Y(n23489) );
  INVXL U14462 ( .A(n23491), .Y(n23466) );
  NOR2XL U14463 ( .A(n23384), .B(n23383), .Y(n23488) );
  INVXL U14464 ( .A(n23862), .Y(n23625) );
  NAND2XL U14465 ( .A(n23384), .B(n23383), .Y(n23490) );
  NAND2XL U14466 ( .A(n23331), .B(n23330), .Y(n23374) );
  INVXL U14467 ( .A(n23376), .Y(n23332) );
  NOR2XL U14468 ( .A(n23287), .B(n23286), .Y(n23372) );
  AOI21XL U14469 ( .A0(n23285), .A1(n23373), .B0(n23378), .Y(n23329) );
  NAND2XL U14470 ( .A(n23287), .B(n23286), .Y(n23375) );
  INVXL U14471 ( .A(n23283), .Y(n23260) );
  NAND2XL U14472 ( .A(n23263), .B(n23262), .Y(n23282) );
  INVXL U14473 ( .A(n23284), .Y(n23264) );
  NAND2XL U14474 ( .A(n23220), .B(n23219), .Y(n23283) );
  INVXL U14475 ( .A(n23382), .Y(n23285) );
  INVXL U14476 ( .A(n23281), .Y(n23261) );
  NAND2XL U14477 ( .A(n23161), .B(n23160), .Y(n23213) );
  INVXL U14478 ( .A(n23215), .Y(n23162) );
  NOR2XL U14479 ( .A(n22104), .B(U0_pipe6[1]), .Y(n23212) );
  INVXL U14480 ( .A(n23217), .Y(n23159) );
  NAND2XL U14481 ( .A(n22104), .B(U0_pipe6[1]), .Y(n23214) );
  AOI21XL U14482 ( .A0(n27007), .A1(n26965), .B0(n27006), .Y(n27052) );
  INVXL U14483 ( .A(n27005), .Y(n27006) );
  NOR2XL U14484 ( .A(n27009), .B(n27008), .Y(n27051) );
  NAND2XL U14485 ( .A(n27009), .B(n27008), .Y(n27050) );
  AOI21XL U14486 ( .A0(n26853), .A1(n26810), .B0(n26852), .Y(n26898) );
  INVXL U14487 ( .A(n26851), .Y(n26852) );
  INVXL U14488 ( .A(n26723), .Y(n26690) );
  INVXL U14489 ( .A(n26720), .Y(n26691) );
  NAND2XL U14490 ( .A(n26693), .B(n26692), .Y(n26721) );
  INVXL U14491 ( .A(n26722), .Y(n26694) );
  INVXL U14492 ( .A(B5_q[0]), .Y(n15985) );
  INVXL U14493 ( .A(B6_q[0]), .Y(n15578) );
  AOI22XL U14494 ( .A0(B6_q[10]), .A1(n15958), .B0(B7_q[10]), .B1(n15982), .Y(
        n15937) );
  AOI22XL U14495 ( .A0(B5_q[10]), .A1(n16344), .B0(B7_q[10]), .B1(n16325), .Y(
        n15731) );
  AOI22XL U14496 ( .A0(B5_q[10]), .A1(n16165), .B0(B7_q[10]), .B1(n16128), .Y(
        n15539) );
  AOI22XL U14497 ( .A0(B5_q[10]), .A1(n16559), .B0(B6_q[10]), .B1(n16570), .Y(
        n15337) );
  AOI22XL U14498 ( .A0(B7_q[11]), .A1(n15982), .B0(B6_q[11]), .B1(n15958), .Y(
        n15933) );
  AOI22XL U14499 ( .A0(B5_q[11]), .A1(n16344), .B0(B6_q[11]), .B1(n16354), .Y(
        n15727) );
  AOI22XL U14500 ( .A0(B4_q[11]), .A1(n7126), .B0(B7_q[11]), .B1(n7127), .Y(
        n15330) );
  AOI22XL U14501 ( .A0(B6_q[12]), .A1(n15958), .B0(B5_q[12]), .B1(n15963), .Y(
        n15929) );
  AOI22XL U14502 ( .A0(B6_q[12]), .A1(n16354), .B0(B5_q[12]), .B1(n16344), .Y(
        n15723) );
  AOI22XL U14503 ( .A0(B7_q[12]), .A1(n16158), .B0(B5_q[12]), .B1(n16165), .Y(
        n15531) );
  AOI22XL U14504 ( .A0(B7_q[12]), .A1(n7127), .B0(B6_q[12]), .B1(n16570), .Y(
        n15322) );
  INVXL U14505 ( .A(B7_q[13]), .Y(n15927) );
  INVXL U14506 ( .A(B4_q[13]), .Y(n15316) );
  AOI22XL U14507 ( .A0(B5_q[14]), .A1(n15963), .B0(B6_q[14]), .B1(n15958), .Y(
        n15921) );
  AOI22XL U14508 ( .A0(B7_q[14]), .A1(n16325), .B0(B6_q[14]), .B1(n5926), .Y(
        n15715) );
  AOI22XL U14509 ( .A0(B5_q[14]), .A1(n16165), .B0(B6_q[14]), .B1(n16143), .Y(
        n15524) );
  AOI22XL U14510 ( .A0(B7_q[14]), .A1(n7127), .B0(B5_q[14]), .B1(n16559), .Y(
        n15306) );
  AOI22XL U14511 ( .A0(B6_q[15]), .A1(n15958), .B0(B7_q[15]), .B1(n5930), .Y(
        n15917) );
  AOI22XL U14512 ( .A0(B6_q[15]), .A1(n16354), .B0(B4_q[15]), .B1(n15687), .Y(
        n15711) );
  AOI22XL U14513 ( .A0(B7_q[15]), .A1(n7127), .B0(B6_q[15]), .B1(n16570), .Y(
        n15299) );
  AOI22XL U14514 ( .A0(B6_q[16]), .A1(n16143), .B0(B5_q[16]), .B1(n16165), .Y(
        n15516) );
  AOI22XL U14515 ( .A0(B7_q[16]), .A1(n7127), .B0(B6_q[16]), .B1(n16570), .Y(
        n15292) );
  AOI22XL U14516 ( .A0(B7_q[17]), .A1(n5930), .B0(B4_q[17]), .B1(n5925), .Y(
        n15909) );
  AOI22XL U14517 ( .A0(B7_q[17]), .A1(n16325), .B0(B4_q[17]), .B1(n15687), .Y(
        n15703) );
  AOI22XL U14518 ( .A0(B6_q[17]), .A1(n16143), .B0(B4_q[17]), .B1(n15557), .Y(
        n15512) );
  AOI22XL U14519 ( .A0(B7_q[17]), .A1(n7127), .B0(B6_q[17]), .B1(n16570), .Y(
        n15284) );
  INVXL U14520 ( .A(B7_q[18]), .Y(n15907) );
  AOI22XL U14521 ( .A0(B6_q[19]), .A1(n15958), .B0(B7_q[19]), .B1(n5930), .Y(
        n15901) );
  AOI22XL U14522 ( .A0(B5_q[19]), .A1(n16165), .B0(B7_q[19]), .B1(n16128), .Y(
        n15505) );
  AOI22XL U14523 ( .A0(B5_q[19]), .A1(n16375), .B0(B6_q[19]), .B1(n16570), .Y(
        n15270) );
  INVXL U14524 ( .A(B7_q[1]), .Y(n15574) );
  INVXL U14525 ( .A(B5_q[20]), .Y(n15899) );
  INVXL U14526 ( .A(B6_q[20]), .Y(n15503) );
  INVXL U14527 ( .A(B4_q[20]), .Y(n15264) );
  AOI22XL U14528 ( .A0(B4_q[21]), .A1(n5925), .B0(B7_q[21]), .B1(n5930), .Y(
        n15893) );
  AOI22XL U14529 ( .A0(B7_q[21]), .A1(n16325), .B0(B6_q[21]), .B1(n16354), .Y(
        n15688) );
  AOI22XL U14530 ( .A0(B5_q[21]), .A1(n16165), .B0(B6_q[21]), .B1(n16143), .Y(
        n15497) );
  AOI22XL U14531 ( .A0(B7_q[21]), .A1(n7127), .B0(B5_q[21]), .B1(n16559), .Y(
        n15254) );
  INVXL U14532 ( .A(B5_q[22]), .Y(n15891) );
  INVXL U14533 ( .A(B6_q[22]), .Y(n15685) );
  INVXL U14534 ( .A(B4_q[22]), .Y(n15248) );
  AOI22XL U14535 ( .A0(B6_q[23]), .A1(n15958), .B0(B5_q[23]), .B1(n15963), .Y(
        n15885) );
  AOI22XL U14536 ( .A0(B7_q[23]), .A1(n16325), .B0(B5_q[23]), .B1(n16344), .Y(
        n15679) );
  AOI22XL U14537 ( .A0(B7_q[23]), .A1(n16128), .B0(B5_q[23]), .B1(n16165), .Y(
        n15489) );
  AOI22XL U14538 ( .A0(B7_q[23]), .A1(n7127), .B0(B6_q[23]), .B1(n16570), .Y(
        n15239) );
  INVXL U14539 ( .A(B7_q[25]), .Y(n15484) );
  INVXL U14540 ( .A(B7_q[26]), .Y(n15480) );
  AOI22XL U14541 ( .A0(B6_q[27]), .A1(n16143), .B0(B7_q[27]), .B1(n16128), .Y(
        n15474) );
  AOI22XL U14542 ( .A0(B5_q[27]), .A1(n16559), .B0(B6_q[27]), .B1(n16570), .Y(
        n14999) );
  INVXL U14543 ( .A(B5_q[28]), .Y(n15867) );
  INVXL U14544 ( .A(B7_q[28]), .Y(n15664) );
  INVXL U14545 ( .A(B4_q[28]), .Y(n15036) );
  AOI22XL U14546 ( .A0(B7_q[29]), .A1(n16128), .B0(B5_q[29]), .B1(n16165), .Y(
        n15467) );
  AOI22XL U14547 ( .A0(B7_q[29]), .A1(n7127), .B0(B6_q[29]), .B1(n16570), .Y(
        n15371) );
  AOI22XL U14548 ( .A0(B7_q[2]), .A1(n15982), .B0(B6_q[2]), .B1(n15958), .Y(
        n15974) );
  AOI22XL U14549 ( .A0(B4_q[2]), .A1(n15687), .B0(B6_q[2]), .B1(n16354), .Y(
        n15763) );
  AOI22XL U14550 ( .A0(B7_q[2]), .A1(n16128), .B0(B4_q[2]), .B1(n15557), .Y(
        n15568) );
  INVXL U14551 ( .A(B6_q[34]), .Y(n15643) );
  INVXL U14552 ( .A(B5_q[34]), .Y(n15843) );
  INVXL U14553 ( .A(B4_q[34]), .Y(n15015) );
  AOI22XL U14554 ( .A0(B4_q[35]), .A1(n5925), .B0(B6_q[35]), .B1(n15958), .Y(
        n15837) );
  AOI22XL U14555 ( .A0(B7_q[35]), .A1(n16128), .B0(B6_q[35]), .B1(n16143), .Y(
        n15448) );
  AOI22XL U14556 ( .A0(B7_q[37]), .A1(n15982), .B0(B4_q[37]), .B1(n5925), .Y(
        n15829) );
  AOI22XL U14557 ( .A0(B6_q[38]), .A1(n15958), .B0(B7_q[38]), .B1(n5930), .Y(
        n15825) );
  AOI22XL U14558 ( .A0(B6_q[38]), .A1(n16143), .B0(B7_q[38]), .B1(n16128), .Y(
        n15436) );
  AOI22XL U14559 ( .A0(B5_q[38]), .A1(n16375), .B0(B6_q[38]), .B1(n16570), .Y(
        n15318) );
  INVXL U14560 ( .A(B5_q[39]), .Y(n15823) );
  INVXL U14561 ( .A(B6_q[39]), .Y(n15434) );
  INVXL U14562 ( .A(B4_q[39]), .Y(n15312) );
  AOI22XL U14563 ( .A0(B4_q[42]), .A1(n5925), .B0(B7_q[42]), .B1(n5930), .Y(
        n15809) );
  AOI22XL U14564 ( .A0(B6_q[42]), .A1(n16293), .B0(B4_q[42]), .B1(n15687), .Y(
        n15612) );
  AOI22XL U14565 ( .A0(B6_q[42]), .A1(n16143), .B0(B7_q[42]), .B1(n16128), .Y(
        n15421) );
  AOI22XL U14566 ( .A0(B7_q[44]), .A1(n15982), .B0(B6_q[44]), .B1(n15958), .Y(
        n15801) );
  AOI22XL U14567 ( .A0(B4_q[44]), .A1(n15557), .B0(B6_q[44]), .B1(n16161), .Y(
        n15414) );
  AOI22XL U14568 ( .A0(B4_q[44]), .A1(n7126), .B0(B7_q[44]), .B1(n7127), .Y(
        n15274) );
  AOI22XL U14569 ( .A0(B6_q[46]), .A1(n15958), .B0(B7_q[46]), .B1(n5930), .Y(
        n15793) );
  AOI22XL U14570 ( .A0(B5_q[46]), .A1(n16344), .B0(B7_q[46]), .B1(n16325), .Y(
        n15597) );
  AOI22XL U14571 ( .A0(B6_q[46]), .A1(n16143), .B0(B7_q[46]), .B1(n16128), .Y(
        n15407) );
  INVXL U14572 ( .A(B5_q[47]), .Y(n15595) );
  INVXL U14573 ( .A(B7_q[47]), .Y(n15791) );
  INVXL U14574 ( .A(B7_q[48]), .Y(n15402) );
  INVXL U14575 ( .A(R7_valid), .Y(n15349) );
  INVXL U14576 ( .A(B7_q[49]), .Y(n15398) );
  INVXL U14577 ( .A(B5_q[4]), .Y(n15758) );
  INVXL U14578 ( .A(B7_q[4]), .Y(n15966) );
  AOI22XL U14579 ( .A0(B6_q[50]), .A1(n15958), .B0(B4_q[50]), .B1(n15969), .Y(
        n15777) );
  AOI22XL U14580 ( .A0(B7_q[50]), .A1(n16325), .B0(B4_q[50]), .B1(n15687), .Y(
        n15583) );
  AOI22XL U14581 ( .A0(B7_q[50]), .A1(n16128), .B0(B4_q[50]), .B1(n15557), .Y(
        n15392) );
  NOR2XL U14582 ( .A(n7305), .B(A_sel_reg[4]), .Y(n14995) );
  AOI22XL U14583 ( .A0(B7_q[50]), .A1(n7127), .B0(B6_q[50]), .B1(n16570), .Y(
        n15229) );
  INVXL U14584 ( .A(R7_valid), .Y(n16501) );
  INVXL U14585 ( .A(R7_valid), .Y(n16461) );
  AOI22XL U14586 ( .A0(B7_q[5]), .A1(n15982), .B0(B4_q[5]), .B1(n15969), .Y(
        n15959) );
  AOI22XL U14587 ( .A0(B6_q[5]), .A1(n16143), .B0(B4_q[5]), .B1(n15557), .Y(
        n15558) );
  AOI22XL U14588 ( .A0(B7_q[6]), .A1(n15982), .B0(B4_q[6]), .B1(n15969), .Y(
        n15954) );
  AOI22XL U14589 ( .A0(B7_q[6]), .A1(n16325), .B0(B4_q[6]), .B1(n15687), .Y(
        n15748) );
  AOI22XL U14590 ( .A0(B6_q[6]), .A1(n16143), .B0(B4_q[6]), .B1(n15557), .Y(
        n15553) );
  INVXL U14591 ( .A(R7_valid), .Y(n16470) );
  INVXL U14592 ( .A(B5_q[7]), .Y(n15745) );
  INVXL U14593 ( .A(B7_q[7]), .Y(n15952) );
  INVXL U14594 ( .A(B5_q[8]), .Y(n15741) );
  CLKINVX3 U14595 ( .A(n15431), .Y(n15495) );
  INVXL U14596 ( .A(B6_q[8]), .Y(n15947) );
  INVXL U14597 ( .A(B4_q[8]), .Y(n15347) );
  AOI22XL U14598 ( .A0(B6_q[9]), .A1(n15958), .B0(B4_q[9]), .B1(n5925), .Y(
        n15941) );
  AOI22XL U14599 ( .A0(B7_q[9]), .A1(n16325), .B0(B4_q[9]), .B1(n15687), .Y(
        n15735) );
  AOI22XL U14600 ( .A0(B6_q[9]), .A1(n16161), .B0(B4_q[9]), .B1(n5933), .Y(
        n15543) );
  AOI22XL U14601 ( .A0(B7_q[9]), .A1(n7127), .B0(B6_q[9]), .B1(n16570), .Y(
        n15341) );
  NAND2XL U14602 ( .A(n21332), .B(n21331), .Y(n21381) );
  NOR2XL U14603 ( .A(n21380), .B(n21382), .Y(n21441) );
  NAND2XL U14604 ( .A(n21387), .B(n21386), .Y(n21442) );
  NOR2XL U14605 ( .A(n21672), .B(n21671), .Y(n21710) );
  NAND2XL U14606 ( .A(n21672), .B(n21671), .Y(n21709) );
  AOI21XL U14607 ( .A0(n21670), .A1(n21633), .B0(n21669), .Y(n21711) );
  INVXL U14608 ( .A(n21668), .Y(n21669) );
  NAND2XL U14609 ( .A(n16936), .B(U1_pipe6[1]), .Y(n17799) );
  NOR2XL U14610 ( .A(n16936), .B(U1_pipe6[1]), .Y(n17797) );
  NAND2XL U14611 ( .A(n17760), .B(n17759), .Y(n17798) );
  INVXL U14612 ( .A(n17800), .Y(n17761) );
  INVXL U14613 ( .A(n17802), .Y(n17758) );
  NOR2XL U14614 ( .A(n17929), .B(n17928), .Y(n17985) );
  NAND2XL U14615 ( .A(n17929), .B(n17928), .Y(n17988) );
  NAND2XL U14616 ( .A(n17947), .B(n17946), .Y(n17987) );
  INVXL U14617 ( .A(n17989), .Y(n17948) );
  AOI21XL U14618 ( .A0(n17927), .A1(n17986), .B0(n17991), .Y(n17945) );
  NAND2XL U14619 ( .A(n17997), .B(n17996), .Y(n18102) );
  NOR2XL U14620 ( .A(n17997), .B(n17996), .Y(n18100) );
  NAND2XL U14621 ( .A(n18087), .B(n18086), .Y(n18101) );
  INVXL U14622 ( .A(n18103), .Y(n18088) );
  INVXL U14623 ( .A(n18438), .Y(n18239) );
  NAND2XL U14624 ( .A(n18241), .B(n18240), .Y(n18321) );
  INVXL U14625 ( .A(n18274), .Y(n18325) );
  INVXL U14626 ( .A(n18319), .Y(n18273) );
  INVXL U14627 ( .A(n18321), .Y(n18272) );
  NAND2XL U14628 ( .A(n18276), .B(n18275), .Y(n18320) );
  INVXL U14629 ( .A(n18322), .Y(n18277) );
  NAND2XL U14630 ( .A(n18620), .B(n18619), .Y(n18690) );
  NOR2XL U14631 ( .A(n18689), .B(n18691), .Y(n18753) );
  NAND2XL U14632 ( .A(n18696), .B(n18695), .Y(n18754) );
  AOI21XL U14633 ( .A0(n18897), .A1(n18851), .B0(n18896), .Y(n18937) );
  INVXL U14634 ( .A(n18895), .Y(n18896) );
  NOR2XL U14635 ( .A(n18899), .B(n18898), .Y(n18936) );
  NAND2XL U14636 ( .A(n18899), .B(n18898), .Y(n18935) );
  NOR2XL U14637 ( .A(n18975), .B(n18974), .Y(n18996) );
  NAND2XL U14638 ( .A(n18975), .B(n18974), .Y(n18995) );
  AOI21XL U14639 ( .A0(n18973), .A1(n18938), .B0(n18972), .Y(n18997) );
  INVXL U14640 ( .A(n18971), .Y(n18972) );
  NAND2XL U14641 ( .A(n20493), .B(n20492), .Y(n20581) );
  NOR2XL U14642 ( .A(n20493), .B(n20492), .Y(n20579) );
  NAND2XL U14643 ( .A(n20535), .B(n20534), .Y(n20580) );
  INVXL U14644 ( .A(n20582), .Y(n20536) );
  INVXL U14645 ( .A(n20584), .Y(n20533) );
  NOR2XL U14646 ( .A(n20680), .B(n20679), .Y(n20780) );
  NAND2XL U14647 ( .A(n20680), .B(n20679), .Y(n20783) );
  NAND2XL U14648 ( .A(n20728), .B(n20727), .Y(n20782) );
  INVXL U14649 ( .A(n20784), .Y(n20729) );
  AOI21XL U14650 ( .A0(n20678), .A1(n20781), .B0(n20786), .Y(n20726) );
  NAND2XL U14651 ( .A(n20792), .B(n20791), .Y(n20881) );
  NOR2XL U14652 ( .A(n20792), .B(n20791), .Y(n20879) );
  NAND2XL U14653 ( .A(n20837), .B(n20836), .Y(n20880) );
  INVXL U14654 ( .A(n20882), .Y(n20838) );
  INVXL U14655 ( .A(n21210), .Y(n20973) );
  NAND2XL U14656 ( .A(n20975), .B(n20974), .Y(n21078) );
  INVXL U14657 ( .A(n21027), .Y(n21082) );
  INVXL U14658 ( .A(n21076), .Y(n21026) );
  NAND2XL U14659 ( .A(n21029), .B(n21028), .Y(n21077) );
  NAND2XL U14660 ( .A(n21321), .B(n21320), .Y(n21370) );
  NOR2XL U14661 ( .A(n21369), .B(n21371), .Y(n21429) );
  NAND2XL U14662 ( .A(n21376), .B(n21375), .Y(n21430) );
  AOI21XL U14663 ( .A0(n21488), .A1(n21436), .B0(n21487), .Y(n21538) );
  INVXL U14664 ( .A(n21486), .Y(n21487) );
  NAND2XL U14665 ( .A(n21541), .B(n21540), .Y(n21580) );
  NOR2XL U14666 ( .A(n21664), .B(n21663), .Y(n21703) );
  NAND2XL U14667 ( .A(n21664), .B(n21663), .Y(n21702) );
  AOI21XL U14668 ( .A0(n21662), .A1(n21625), .B0(n21661), .Y(n21704) );
  INVXL U14669 ( .A(n21660), .Y(n21661) );
  AOI21XL U14670 ( .A0(n17451), .A1(n17450), .B0(n17449), .Y(n17774) );
  OR2XL U14671 ( .A(U1_pipe15[1]), .B(U1_pipe14[1]), .Y(n17451) );
  AND2XL U14672 ( .A(U1_pipe15[1]), .B(U1_pipe14[1]), .Y(n17449) );
  OR2XL U14673 ( .A(n28911), .B(U1_pipe14[0]), .Y(n17450) );
  NOR2XL U14674 ( .A(n17447), .B(n28903), .Y(n17773) );
  NAND2XL U14675 ( .A(n17447), .B(n28903), .Y(n17772) );
  NAND2XL U14676 ( .A(n17776), .B(n17775), .Y(n17868) );
  NOR2XL U14677 ( .A(n17776), .B(n17775), .Y(n17866) );
  NAND2XL U14678 ( .A(n17821), .B(n17820), .Y(n17867) );
  INVXL U14679 ( .A(n17869), .Y(n17822) );
  INVXL U14680 ( .A(n17871), .Y(n17819) );
  NOR2XL U14681 ( .A(n17965), .B(n17964), .Y(n18070) );
  NAND2XL U14682 ( .A(n17965), .B(n17964), .Y(n18073) );
  NAND2XL U14683 ( .A(n18019), .B(n18018), .Y(n18072) );
  INVXL U14684 ( .A(n18074), .Y(n18020) );
  AOI21XL U14685 ( .A0(n17963), .A1(n18071), .B0(n18076), .Y(n18017) );
  NAND2XL U14686 ( .A(n18082), .B(n18081), .Y(n18168) );
  NOR2XL U14687 ( .A(n18082), .B(n18081), .Y(n18166) );
  NAND2XL U14688 ( .A(n18121), .B(n18120), .Y(n18167) );
  INVXL U14689 ( .A(n18169), .Y(n18122) );
  NAND2XL U14690 ( .A(n18269), .B(n18268), .Y(n18368) );
  INVXL U14691 ( .A(n18312), .Y(n18372) );
  NAND2XL U14692 ( .A(n18314), .B(n18313), .Y(n18367) );
  NAND2XL U14693 ( .A(n18517), .B(n18516), .Y(n18554) );
  NAND2XL U14694 ( .A(n18608), .B(n18607), .Y(n18657) );
  NOR2XL U14695 ( .A(n18656), .B(n18658), .Y(n18716) );
  NAND2XL U14696 ( .A(n18663), .B(n18662), .Y(n18717) );
  NOR2XL U14697 ( .A(n18951), .B(n18950), .Y(n18989) );
  NAND2XL U14698 ( .A(n18951), .B(n18950), .Y(n18988) );
  AOI21XL U14699 ( .A0(n18949), .A1(n18914), .B0(n18948), .Y(n18990) );
  INVXL U14700 ( .A(n18947), .Y(n18948) );
  NAND2XL U14701 ( .A(n17170), .B(U1_pipe4[1]), .Y(n17810) );
  NOR2XL U14702 ( .A(n17170), .B(U1_pipe4[1]), .Y(n17808) );
  NAND2XL U14703 ( .A(n17767), .B(n17766), .Y(n17809) );
  INVXL U14704 ( .A(n17811), .Y(n17768) );
  INVXL U14705 ( .A(n17813), .Y(n17765) );
  NAND2XL U14706 ( .A(n17816), .B(n17815), .Y(n17907) );
  INVXL U14707 ( .A(n17905), .Y(n17859) );
  INVXL U14708 ( .A(n17907), .Y(n17858) );
  NAND2XL U14709 ( .A(n17861), .B(n17860), .Y(n17906) );
  INVXL U14710 ( .A(n17908), .Y(n17862) );
  INVXL U14711 ( .A(n18011), .Y(n17909) );
  NOR2XL U14712 ( .A(n17911), .B(n17910), .Y(n18001) );
  NAND2XL U14713 ( .A(n17911), .B(n17910), .Y(n18004) );
  NAND2XL U14714 ( .A(n17954), .B(n17953), .Y(n18003) );
  INVXL U14715 ( .A(n18005), .Y(n17955) );
  AOI21XL U14716 ( .A0(n17909), .A1(n18002), .B0(n18007), .Y(n17952) );
  NAND2XL U14717 ( .A(n18013), .B(n18012), .Y(n18112) );
  NOR2XL U14718 ( .A(n18013), .B(n18012), .Y(n18110) );
  NAND2XL U14719 ( .A(n18065), .B(n18064), .Y(n18111) );
  INVXL U14720 ( .A(n18113), .Y(n18066) );
  INVXL U14721 ( .A(n18457), .Y(n18217) );
  NAND2XL U14722 ( .A(n18338), .B(n18337), .Y(n18447) );
  INVXL U14723 ( .A(n18443), .Y(n18387) );
  INVXL U14724 ( .A(n18447), .Y(n18386) );
  NAND2XL U14725 ( .A(n18390), .B(n18389), .Y(n18446) );
  INVXL U14726 ( .A(n18448), .Y(n18391) );
  INVXL U14727 ( .A(n18444), .Y(n18335) );
  INVXL U14728 ( .A(n18450), .Y(n18334) );
  NAND2XL U14729 ( .A(n18632), .B(n18631), .Y(n18679) );
  NOR2XL U14730 ( .A(n18678), .B(n18680), .Y(n18741) );
  NAND2XL U14731 ( .A(n18685), .B(n18684), .Y(n18742) );
  NOR2XL U14732 ( .A(n18967), .B(n18966), .Y(n19003) );
  NAND2XL U14733 ( .A(n18967), .B(n18966), .Y(n19002) );
  AOI21XL U14734 ( .A0(n18965), .A1(n18930), .B0(n18964), .Y(n19004) );
  INVXL U14735 ( .A(n18963), .Y(n18964) );
  NAND2XL U14736 ( .A(n20501), .B(n20500), .Y(n20562) );
  NOR2XL U14737 ( .A(n20501), .B(n20500), .Y(n20560) );
  NAND2XL U14738 ( .A(n20542), .B(n20541), .Y(n20561) );
  INVXL U14739 ( .A(n20563), .Y(n20543) );
  INVXL U14740 ( .A(n20565), .Y(n20540) );
  NOR2XL U14741 ( .A(n20690), .B(n20689), .Y(n20758) );
  NAND2XL U14742 ( .A(n20690), .B(n20689), .Y(n20761) );
  NAND2XL U14743 ( .A(n20705), .B(n20704), .Y(n20760) );
  INVXL U14744 ( .A(n20762), .Y(n20706) );
  AOI21XL U14745 ( .A0(n20688), .A1(n20759), .B0(n20764), .Y(n20703) );
  NAND2XL U14746 ( .A(n20770), .B(n20769), .Y(n20891) );
  NOR2XL U14747 ( .A(n20770), .B(n20769), .Y(n20889) );
  NAND2XL U14748 ( .A(n20843), .B(n20842), .Y(n20890) );
  INVXL U14749 ( .A(n20892), .Y(n20844) );
  INVXL U14750 ( .A(n21258), .Y(n20986) );
  NAND2XL U14751 ( .A(n20988), .B(n20987), .Y(n21089) );
  INVXL U14752 ( .A(n21036), .Y(n21093) );
  NAND2XL U14753 ( .A(n21038), .B(n21037), .Y(n21088) );
  NAND2XL U14754 ( .A(n21355), .B(n21354), .Y(n21403) );
  NOR2XL U14755 ( .A(n21402), .B(n21404), .Y(n21465) );
  NAND2XL U14756 ( .A(n21409), .B(n21408), .Y(n21466) );
  NOR2XL U14757 ( .A(n21592), .B(n21591), .Y(n21647) );
  NAND2XL U14758 ( .A(n21592), .B(n21591), .Y(n21646) );
  NOR2XL U14759 ( .A(n21688), .B(n21687), .Y(n21724) );
  NAND2XL U14760 ( .A(n21688), .B(n21687), .Y(n21723) );
  INVXL U14761 ( .A(n21684), .Y(n21685) );
  NAND2XL U14762 ( .A(n17746), .B(U1_pipe10[1]), .Y(n17828) );
  NOR2XL U14763 ( .A(n17746), .B(U1_pipe10[1]), .Y(n17826) );
  NAND2XL U14764 ( .A(n17782), .B(n17781), .Y(n17827) );
  INVXL U14765 ( .A(n17829), .Y(n17783) );
  INVXL U14766 ( .A(n17831), .Y(n17780) );
  NOR2XL U14767 ( .A(n17901), .B(n17900), .Y(n18024) );
  NAND2XL U14768 ( .A(n17901), .B(n17900), .Y(n18027) );
  NAND2XL U14769 ( .A(n17971), .B(n17970), .Y(n18026) );
  INVXL U14770 ( .A(n18028), .Y(n17972) );
  AOI21XL U14771 ( .A0(n17899), .A1(n18025), .B0(n18030), .Y(n17969) );
  INVXL U14772 ( .A(n18129), .Y(n18060) );
  NAND2XL U14773 ( .A(n18133), .B(n18132), .Y(n18199) );
  INVXL U14774 ( .A(n18196), .Y(n18177) );
  INVXL U14775 ( .A(n18197), .Y(n18131) );
  INVXL U14776 ( .A(n18202), .Y(n18130) );
  NAND2XL U14777 ( .A(n18206), .B(n18205), .Y(n18343) );
  INVXL U14778 ( .A(n18292), .Y(n18347) );
  NAND2XL U14779 ( .A(n18294), .B(n18293), .Y(n18342) );
  NAND2XL U14780 ( .A(n18728), .B(n18672), .Y(n18733) );
  AOI21XL U14781 ( .A0(n18731), .A1(n18672), .B0(n18730), .Y(n18732) );
  INVXL U14782 ( .A(n18729), .Y(n18730) );
  AOI21XL U14783 ( .A0(n18800), .A1(n18735), .B0(n18799), .Y(n18834) );
  INVXL U14784 ( .A(n18798), .Y(n18799) );
  NOR2XL U14785 ( .A(n18802), .B(n18801), .Y(n18833) );
  NAND2XL U14786 ( .A(n18802), .B(n18801), .Y(n18832) );
  NOR2XL U14787 ( .A(n18959), .B(n18958), .Y(n19010) );
  NAND2XL U14788 ( .A(n18959), .B(n18958), .Y(n19009) );
  AOI21XL U14789 ( .A0(n18957), .A1(n18922), .B0(n18956), .Y(n19011) );
  INVXL U14790 ( .A(n18955), .Y(n18956) );
  NAND2XL U14791 ( .A(n20478), .B(n20477), .Y(n20592) );
  NOR2XL U14792 ( .A(n20478), .B(n20477), .Y(n20590) );
  NAND2XL U14793 ( .A(n20517), .B(n20516), .Y(n20591) );
  INVXL U14794 ( .A(n20593), .Y(n20518) );
  INVXL U14795 ( .A(n20595), .Y(n20515) );
  NOR2XL U14796 ( .A(n20663), .B(n20662), .Y(n20796) );
  NAND2XL U14797 ( .A(n20663), .B(n20662), .Y(n20799) );
  NAND2XL U14798 ( .A(n20735), .B(n20734), .Y(n20798) );
  INVXL U14799 ( .A(n20800), .Y(n20736) );
  AOI21XL U14800 ( .A0(n20661), .A1(n20797), .B0(n20802), .Y(n20733) );
  NAND2XL U14801 ( .A(n20808), .B(n20807), .Y(n20862) );
  NOR2XL U14802 ( .A(n20808), .B(n20807), .Y(n20860) );
  NAND2XL U14803 ( .A(n20821), .B(n20820), .Y(n20861) );
  INVXL U14804 ( .A(n20863), .Y(n20822) );
  INVXL U14805 ( .A(n21230), .Y(n21008) );
  NAND2XL U14806 ( .A(n19705), .B(U1_pipe0[1]), .Y(n20524) );
  NOR2XL U14807 ( .A(n19705), .B(U1_pipe0[1]), .Y(n20522) );
  NAND2XL U14808 ( .A(n20484), .B(n20483), .Y(n20523) );
  INVXL U14809 ( .A(n20525), .Y(n20485) );
  INVXL U14810 ( .A(n20527), .Y(n20482) );
  NOR2XL U14811 ( .A(n20625), .B(n20624), .Y(n20710) );
  NAND2XL U14812 ( .A(n20625), .B(n20624), .Y(n20713) );
  NAND2XL U14813 ( .A(n20669), .B(n20668), .Y(n20712) );
  INVXL U14814 ( .A(n20714), .Y(n20670) );
  NAND2XL U14815 ( .A(n20722), .B(n20721), .Y(n20828) );
  NOR2XL U14816 ( .A(n20722), .B(n20721), .Y(n20826) );
  NAND2XL U14817 ( .A(n20775), .B(n20774), .Y(n20827) );
  INVXL U14818 ( .A(n20829), .Y(n20776) );
  INVXL U14819 ( .A(n21161), .Y(n20927) );
  NAND2XL U14820 ( .A(n20929), .B(n20928), .Y(n21045) );
  INVXL U14821 ( .A(n20993), .Y(n21049) );
  INVXL U14822 ( .A(n21043), .Y(n20992) );
  NAND2XL U14823 ( .A(n20995), .B(n20994), .Y(n21044) );
  NAND2XL U14824 ( .A(n21344), .B(n21343), .Y(n21392) );
  NOR2XL U14825 ( .A(n21391), .B(n21393), .Y(n21453) );
  NAND2XL U14826 ( .A(n21398), .B(n21397), .Y(n21454) );
  NOR2XL U14827 ( .A(n21680), .B(n21679), .Y(n21717) );
  NAND2XL U14828 ( .A(n21680), .B(n21679), .Y(n21716) );
  AOI21XL U14829 ( .A0(n21678), .A1(n21641), .B0(n21677), .Y(n21718) );
  INVXL U14830 ( .A(n21676), .Y(n21677) );
  NOR2X1 U14831 ( .A(n26038), .B(n26037), .Y(n26142) );
  AOI21XL U14832 ( .A0(n26034), .A1(n26143), .B0(n26148), .Y(n26079) );
  INVXL U14833 ( .A(n26347), .Y(n26240) );
  INVXL U14834 ( .A(n26817), .Y(n26763) );
  NOR2XL U14835 ( .A(U2_A_i_d[0]), .B(n21730), .Y(n23131) );
  NAND2XL U14836 ( .A(U2_A_i_d[0]), .B(n21730), .Y(n23167) );
  NAND2XL U14837 ( .A(n23179), .B(n23178), .Y(n23270) );
  NOR2XL U14838 ( .A(n23179), .B(n23178), .Y(n23268) );
  INVXL U14839 ( .A(n23271), .Y(n23228) );
  INVXL U14840 ( .A(n23573), .Y(n23528) );
  INVXL U14841 ( .A(n23685), .Y(n23637) );
  INVXL U14842 ( .A(n23682), .Y(n23575) );
  NAND2X1 U14843 ( .A(n23744), .B(n23745), .Y(n23789) );
  INVXL U14844 ( .A(n23927), .Y(n23874) );
  INVXL U14845 ( .A(n24036), .Y(n23980) );
  INVXL U14846 ( .A(n24039), .Y(n23985) );
  INVXL U14847 ( .A(n24157), .Y(n24095) );
  INVX1 U14848 ( .A(n24205), .Y(n24158) );
  INVXL U14849 ( .A(n24200), .Y(n24201) );
  NAND2XL U14850 ( .A(n20510), .B(n20509), .Y(n20548) );
  INVXL U14851 ( .A(n20550), .Y(n20511) );
  NAND2XL U14852 ( .A(n20470), .B(U2_A_r_d[1]), .Y(n20549) );
  INVXL U14853 ( .A(n20553), .Y(n20505) );
  INVXL U14854 ( .A(n20750), .Y(n20649) );
  INVXL U14855 ( .A(n20950), .Y(n20900) );
  OAI21XL U14856 ( .A0(n20958), .A1(n20853), .B0(n20852), .Y(n20901) );
  INVXL U14857 ( .A(n20951), .Y(n20853) );
  INVXL U14858 ( .A(n21063), .Y(n21014) );
  INVXL U14859 ( .A(n21066), .Y(n21020) );
  INVXL U14860 ( .A(n21175), .Y(n21119) );
  INVXL U14861 ( .A(n21179), .Y(n21118) );
  INVXL U14862 ( .A(n21176), .Y(n21068) );
  INVXL U14863 ( .A(n21182), .Y(n21067) );
  INVXL U14864 ( .A(n21304), .Y(n21265) );
  INVXL U14865 ( .A(n21307), .Y(n21269) );
  INVXL U14866 ( .A(n21417), .Y(n21365) );
  INVX1 U14867 ( .A(n21481), .Y(n7404) );
  INVX1 U14868 ( .A(n21482), .Y(n7405) );
  INVXL U14869 ( .A(n21527), .Y(n21421) );
  INVXL U14870 ( .A(n21612), .Y(n21613) );
  INVXL U14871 ( .A(n26991), .Y(n21655) );
  INVXL U14872 ( .A(n26990), .Y(n21654) );
  INVXL U14873 ( .A(n21692), .Y(n7414) );
  INVXL U14874 ( .A(n27033), .Y(n21697) );
  INVXL U14875 ( .A(n27032), .Y(n21696) );
  NOR2XL U14876 ( .A(n16604), .B(n16619), .Y(n16622) );
  NAND2XL U14877 ( .A(n17792), .B(n17791), .Y(n17838) );
  INVXL U14878 ( .A(n17840), .Y(n17793) );
  NAND2XL U14879 ( .A(n17754), .B(U2_A_i_d[1]), .Y(n17839) );
  INVXL U14880 ( .A(n17843), .Y(n17787) );
  AOI21XL U14881 ( .A0(n17937), .A1(n18041), .B0(n18046), .Y(n17976) );
  INVXL U14882 ( .A(n18139), .Y(n18096) );
  INVXL U14883 ( .A(n18248), .Y(n18192) );
  INVXL U14884 ( .A(n18250), .Y(n18140) );
  INVXL U14885 ( .A(n18591), .Y(n18545) );
  INVXL U14886 ( .A(n18704), .Y(n18654) );
  INVXL U14887 ( .A(n18807), .Y(n18709) );
  INVXL U14888 ( .A(n24373), .Y(n18984) );
  INVXL U14889 ( .A(n24372), .Y(n18983) );
  NAND2XL U14890 ( .A(n25850), .B(n25849), .Y(n25938) );
  NAND2XL U14891 ( .A(n25890), .B(n25889), .Y(n25937) );
  INVXL U14892 ( .A(n25939), .Y(n25891) );
  INVXL U14893 ( .A(n25942), .Y(n25886) );
  INVXL U14894 ( .A(n26152), .Y(n26034) );
  NOR2XL U14895 ( .A(n19045), .B(n19060), .Y(n19063) );
  NOR2XL U14896 ( .A(U2_A_r_d[0]), .B(n24409), .Y(n25799) );
  NAND2XL U14897 ( .A(U2_A_r_d[0]), .B(n24409), .Y(n25838) );
  INVXL U14898 ( .A(n24714), .Y(n24716) );
  NAND2XL U14899 ( .A(n24721), .B(n24720), .Y(n24998) );
  NOR2X1 U14900 ( .A(n24641), .B(n24664), .Y(n25011) );
  NAND2XL U14901 ( .A(n24745), .B(n24744), .Y(n25020) );
  INVXL U14902 ( .A(n25007), .Y(n7561) );
  INVXL U14903 ( .A(n24802), .Y(n25062) );
  INVXL U14904 ( .A(n25093), .Y(n25104) );
  NAND2XL U14905 ( .A(n24851), .B(n25448), .Y(n25111) );
  NAND2XL U14906 ( .A(n22454), .B(U2_A_r_d[25]), .Y(n24865) );
  NOR2X1 U14907 ( .A(n24875), .B(n24434), .Y(n7272) );
  NAND2X1 U14908 ( .A(n14146), .B(n7075), .Y(n24445) );
  INVXL U14909 ( .A(n24899), .Y(n24902) );
  NAND2XL U14910 ( .A(n14025), .B(U2_A_r_d[7]), .Y(n24946) );
  INVXL U14911 ( .A(n24964), .Y(n24975) );
  INVXL U14912 ( .A(n22050), .Y(n22376) );
  INVXL U14913 ( .A(n22406), .Y(n22416) );
  INVXL U14914 ( .A(n22218), .Y(n22221) );
  INVXL U14915 ( .A(n22219), .Y(n22220) );
  INVXL U14916 ( .A(n22238), .Y(n22262) );
  INVXL U14917 ( .A(n22264), .Y(n22277) );
  INVXL U14918 ( .A(n22279), .Y(n22286) );
  AND2XL U14919 ( .A(n25458), .B(U2_A_i_d[0]), .Y(n22291) );
  INVXL U14920 ( .A(n24752), .Y(n24755) );
  INVXL U14921 ( .A(n24753), .Y(n24754) );
  INVXL U14922 ( .A(n24771), .Y(n24766) );
  NAND2XL U14923 ( .A(n24781), .B(n24780), .Y(n25052) );
  NAND2XL U14924 ( .A(n24798), .B(n24797), .Y(n25063) );
  INVXL U14925 ( .A(n24796), .Y(n24798) );
  INVXL U14926 ( .A(n24825), .Y(n24818) );
  INVXL U14927 ( .A(n24819), .Y(n24821) );
  INVXL U14928 ( .A(n24810), .Y(n24828) );
  INVXL U14929 ( .A(n24817), .Y(n24826) );
  INVXL U14930 ( .A(n24833), .Y(n24835) );
  INVXL U14931 ( .A(n24830), .Y(n24841) );
  AND2XL U14932 ( .A(n24591), .B(n24590), .Y(n24592) );
  NAND2XL U14933 ( .A(n8850), .B(n24843), .Y(n25108) );
  NAND2XL U14934 ( .A(n24847), .B(n25106), .Y(n25112) );
  INVXL U14935 ( .A(n24424), .Y(n24426) );
  INVXL U14936 ( .A(n24430), .Y(n24433) );
  NAND2XL U14937 ( .A(n24469), .B(n24468), .Y(n24893) );
  NAND2XL U14938 ( .A(n24473), .B(n24890), .Y(n24896) );
  NAND2XL U14939 ( .A(n24484), .B(n24483), .Y(n24905) );
  NAND2XL U14940 ( .A(n24495), .B(n24494), .Y(n24913) );
  NAND2X1 U14941 ( .A(n24503), .B(n7588), .Y(n7587) );
  NOR2XL U14942 ( .A(n24505), .B(n7603), .Y(n7588) );
  NAND2XL U14943 ( .A(n24509), .B(n24508), .Y(n24923) );
  NAND2XL U14944 ( .A(n24525), .B(n24524), .Y(n24934) );
  NOR2XL U14945 ( .A(n24547), .B(n24545), .Y(n24539) );
  OAI21XL U14946 ( .A0(n24553), .A1(n24547), .B0(n24548), .Y(n24538) );
  NAND2XL U14947 ( .A(n14067), .B(U2_A_r_d[7]), .Y(n24540) );
  NAND2XL U14948 ( .A(n14066), .B(U2_A_r_d[6]), .Y(n24548) );
  INVXL U14949 ( .A(n24537), .Y(n24556) );
  INVXL U14950 ( .A(n24545), .Y(n24554) );
  INVXL U14951 ( .A(n24559), .Y(n24561) );
  INVXL U14952 ( .A(n24558), .Y(n24569) );
  INVXL U14953 ( .A(n24578), .Y(n13351) );
  NAND2XL U14954 ( .A(n14061), .B(U2_A_r_d[2]), .Y(n24572) );
  NAND2XL U14955 ( .A(n14020), .B(U2_A_r_d[2]), .Y(n24978) );
  INVXL U14956 ( .A(n25574), .Y(n25577) );
  INVXL U14957 ( .A(n25594), .Y(n25617) );
  INVXL U14958 ( .A(n25457), .Y(n25627) );
  INVXL U14959 ( .A(n25634), .Y(n25641) );
  AND2XL U14960 ( .A(n25458), .B(U2_A_r_d[0]), .Y(n25646) );
  XOR2XL U14961 ( .A(n12359), .B(n12358), .Y(n12360) );
  INVXL U14962 ( .A(n21957), .Y(n21960) );
  INVXL U14963 ( .A(n22044), .Y(n22046) );
  NAND2XL U14964 ( .A(n14527), .B(n22887), .Y(n22061) );
  INVXL U14965 ( .A(n22065), .Y(n22074) );
  NOR2XL U14966 ( .A(n14521), .B(n22890), .Y(n22080) );
  INVXL U14967 ( .A(n22078), .Y(n22089) );
  INVXL U14968 ( .A(n22098), .Y(n14517) );
  AND2XL U14969 ( .A(n14515), .B(n22892), .Y(n14516) );
  NAND2XL U14970 ( .A(n22093), .B(n22092), .Y(n22419) );
  INVXL U14971 ( .A(n22091), .Y(n22093) );
  NAND2XL U14972 ( .A(n5768), .B(n22097), .Y(n22422) );
  NAND2XL U14973 ( .A(n21818), .B(n22174), .Y(n22183) );
  INVXL U14974 ( .A(n22175), .Y(n21818) );
  INVXL U14975 ( .A(n21822), .Y(n21825) );
  NAND2XL U14976 ( .A(n21826), .B(n22170), .Y(n22188) );
  NAND2XL U14977 ( .A(n22168), .B(n22166), .Y(n22193) );
  NAND2XL U14978 ( .A(n22155), .B(n22152), .Y(n22213) );
  NAND2XL U14979 ( .A(n22149), .B(n22146), .Y(n22224) );
  INVXL U14980 ( .A(n21860), .Y(n21863) );
  INVXL U14981 ( .A(n21861), .Y(n21862) );
  NAND2XL U14982 ( .A(n22140), .B(n22222), .Y(n22227) );
  NAND2XL U14983 ( .A(n8057), .B(n22144), .Y(n22232) );
  NAND2XL U14984 ( .A(n22116), .B(n22114), .Y(n22243) );
  NOR2XL U14985 ( .A(n21750), .B(n21916), .Y(n21912) );
  NAND2XL U14986 ( .A(n22134), .B(n22132), .Y(n22267) );
  INVXL U14987 ( .A(n21910), .Y(n21925) );
  NAND2XL U14988 ( .A(n21930), .B(n22126), .Y(n22282) );
  INVXL U14989 ( .A(n22127), .Y(n21930) );
  INVXL U14990 ( .A(n21927), .Y(n21936) );
  NAND2XL U14991 ( .A(n21934), .B(n22280), .Y(n22285) );
  INVXL U14992 ( .A(n22281), .Y(n21934) );
  NAND2XL U14993 ( .A(n21938), .B(n22124), .Y(n22289) );
  INVXL U14994 ( .A(n22125), .Y(n21938) );
  NAND2XL U14995 ( .A(n21942), .B(n22122), .Y(n22292) );
  NAND2XL U14996 ( .A(n21963), .B(n21962), .Y(n22306) );
  NAND2XL U14997 ( .A(n21974), .B(n22309), .Y(n22314) );
  INVXL U14998 ( .A(n22320), .Y(n22321) );
  NAND2XL U14999 ( .A(n21992), .B(n21991), .Y(n22332) );
  INVXL U15000 ( .A(n22338), .Y(n22339) );
  NAND2XL U15001 ( .A(n22030), .B(n22029), .Y(n22366) );
  AND2XL U15002 ( .A(n14016), .B(U2_A_r_d[0]), .Y(n24983) );
  NAND2XL U15003 ( .A(n5778), .B(n24577), .Y(n24984) );
  AND2XL U15004 ( .A(n14386), .B(U2_A_r_d[11]), .Y(n25210) );
  NAND2XL U15005 ( .A(n6980), .B(n25481), .Y(n25598) );
  NOR2XL U15006 ( .A(n14344), .B(n25247), .Y(n25241) );
  NAND2XL U15007 ( .A(n25242), .B(n25469), .Y(n25622) );
  INVXL U15008 ( .A(n25239), .Y(n25258) );
  NAND2XL U15009 ( .A(n25627), .B(n25625), .Y(n25631) );
  NAND2XL U15010 ( .A(n25264), .B(n25463), .Y(n25637) );
  INVXL U15011 ( .A(n25260), .Y(n25272) );
  NAND2XL U15012 ( .A(n25276), .B(n25461), .Y(n25644) );
  INVXL U15013 ( .A(n25462), .Y(n25276) );
  NAND2XL U15014 ( .A(n25280), .B(n25459), .Y(n25647) );
  NAND2XL U15015 ( .A(n5858), .B(n24684), .Y(n22985) );
  INVXL U15016 ( .A(n23026), .Y(n23029) );
  NAND2BX1 U15017 ( .AN(n7410), .B(n22935), .Y(n23043) );
  INVXL U15018 ( .A(n23104), .Y(n23113) );
  AND2XL U15019 ( .A(n22894), .B(n24590), .Y(n8002) );
  INVXL U15020 ( .A(n22751), .Y(n22754) );
  NAND2XL U15021 ( .A(n14146), .B(U2_A_i_d[21]), .Y(n22759) );
  INVXL U15022 ( .A(n22783), .Y(n22786) );
  NAND2XL U15023 ( .A(n14067), .B(U2_A_i_d[7]), .Y(n22841) );
  NAND2XL U15024 ( .A(n14066), .B(U2_A_i_d[6]), .Y(n22849) );
  NAND2XL U15025 ( .A(n14065), .B(U2_A_i_d[5]), .Y(n22855) );
  INVXL U15026 ( .A(n22838), .Y(n22858) );
  INVXL U15027 ( .A(n22861), .Y(n22863) );
  INVXL U15028 ( .A(n22860), .Y(n22871) );
  INVXL U15029 ( .A(n22880), .Y(n14060) );
  NAND2XL U15030 ( .A(n14061), .B(U2_A_i_d[2]), .Y(n22874) );
  INVXL U15031 ( .A(n25292), .Y(n25294) );
  INVXL U15032 ( .A(n25302), .Y(n25304) );
  NOR2X1 U15033 ( .A(n14550), .B(n24641), .Y(n25684) );
  AOI2BB1X2 U15034 ( .A0N(n25693), .A1N(n25680), .B0(n25682), .Y(n25689) );
  INVXL U15035 ( .A(n25700), .Y(n25701) );
  NAND2XL U15036 ( .A(n24615), .B(n13114), .Y(n25742) );
  INVXL U15037 ( .A(n25741), .Y(n25743) );
  INVXL U15038 ( .A(n25775), .Y(n25782) );
  AND2XL U15039 ( .A(n25448), .B(n13098), .Y(n25788) );
  NOR2XL U15040 ( .A(n7410), .B(n22935), .Y(n12606) );
  INVX1 U15041 ( .A(n22657), .Y(n22685) );
  NAND2XL U15042 ( .A(n24600), .B(n22890), .Y(n22714) );
  NAND2XL U15043 ( .A(n22710), .B(n22709), .Y(n23107) );
  INVXL U15044 ( .A(n22708), .Y(n22710) );
  NAND2XL U15045 ( .A(n22715), .B(n22714), .Y(n23111) );
  INVXL U15046 ( .A(n22713), .Y(n22715) );
  INVXL U15047 ( .A(n22707), .Y(n22716) );
  NOR2XL U15048 ( .A(n24590), .B(n22892), .Y(n22718) );
  NAND2XL U15049 ( .A(n24590), .B(n22892), .Y(n22723) );
  NAND2XL U15050 ( .A(n22720), .B(n22719), .Y(n23115) );
  NAND2XL U15051 ( .A(n24851), .B(n22727), .Y(n22725) );
  NAND2XL U15052 ( .A(n22724), .B(n22723), .Y(n23119) );
  NAND2XL U15053 ( .A(n22454), .B(U2_A_i_d[25]), .Y(n22463) );
  NAND2BX1 U15054 ( .AN(n22474), .B(n7612), .Y(n7611) );
  INVXL U15055 ( .A(n22468), .Y(n22470) );
  NAND2XL U15056 ( .A(n22494), .B(n22493), .Y(n22775) );
  NAND2XL U15057 ( .A(n22506), .B(n22505), .Y(n22789) );
  INVXL U15058 ( .A(n22500), .Y(n22503) );
  INVXL U15059 ( .A(n22501), .Y(n22502) );
  NAND2XL U15060 ( .A(n22515), .B(n22514), .Y(n22799) );
  NAND2XL U15061 ( .A(n22526), .B(n22525), .Y(n22812) );
  NAND2XL U15062 ( .A(n22537), .B(n22536), .Y(n22826) );
  INVXL U15063 ( .A(n22535), .Y(n22537) );
  INVXL U15064 ( .A(n22521), .Y(n22547) );
  NOR2XL U15065 ( .A(n22558), .B(n22556), .Y(n22551) );
  INVXL U15066 ( .A(n22549), .Y(n22567) );
  INVXL U15067 ( .A(n22570), .Y(n22572) );
  INVXL U15068 ( .A(n22569), .Y(n22580) );
  NAND2XL U15069 ( .A(n14021), .B(U2_A_i_d[3]), .Y(n22577) );
  NAND2XL U15070 ( .A(n14020), .B(U2_A_i_d[2]), .Y(n22583) );
  AND2XL U15071 ( .A(n14016), .B(U2_A_i_d[0]), .Y(n22589) );
  NAND2XL U15072 ( .A(n14017), .B(n22588), .Y(n22879) );
  INVXL U15073 ( .A(n25395), .Y(n25388) );
  NAND2XL U15074 ( .A(n14536), .B(n24615), .Y(n25390) );
  INVXL U15075 ( .A(n25387), .Y(n25396) );
  INVXL U15076 ( .A(n25419), .Y(n25412) );
  INVXL U15077 ( .A(n25413), .Y(n25415) );
  INVXL U15078 ( .A(n25404), .Y(n25422) );
  INVXL U15079 ( .A(n25411), .Y(n25420) );
  NAND2XL U15080 ( .A(n25429), .B(n25428), .Y(n25778) );
  INVXL U15081 ( .A(n25424), .Y(n25435) );
  INVXL U15082 ( .A(n25445), .Y(n12364) );
  NAND2XL U15083 ( .A(n25439), .B(n25438), .Y(n25785) );
  INVXL U15084 ( .A(n25437), .Y(n25439) );
  NOR2XL U15085 ( .A(n25449), .B(n25448), .Y(n25445) );
  INVXL U15086 ( .A(n25137), .Y(n25139) );
  NAND2XL U15087 ( .A(n25141), .B(n25518), .Y(n25539) );
  NAND2XL U15088 ( .A(n25513), .B(n25542), .Y(n25547) );
  AND2XL U15089 ( .A(n14453), .B(U2_A_r_d[19]), .Y(n25160) );
  OAI21XL U15090 ( .A0(n25170), .A1(n25159), .B0(n25158), .Y(n25168) );
  INVXL U15091 ( .A(n25182), .Y(n25185) );
  INVXL U15092 ( .A(n25183), .Y(n25184) );
  NAND2XL U15093 ( .A(n25493), .B(n25491), .Y(n25588) );
  INVXL U15094 ( .A(n19847), .Y(n19850) );
  NAND2X1 U15095 ( .A(n19824), .B(n7529), .Y(n7528) );
  AND2X1 U15096 ( .A(n19775), .B(U1_A_r_d0[23]), .Y(n19780) );
  INVXL U15097 ( .A(n20176), .Y(n19955) );
  AND2XL U15098 ( .A(n14908), .B(n19954), .Y(n8010) );
  INVXL U15099 ( .A(n20156), .Y(n20167) );
  NAND2XL U15100 ( .A(n19966), .B(n19965), .Y(n20151) );
  NAND2XL U15101 ( .A(n19970), .B(n19969), .Y(n20139) );
  INVXL U15102 ( .A(n20079), .Y(n20082) );
  AND2XL U15103 ( .A(n13665), .B(U1_A_i_d0[0]), .Y(n17294) );
  NOR2XL U15104 ( .A(n13670), .B(U1_A_i_d0[3]), .Y(n17283) );
  INVXL U15105 ( .A(n17277), .Y(n17286) );
  INVXL U15106 ( .A(n17243), .Y(n17252) );
  OAI21XL U15107 ( .A0(n17257), .A1(n17242), .B0(n17255), .Y(n17253) );
  INVXL U15108 ( .A(n17239), .Y(n17235) );
  OAI21X2 U15109 ( .A0(n13719), .A1(n7701), .B0(n7700), .Y(n17209) );
  INVX1 U15110 ( .A(n13721), .Y(n7701) );
  NAND2XL U15111 ( .A(n19507), .B(n16932), .Y(n17443) );
  INVXL U15112 ( .A(n17424), .Y(n17426) );
  INVXL U15113 ( .A(n17423), .Y(n17434) );
  NAND2X1 U15114 ( .A(n5869), .B(n7520), .Y(n17364) );
  NAND2BX1 U15115 ( .AN(n19544), .B(n5862), .Y(n17359) );
  INVX1 U15116 ( .A(n17322), .Y(n7782) );
  NAND2X1 U15117 ( .A(n5868), .B(n5865), .Y(n17345) );
  INVXL U15118 ( .A(n17306), .Y(n7552) );
  NOR2X1 U15119 ( .A(n13560), .B(n7501), .Y(n13561) );
  NAND2BX1 U15120 ( .AN(n17325), .B(n7554), .Y(n7553) );
  NAND2BX1 U15121 ( .AN(n7861), .B(n7863), .Y(n14108) );
  NOR2X1 U15122 ( .A(n19568), .B(n7863), .Y(n14107) );
  NAND2XL U15123 ( .A(n14866), .B(n20175), .Y(n20456) );
  NAND2XL U15124 ( .A(n20171), .B(n20170), .Y(n20453) );
  OAI21XL U15125 ( .A0(n20428), .A1(n20434), .B0(n20429), .Y(n20420) );
  NOR2X1 U15126 ( .A(n14945), .B(n20005), .Y(n20367) );
  NAND2X1 U15127 ( .A(n7843), .B(n19999), .Y(n20355) );
  NAND2X1 U15128 ( .A(n20386), .B(n20310), .Y(n7445) );
  NAND2XL U15129 ( .A(n20072), .B(n20071), .Y(n20357) );
  NAND2XL U15130 ( .A(n20324), .B(n20322), .Y(n20346) );
  INVXL U15131 ( .A(n20327), .Y(n20042) );
  INVXL U15132 ( .A(n20337), .Y(n20335) );
  NAND2XL U15133 ( .A(n9570), .B(n17293), .Y(n17591) );
  INVXL U15134 ( .A(n17592), .Y(n9400) );
  NAND2XL U15135 ( .A(n17290), .B(n17289), .Y(n17587) );
  INVXL U15136 ( .A(n17288), .Y(n17290) );
  NAND2XL U15137 ( .A(n9658), .B(U1_A_i_d0[3]), .Y(n17577) );
  NAND2XL U15138 ( .A(n17280), .B(n17279), .Y(n17579) );
  INVXL U15139 ( .A(n17576), .Y(n17585) );
  INVXL U15140 ( .A(n17564), .Y(n17567) );
  INVXL U15141 ( .A(n17565), .Y(n17566) );
  NAND2XL U15142 ( .A(n17270), .B(n17269), .Y(n17568) );
  NAND2XL U15143 ( .A(n9665), .B(U1_A_i_d0[6]), .Y(n9415) );
  NAND2XL U15144 ( .A(n17263), .B(n17262), .Y(n17560) );
  INVXL U15145 ( .A(n17557), .Y(n17574) );
  INVXL U15146 ( .A(n17245), .Y(n17247) );
  NAND2XL U15147 ( .A(n6996), .B(n17225), .Y(n17518) );
  NAND2XL U15148 ( .A(n17217), .B(n17216), .Y(n17508) );
  INVXL U15149 ( .A(n17502), .Y(n17505) );
  AND2X2 U15150 ( .A(U1_A_i_d0[19]), .B(n9512), .Y(n17481) );
  NAND2XL U15151 ( .A(n13728), .B(n13727), .Y(n17483) );
  INVXL U15152 ( .A(n17739), .Y(n12863) );
  INVXL U15153 ( .A(n17719), .Y(n17730) );
  INVXL U15154 ( .A(n17610), .Y(n17611) );
  NAND2X1 U15155 ( .A(n17609), .B(n7969), .Y(n17604) );
  AND2XL U15156 ( .A(n19711), .B(U1_A_r_d0[1]), .Y(n19712) );
  INVXL U15157 ( .A(n19947), .Y(n19713) );
  NAND2XL U15158 ( .A(n19717), .B(U1_A_r_d0[3]), .Y(n19928) );
  NOR2XL U15159 ( .A(n19717), .B(U1_A_r_d0[3]), .Y(n19929) );
  INVXL U15160 ( .A(n19927), .Y(n19938) );
  INVXL U15161 ( .A(n19906), .Y(n19925) );
  AND2XL U15162 ( .A(n13665), .B(U1_A_r_d0[0]), .Y(n19501) );
  INVXL U15163 ( .A(n17103), .Y(n17097) );
  INVXL U15164 ( .A(n17084), .Y(n17085) );
  INVXL U15165 ( .A(n17083), .Y(n17086) );
  INVX1 U15166 ( .A(n14006), .Y(n7821) );
  NAND2X1 U15167 ( .A(n14962), .B(n20050), .Y(n17063) );
  NAND2X1 U15168 ( .A(n14968), .B(n20032), .Y(n16790) );
  NAND2BX1 U15169 ( .AN(n13988), .B(n7508), .Y(n7507) );
  NAND2BXL U15170 ( .AN(n16789), .B(n13987), .Y(n7510) );
  AND2XL U15171 ( .A(n19711), .B(U1_A_i_d0[1]), .Y(n8642) );
  NAND2XL U15172 ( .A(n19717), .B(U1_A_i_d0[3]), .Y(n16758) );
  NOR2XL U15173 ( .A(n19717), .B(U1_A_i_d0[3]), .Y(n16759) );
  INVXL U15174 ( .A(n16757), .Y(n16768) );
  INVXL U15175 ( .A(n16702), .Y(n16734) );
  INVXL U15176 ( .A(n16678), .Y(n16681) );
  INVXL U15177 ( .A(n16679), .Y(n16680) );
  NAND2XL U15178 ( .A(n16645), .B(n16644), .Y(n16947) );
  INVXL U15179 ( .A(n16929), .Y(n14910) );
  AND2XL U15180 ( .A(n14908), .B(n14907), .Y(n14909) );
  INVXL U15181 ( .A(n16909), .Y(n16920) );
  OAI21XL U15182 ( .A0(n16898), .A1(n16904), .B0(n16899), .Y(n16890) );
  NAND2XL U15183 ( .A(n13881), .B(n16865), .Y(n17114) );
  NAND2XL U15184 ( .A(n7018), .B(n16861), .Y(n17111) );
  INVXL U15185 ( .A(n16834), .Y(n16835) );
  AND2X2 U15186 ( .A(n14956), .B(n14955), .Y(n16824) );
  INVX1 U15187 ( .A(n16788), .Y(n7838) );
  NAND2XL U15188 ( .A(n12287), .B(n19946), .Y(n20305) );
  NAND2XL U15189 ( .A(n19942), .B(n19941), .Y(n20302) );
  INVXL U15190 ( .A(n19940), .Y(n19942) );
  NAND2XL U15191 ( .A(n19932), .B(n19931), .Y(n20295) );
  INVXL U15192 ( .A(n19930), .Y(n19932) );
  INVXL U15193 ( .A(n20292), .Y(n20299) );
  NAND2XL U15194 ( .A(n12286), .B(n19909), .Y(n20280) );
  INVXL U15195 ( .A(n20253), .Y(n20275) );
  NAND2XL U15196 ( .A(n19878), .B(n19877), .Y(n20257) );
  NAND2XL U15197 ( .A(n12310), .B(n19864), .Y(n20247) );
  NAND2XL U15198 ( .A(n19854), .B(n19853), .Y(n20238) );
  INVXL U15199 ( .A(n20232), .Y(n20235) );
  NAND2XL U15200 ( .A(n19756), .B(U1_A_r_d0[17]), .Y(n20223) );
  NAND2XL U15201 ( .A(n19839), .B(n19838), .Y(n20226) );
  INVXL U15202 ( .A(n20212), .Y(n20213) );
  INVXL U15203 ( .A(n20211), .Y(n20214) );
  NAND2XL U15204 ( .A(n19814), .B(n19813), .Y(n20202) );
  NAND2XL U15205 ( .A(n19807), .B(n19806), .Y(n20197) );
  NAND2X1 U15206 ( .A(n12330), .B(n19797), .Y(n7303) );
  NAND2XL U15207 ( .A(n13666), .B(n19227), .Y(n19502) );
  INVXL U15208 ( .A(n19228), .Y(n9654) );
  NAND2XL U15209 ( .A(n19223), .B(n19222), .Y(n19499) );
  INVXL U15210 ( .A(n19221), .Y(n19223) );
  NAND2XL U15211 ( .A(n9658), .B(U1_A_r_d0[3]), .Y(n19208) );
  INVXL U15212 ( .A(n19207), .Y(n19219) );
  NAND2XL U15213 ( .A(n9665), .B(U1_A_r_d0[6]), .Y(n9666) );
  INVXL U15214 ( .A(n19186), .Y(n19205) );
  AND2XL U15215 ( .A(n9680), .B(U1_A_r_d0[11]), .Y(n19155) );
  INVXL U15216 ( .A(n19374), .Y(n14737) );
  AND2XL U15217 ( .A(n14734), .B(n19373), .Y(n14735) );
  INVXL U15218 ( .A(n19355), .Y(n19366) );
  NAND2XL U15219 ( .A(n7357), .B(n19519), .Y(n19345) );
  NOR2XL U15220 ( .A(n19344), .B(n19342), .Y(n19336) );
  OR2X2 U15221 ( .A(n14755), .B(n19520), .Y(n19338) );
  NAND2XL U15222 ( .A(n14755), .B(n19520), .Y(n19337) );
  INVXL U15223 ( .A(n19334), .Y(n19353) );
  INVX1 U15224 ( .A(n19301), .Y(n19332) );
  NAND2XL U15225 ( .A(n19542), .B(n14826), .Y(n19292) );
  INVXL U15226 ( .A(n19276), .Y(n19279) );
  NAND2XL U15227 ( .A(n7861), .B(n20333), .Y(n7855) );
  NAND2XL U15228 ( .A(n8510), .B(n16776), .Y(n17047) );
  NAND2XL U15229 ( .A(n16772), .B(n16771), .Y(n17044) );
  INVXL U15230 ( .A(n16770), .Y(n16772) );
  NAND2XL U15231 ( .A(n16762), .B(n16761), .Y(n17037) );
  INVXL U15232 ( .A(n16760), .Y(n16762) );
  INVXL U15233 ( .A(n17034), .Y(n17041) );
  NOR2X1 U15234 ( .A(n6583), .B(n16753), .Y(n17020) );
  NAND2XL U15235 ( .A(n16740), .B(n16739), .Y(n17021) );
  NAND2XL U15236 ( .A(n8553), .B(n16712), .Y(n17001) );
  NAND2XL U15237 ( .A(n16708), .B(n16707), .Y(n16998) );
  NAND2XL U15238 ( .A(n8174), .B(n16670), .Y(n16970) );
  NAND2XL U15239 ( .A(n8148), .B(n16648), .Y(n16952) );
  AOI21XL U15240 ( .A0(n16957), .A1(n8616), .B0(n8615), .Y(n8617) );
  NAND2XL U15241 ( .A(n13833), .B(n16928), .Y(n17164) );
  NAND2XL U15242 ( .A(n16924), .B(n16923), .Y(n17161) );
  INVXL U15243 ( .A(n16922), .Y(n16924) );
  NAND2XL U15244 ( .A(n16914), .B(n16913), .Y(n17154) );
  INVXL U15245 ( .A(n16912), .Y(n16914) );
  INVXL U15246 ( .A(n17151), .Y(n17158) );
  INVXL U15247 ( .A(n17131), .Y(n17149) );
  INVXL U15248 ( .A(n17107), .Y(n17129) );
  NAND2XL U15249 ( .A(n16877), .B(n16876), .Y(n17122) );
  INVXL U15250 ( .A(n16881), .Y(n17121) );
  NAND2XL U15251 ( .A(n19482), .B(n19480), .Y(n19486) );
  INVXL U15252 ( .A(n19203), .Y(n19482) );
  NAND2XL U15253 ( .A(n13664), .B(n19189), .Y(n19477) );
  INVXL U15254 ( .A(n19178), .Y(n19464) );
  NAND2XL U15255 ( .A(n19134), .B(n19133), .Y(n19437) );
  INVXL U15256 ( .A(n7688), .Y(n19133) );
  NAND2XL U15257 ( .A(n19119), .B(n19118), .Y(n19425) );
  NOR2X1 U15258 ( .A(n13702), .B(U1_A_r_d0[19]), .Y(n19415) );
  AOI21X1 U15259 ( .A0(n19429), .A1(n19413), .B0(n19412), .Y(n19420) );
  NAND2XL U15260 ( .A(n19506), .B(n19693), .Y(n19699) );
  NAND2XL U15261 ( .A(n19507), .B(n20179), .Y(n19698) );
  NAND2XL U15262 ( .A(n19511), .B(n19508), .Y(n19695) );
  NAND2XL U15263 ( .A(n19359), .B(n19514), .Y(n19687) );
  INVXL U15264 ( .A(n19664), .Y(n19682) );
  INVXL U15265 ( .A(n19531), .Y(n19642) );
  INVX1 U15266 ( .A(n19539), .Y(n19631) );
  NAND2XL U15267 ( .A(n19548), .B(n19545), .Y(n19621) );
  NAND2XL U15268 ( .A(n19538), .B(n19609), .Y(n19614) );
  NAND2X1 U15269 ( .A(n7843), .B(n19272), .Y(n19609) );
  NAND2BX1 U15270 ( .AN(n19553), .B(n14835), .Y(n19605) );
  INVXL U15271 ( .A(n19562), .Y(n19244) );
  NAND2XL U15272 ( .A(n13670), .B(U1_A_r_d0[3]), .Y(n19490) );
  NOR2XL U15273 ( .A(n13670), .B(U1_A_r_d0[3]), .Y(n19491) );
  NAND2XL U15274 ( .A(n19212), .B(n19211), .Y(n19492) );
  INVXL U15275 ( .A(n19489), .Y(n19496) );
  NAND2XL U15276 ( .A(n11974), .B(cnt[0]), .Y(n28629) );
  NAND3XL U15277 ( .A(n11974), .B(cnt[1]), .C(cnt[0]), .Y(n28633) );
  NAND3BXL U15278 ( .AN(n11949), .B(cnt[8]), .C(n27814), .Y(n11638) );
  NOR2XL U15279 ( .A(cs[0]), .B(n5808), .Y(n11948) );
  NOR2XL U15280 ( .A(cs[2]), .B(n11633), .Y(n11951) );
  AOI31XL U15281 ( .A0(n11974), .A1(n11973), .A2(n11972), .B0(n28631), .Y(
        n11980) );
  INVXL U15282 ( .A(n14978), .Y(n11647) );
  NOR2BXL U15283 ( .AN(n11613), .B(n28706), .Y(n11648) );
  AOI22XL U15284 ( .A0(n5840), .A1(CQ1[9]), .B0(Q5[9]), .B1(n27211), .Y(n27552) );
  INVXL U15285 ( .A(n27115), .Y(n27555) );
  OAI22XL U15286 ( .A0(n27814), .A1(Q4[9]), .B0(CQ1[9]), .B1(n27976), .Y(
        n27115) );
  AOI22XL U15287 ( .A0(n5840), .A1(CQ1[8]), .B0(Q5[8]), .B1(n27211), .Y(n27546) );
  INVXL U15288 ( .A(n27112), .Y(n27549) );
  OAI22XL U15289 ( .A0(n27814), .A1(Q4[8]), .B0(CQ1[8]), .B1(n27976), .Y(
        n27112) );
  INVXL U15290 ( .A(n27109), .Y(n27543) );
  OAI22XL U15291 ( .A0(n27814), .A1(Q4[7]), .B0(CQ1[7]), .B1(n27976), .Y(
        n27109) );
  AOI22XL U15292 ( .A0(n5840), .A1(CQ1[6]), .B0(Q5[6]), .B1(n27213), .Y(n27534) );
  INVXL U15293 ( .A(n27106), .Y(n27537) );
  OAI22XL U15294 ( .A0(n27814), .A1(Q4[6]), .B0(CQ1[6]), .B1(n27976), .Y(
        n27106) );
  INVXL U15295 ( .A(n27103), .Y(n27531) );
  OAI22XL U15296 ( .A0(n27814), .A1(Q4[5]), .B0(CQ1[5]), .B1(n27976), .Y(
        n27103) );
  OAI21XL U15297 ( .A0(Q6[53]), .A1(OP_done1), .B0(n27278), .Y(n27813) );
  NAND2XL U15298 ( .A(Q4[53]), .B(n27976), .Y(n27277) );
  OAI21XL U15299 ( .A0(Q6[52]), .A1(OP_done1), .B0(n27274), .Y(n27807) );
  NAND2XL U15300 ( .A(Q4[52]), .B(n27976), .Y(n27273) );
  OAI21XL U15301 ( .A0(Q5[52]), .A1(OP_done1), .B0(n27274), .Y(n27802) );
  AOI22XL U15302 ( .A0(n7123), .A1(CQ1[4]), .B0(Q6[4]), .B1(n28922), .Y(n27522) );
  INVXL U15303 ( .A(n27100), .Y(n27525) );
  OAI22XL U15304 ( .A0(n27814), .A1(Q4[4]), .B0(CQ1[4]), .B1(n27976), .Y(
        n27100) );
  OAI21XL U15305 ( .A0(Q5[51]), .A1(OP_done1), .B0(n27270), .Y(n27796) );
  NAND2XL U15306 ( .A(Q4[51]), .B(n27976), .Y(n27269) );
  OAI21XL U15307 ( .A0(Q5[50]), .A1(OP_done1), .B0(n27266), .Y(n27795) );
  NAND2XL U15308 ( .A(Q4[50]), .B(OP2_done0), .Y(n27265) );
  OAI21XL U15309 ( .A0(Q5[49]), .A1(n5840), .B0(n27261), .Y(n27784) );
  NAND2XL U15310 ( .A(Q4[49]), .B(OP2_done0), .Y(n27260) );
  NAND2XL U15311 ( .A(Q4[48]), .B(OP2_done0), .Y(n27256) );
  OAI21XL U15312 ( .A0(Q6[48]), .A1(n5927), .B0(n27257), .Y(n27778) );
  OAI21XL U15313 ( .A0(Q6[47]), .A1(n5927), .B0(n27253), .Y(n27777) );
  NAND2XL U15314 ( .A(Q4[47]), .B(n27976), .Y(n27252) );
  OAI21XL U15315 ( .A0(Q6[46]), .A1(n5840), .B0(n27249), .Y(n27765) );
  NAND2XL U15316 ( .A(Q4[46]), .B(OP2_done0), .Y(n27248) );
  OAI21XL U15317 ( .A0(Q6[45]), .A1(n7123), .B0(n27245), .Y(n27759) );
  NAND2XL U15318 ( .A(Q4[45]), .B(n27976), .Y(n27244) );
  OAI21XL U15319 ( .A0(Q5[44]), .A1(OP_done1), .B0(n27241), .Y(n27758) );
  NAND2XL U15320 ( .A(Q4[44]), .B(n27976), .Y(n27240) );
  OAI21XL U15321 ( .A0(Q6[44]), .A1(n5840), .B0(n27241), .Y(n27753) );
  OAI21XL U15322 ( .A0(Q6[43]), .A1(n7123), .B0(n27237), .Y(n27747) );
  NAND2XL U15323 ( .A(Q4[43]), .B(n27976), .Y(n27235) );
  OAI21XL U15324 ( .A0(Q5[42]), .A1(OP_done1), .B0(n27232), .Y(n27746) );
  NAND2XL U15325 ( .A(Q4[42]), .B(n27976), .Y(n27231) );
  AOI22XL U15326 ( .A0(n7123), .A1(CQ1[3]), .B0(Q6[3]), .B1(n28922), .Y(n27516) );
  INVXL U15327 ( .A(n27097), .Y(n27519) );
  OAI22XL U15328 ( .A0(n28921), .A1(Q4[3]), .B0(CQ1[3]), .B1(n27976), .Y(
        n27097) );
  OAI21XL U15329 ( .A0(Q5[41]), .A1(n5927), .B0(n27228), .Y(n27735) );
  NAND2XL U15330 ( .A(Q4[41]), .B(n27976), .Y(n27227) );
  OAI21XL U15331 ( .A0(Q6[40]), .A1(n5927), .B0(n27224), .Y(n27729) );
  NAND2XL U15332 ( .A(Q4[40]), .B(n27976), .Y(n27223) );
  NAND2XL U15333 ( .A(Q4[39]), .B(n27976), .Y(n27219) );
  OAI21XL U15334 ( .A0(Q6[39]), .A1(n5927), .B0(n27220), .Y(n27723) );
  AOI22XL U15335 ( .A0(n5840), .A1(CQ1[36]), .B0(Q5[38]), .B1(n28922), .Y(
        n27717) );
  INVXL U15336 ( .A(n27216), .Y(n27720) );
  OAI22XL U15337 ( .A0(n27814), .A1(Q4[38]), .B0(CQ1[36]), .B1(n27976), .Y(
        n27216) );
  INVXL U15338 ( .A(n27212), .Y(n27714) );
  OAI22XL U15339 ( .A0(n28921), .A1(Q4[37]), .B0(CQ1[35]), .B1(OP2_done0), .Y(
        n27212) );
  INVXL U15340 ( .A(n27208), .Y(n27708) );
  OAI22XL U15341 ( .A0(n27814), .A1(Q4[36]), .B0(CQ1[34]), .B1(n27976), .Y(
        n27208) );
  AOI22XL U15342 ( .A0(n5840), .A1(CQ1[33]), .B0(Q6[35]), .B1(n28922), .Y(
        n27704) );
  INVXL U15343 ( .A(n27204), .Y(n27702) );
  OAI22XL U15344 ( .A0(n27814), .A1(Q4[35]), .B0(CQ1[33]), .B1(OP2_done0), .Y(
        n27204) );
  AOI22XL U15345 ( .A0(n5840), .A1(CQ1[32]), .B0(Q6[34]), .B1(n27213), .Y(
        n27693) );
  INVXL U15346 ( .A(n27201), .Y(n27696) );
  OAI22XL U15347 ( .A0(n27814), .A1(Q4[34]), .B0(CQ1[32]), .B1(n27976), .Y(
        n27201) );
  INVXL U15348 ( .A(n27198), .Y(n27690) );
  OAI22XL U15349 ( .A0(n27814), .A1(Q4[33]), .B0(CQ1[31]), .B1(n27976), .Y(
        n27198) );
  AOI22XL U15350 ( .A0(n5840), .A1(CQ1[30]), .B0(Q5[32]), .B1(n27211), .Y(
        n27680) );
  INVXL U15351 ( .A(n27195), .Y(n27683) );
  OAI22XL U15352 ( .A0(n27814), .A1(Q4[32]), .B0(CQ1[30]), .B1(n27976), .Y(
        n27195) );
  INVXL U15353 ( .A(n27094), .Y(n27513) );
  OAI22XL U15354 ( .A0(n27814), .A1(Q4[2]), .B0(CQ1[2]), .B1(n27976), .Y(
        n27094) );
  INVXL U15355 ( .A(n27192), .Y(n27677) );
  OAI22XL U15356 ( .A0(n28921), .A1(Q4[31]), .B0(CQ1[29]), .B1(n27976), .Y(
        n27192) );
  INVXL U15357 ( .A(n27189), .Y(n27671) );
  OAI22XL U15358 ( .A0(n27814), .A1(Q4[30]), .B0(CQ1[28]), .B1(n27976), .Y(
        n27189) );
  AOI22XL U15359 ( .A0(n5840), .A1(CQ1[27]), .B0(Q6[29]), .B1(n28922), .Y(
        n27662) );
  INVXL U15360 ( .A(n27186), .Y(n27665) );
  OAI22XL U15361 ( .A0(n27814), .A1(Q4[29]), .B0(CQ1[27]), .B1(OP2_done0), .Y(
        n27186) );
  AOI22XL U15362 ( .A0(n5840), .A1(CQ1[26]), .B0(Q5[28]), .B1(n28922), .Y(
        n27656) );
  INVXL U15363 ( .A(n27183), .Y(n27659) );
  OAI22XL U15364 ( .A0(n27814), .A1(Q4[28]), .B0(CQ1[26]), .B1(n27976), .Y(
        n27183) );
  OAI21XL U15365 ( .A0(Q6[25]), .A1(n5840), .B0(n27180), .Y(n27650) );
  NAND2XL U15366 ( .A(Q4[25]), .B(n27976), .Y(n27179) );
  OAI21XL U15367 ( .A0(Q5[24]), .A1(n5927), .B0(n27176), .Y(n27644) );
  NAND2XL U15368 ( .A(Q4[24]), .B(n27976), .Y(n27175) );
  OAI21XL U15369 ( .A0(Q5[23]), .A1(n5840), .B0(n27172), .Y(n27643) );
  NAND2XL U15370 ( .A(Q4[23]), .B(n27976), .Y(n27171) );
  NAND2XL U15371 ( .A(Q4[22]), .B(n27976), .Y(n27167) );
  OAI21XL U15372 ( .A0(Q6[22]), .A1(OP_done1), .B0(n27168), .Y(n27637) );
  NAND2XL U15373 ( .A(Q4[21]), .B(n27976), .Y(n27163) );
  OAI21XL U15374 ( .A0(Q6[20]), .A1(OP_done1), .B0(n27159), .Y(n27619) );
  NAND2XL U15375 ( .A(Q4[20]), .B(n27976), .Y(n27158) );
  INVXL U15376 ( .A(n27091), .Y(n27507) );
  OAI22XL U15377 ( .A0(n27814), .A1(Q4[1]), .B0(CQ1[1]), .B1(n27976), .Y(
        n27091) );
  OAI21XL U15378 ( .A0(Q5[19]), .A1(OP_done1), .B0(n27155), .Y(n27613) );
  NAND2XL U15379 ( .A(Q4[19]), .B(n27976), .Y(n27154) );
  OAI21XL U15380 ( .A0(Q6[18]), .A1(OP_done1), .B0(n27151), .Y(n27607) );
  NAND2XL U15381 ( .A(Q4[18]), .B(n27976), .Y(n27150) );
  OAI21XL U15382 ( .A0(Q5[17]), .A1(n5840), .B0(n27147), .Y(n27601) );
  NAND2XL U15383 ( .A(Q4[17]), .B(n27976), .Y(n27146) );
  NAND2XL U15384 ( .A(Q4[16]), .B(n27976), .Y(n27142) );
  OAI21XL U15385 ( .A0(Q6[16]), .A1(n5840), .B0(n27143), .Y(n27595) );
  OAI21XL U15386 ( .A0(Q6[15]), .A1(n5840), .B0(n27139), .Y(n27589) );
  NAND2XL U15387 ( .A(Q4[15]), .B(n27976), .Y(n27138) );
  OAI21XL U15388 ( .A0(Q5[14]), .A1(n5840), .B0(n27135), .Y(n27583) );
  OAI21XL U15389 ( .A0(n28958), .A1(n27976), .B0(n27134), .Y(n27586) );
  NAND2XL U15390 ( .A(Q4[14]), .B(n27976), .Y(n27134) );
  OAI21XL U15391 ( .A0(Q5[13]), .A1(n5927), .B0(n27131), .Y(n27582) );
  OAI21XL U15392 ( .A0(n28957), .A1(OP2_done0), .B0(n27130), .Y(n27580) );
  NAND2XL U15393 ( .A(Q4[13]), .B(n27976), .Y(n27130) );
  OAI21XL U15394 ( .A0(Q6[13]), .A1(n5927), .B0(n27131), .Y(n27577) );
  OAI21XL U15395 ( .A0(Q6[12]), .A1(n5927), .B0(n27127), .Y(n27571) );
  OAI21XL U15396 ( .A0(n28956), .A1(n27976), .B0(n27126), .Y(n27574) );
  NAND2XL U15397 ( .A(Q4[12]), .B(n27976), .Y(n27126) );
  OAI21XL U15398 ( .A0(Q6[11]), .A1(n5927), .B0(n27123), .Y(n27565) );
  NAND2XL U15399 ( .A(Q4[11]), .B(n27976), .Y(n27121) );
  AOI22XL U15400 ( .A0(n5840), .A1(CQ1[10]), .B0(Q6[10]), .B1(n27211), .Y(
        n27564) );
  INVXL U15401 ( .A(n27118), .Y(n27562) );
  OAI22XL U15402 ( .A0(n27814), .A1(Q4[10]), .B0(CQ1[10]), .B1(n27976), .Y(
        n27118) );
  AOI22XL U15403 ( .A0(n7123), .A1(CQ1[0]), .B0(Q5[0]), .B1(n27213), .Y(n27498) );
  INVXL U15404 ( .A(n27087), .Y(n27501) );
  OAI22XL U15405 ( .A0(n27814), .A1(Q4[0]), .B0(CQ1[0]), .B1(n27976), .Y(
        n27087) );
  OR2X2 U15406 ( .A(n28707), .B(A_sel_reg[0]), .Y(n7354) );
  NOR2XL U15407 ( .A(n11896), .B(n28665), .Y(n28657) );
  AOI21XL U15408 ( .A0(n27976), .A1(Q3[9]), .B0(n27852), .Y(n28347) );
  OAI2BB1XL U15409 ( .A0N(n27976), .A1N(Q0[9]), .B0(n27851), .Y(n28350) );
  AOI21XL U15410 ( .A0(n27976), .A1(Q3[8]), .B0(n27848), .Y(n28340) );
  OAI2BB1XL U15411 ( .A0N(n27976), .A1N(Q0[8]), .B0(n27847), .Y(n28343) );
  AOI21XL U15412 ( .A0(OP2_done0), .A1(Q3[7]), .B0(n27844), .Y(n28333) );
  OAI2BB1XL U15413 ( .A0N(n27976), .A1N(Q0[7]), .B0(n27843), .Y(n28336) );
  AOI21XL U15414 ( .A0(OP2_done0), .A1(Q3[6]), .B0(n27840), .Y(n28326) );
  OAI2BB1XL U15415 ( .A0N(n27976), .A1N(Q0[6]), .B0(n27839), .Y(n28329) );
  AOI21XL U15416 ( .A0(OP2_done0), .A1(Q3[5]), .B0(n27836), .Y(n28318) );
  OAI2BB1XL U15417 ( .A0N(n27976), .A1N(Q0[5]), .B0(n27835), .Y(n28321) );
  OAI21XL U15418 ( .A0(Q2[53]), .A1(n28053), .B0(n28052), .Y(n28622) );
  OAI2BB1XL U15419 ( .A0N(Q0[53]), .A1N(OP2_done0), .B0(n28051), .Y(n28626) );
  OAI21XL U15420 ( .A0(Q1[53]), .A1(n28053), .B0(n28052), .Y(n28628) );
  OAI21XL U15421 ( .A0(Q2[52]), .A1(n28047), .B0(n28046), .Y(n28621) );
  OAI2BB1XL U15422 ( .A0N(Q0[52]), .A1N(n27976), .B0(n28045), .Y(n28619) );
  OAI21XL U15423 ( .A0(Q1[52]), .A1(n28047), .B0(n28046), .Y(n28616) );
  AOI21XL U15424 ( .A0(OP2_done0), .A1(Q3[4]), .B0(n27832), .Y(n28311) );
  OAI2BB1XL U15425 ( .A0N(n27976), .A1N(Q0[4]), .B0(n27831), .Y(n28314) );
  OAI21XL U15426 ( .A0(Q2[51]), .A1(n28042), .B0(n28041), .Y(n28615) );
  OAI21XL U15427 ( .A0(Q1[51]), .A1(n28042), .B0(n28041), .Y(n28610) );
  OAI2BB1XL U15428 ( .A0N(Q0[51]), .A1N(n27976), .B0(n28040), .Y(n28613) );
  OAI21XL U15429 ( .A0(Q1[50]), .A1(n28037), .B0(n28036), .Y(n28604) );
  OAI2BB1XL U15430 ( .A0N(Q0[50]), .A1N(n27976), .B0(n28035), .Y(n28607) );
  OAI21XL U15431 ( .A0(Q2[50]), .A1(n28037), .B0(n28036), .Y(n28609) );
  OAI21XL U15432 ( .A0(Q1[49]), .A1(n28032), .B0(n28031), .Y(n28598) );
  OAI2BB1XL U15433 ( .A0N(Q0[49]), .A1N(n27976), .B0(n28030), .Y(n28601) );
  OAI21XL U15434 ( .A0(Q2[49]), .A1(n28032), .B0(n28031), .Y(n28603) );
  OAI21XL U15435 ( .A0(Q1[48]), .A1(n28027), .B0(n28026), .Y(n28592) );
  OAI2BB1XL U15436 ( .A0N(Q0[48]), .A1N(n27976), .B0(n28025), .Y(n28595) );
  OAI21XL U15437 ( .A0(Q2[48]), .A1(n28027), .B0(n28026), .Y(n28597) );
  OAI21XL U15438 ( .A0(Q1[47]), .A1(n28022), .B0(n28021), .Y(n28591) );
  OAI21XL U15439 ( .A0(Q2[47]), .A1(n28022), .B0(n28021), .Y(n28586) );
  OAI2BB1XL U15440 ( .A0N(Q0[47]), .A1N(n27976), .B0(n28020), .Y(n28589) );
  OAI21XL U15441 ( .A0(Q2[46]), .A1(n28017), .B0(n28016), .Y(n28580) );
  OAI2BB1XL U15442 ( .A0N(Q0[46]), .A1N(OP2_done0), .B0(n28015), .Y(n28583) );
  OAI21XL U15443 ( .A0(Q1[46]), .A1(n28017), .B0(n28016), .Y(n28585) );
  OAI21XL U15444 ( .A0(Q1[45]), .A1(n28012), .B0(n28011), .Y(n28573) );
  OAI2BB1XL U15445 ( .A0N(Q0[45]), .A1N(OP2_done0), .B0(n28010), .Y(n28576) );
  OAI21XL U15446 ( .A0(Q2[45]), .A1(n28012), .B0(n28011), .Y(n28578) );
  OAI21XL U15447 ( .A0(Q1[44]), .A1(n28007), .B0(n28006), .Y(n28567) );
  OAI2BB1XL U15448 ( .A0N(Q0[44]), .A1N(n27976), .B0(n28005), .Y(n28570) );
  OAI21XL U15449 ( .A0(Q2[44]), .A1(n28007), .B0(n28006), .Y(n28572) );
  OAI21XL U15450 ( .A0(Q2[43]), .A1(n28002), .B0(n28001), .Y(n28566) );
  OAI21XL U15451 ( .A0(Q1[43]), .A1(n28002), .B0(n28001), .Y(n28561) );
  OAI2BB1XL U15452 ( .A0N(Q0[43]), .A1N(n27976), .B0(n28000), .Y(n28564) );
  OAI21XL U15453 ( .A0(Q2[42]), .A1(n27997), .B0(n27996), .Y(n28560) );
  OAI2BB1XL U15454 ( .A0N(Q0[42]), .A1N(n27976), .B0(n27995), .Y(n28558) );
  OAI21XL U15455 ( .A0(Q1[42]), .A1(n27997), .B0(n27996), .Y(n28554) );
  AOI21XL U15456 ( .A0(OP2_done0), .A1(Q3[3]), .B0(n27828), .Y(n28304) );
  OAI2BB1XL U15457 ( .A0N(n27976), .A1N(Q0[3]), .B0(n27827), .Y(n28307) );
  OAI21XL U15458 ( .A0(Q1[41]), .A1(n27992), .B0(n27991), .Y(n28547) );
  OAI2BB1XL U15459 ( .A0N(Q0[41]), .A1N(n27976), .B0(n27990), .Y(n28551) );
  OAI21XL U15460 ( .A0(Q2[41]), .A1(n27992), .B0(n27991), .Y(n28553) );
  OAI21XL U15461 ( .A0(Q1[40]), .A1(n27987), .B0(n27986), .Y(n28546) );
  OAI2BB1XL U15462 ( .A0N(Q0[40]), .A1N(n27976), .B0(n27985), .Y(n28544) );
  OAI21XL U15463 ( .A0(Q2[40]), .A1(n27987), .B0(n27986), .Y(n28540) );
  OAI21XL U15464 ( .A0(Q2[39]), .A1(n27982), .B0(n27981), .Y(n28533) );
  OAI2BB1XL U15465 ( .A0N(Q0[39]), .A1N(OP2_done0), .B0(n27980), .Y(n28537) );
  OAI21XL U15466 ( .A0(Q1[39]), .A1(n27982), .B0(n27981), .Y(n28539) );
  AOI21XL U15467 ( .A0(n27976), .A1(Q3[38]), .B0(n27977), .Y(n28527) );
  OAI2BB1XL U15468 ( .A0N(n27976), .A1N(Q0[38]), .B0(n27975), .Y(n28530) );
  AOI21XL U15469 ( .A0(OP2_done0), .A1(Q3[37]), .B0(n27972), .Y(n28520) );
  OAI2BB1XL U15470 ( .A0N(n27976), .A1N(Q0[37]), .B0(n27971), .Y(n28523) );
  AOI21XL U15471 ( .A0(n27976), .A1(Q3[36]), .B0(n27968), .Y(n28513) );
  OAI2BB1XL U15472 ( .A0N(n27976), .A1N(Q0[36]), .B0(n27967), .Y(n28516) );
  AOI21XL U15473 ( .A0(OP2_done0), .A1(Q3[35]), .B0(n27964), .Y(n28506) );
  OAI2BB1XL U15474 ( .A0N(n27976), .A1N(Q0[35]), .B0(n27963), .Y(n28509) );
  AOI21XL U15475 ( .A0(OP2_done0), .A1(Q3[34]), .B0(n27960), .Y(n28499) );
  OAI2BB1XL U15476 ( .A0N(n27976), .A1N(Q0[34]), .B0(n27958), .Y(n28502) );
  AOI21XL U15477 ( .A0(n27976), .A1(Q3[33]), .B0(n27955), .Y(n28492) );
  OAI2BB1XL U15478 ( .A0N(n27976), .A1N(Q0[33]), .B0(n27954), .Y(n28495) );
  AOI21XL U15479 ( .A0(n27976), .A1(Q3[32]), .B0(n27951), .Y(n28485) );
  OAI2BB1XL U15480 ( .A0N(n27976), .A1N(Q0[32]), .B0(n27950), .Y(n28488) );
  AOI21XL U15481 ( .A0(OP2_done0), .A1(Q3[2]), .B0(n27824), .Y(n28297) );
  OAI2BB1XL U15482 ( .A0N(n27976), .A1N(Q0[2]), .B0(n27823), .Y(n28300) );
  AOI21XL U15483 ( .A0(n27976), .A1(Q3[31]), .B0(n27947), .Y(n28478) );
  OAI2BB1XL U15484 ( .A0N(n27976), .A1N(Q0[31]), .B0(n27946), .Y(n28481) );
  AOI21XL U15485 ( .A0(n27976), .A1(Q3[30]), .B0(n27943), .Y(n28471) );
  OAI2BB1XL U15486 ( .A0N(n27976), .A1N(Q0[30]), .B0(n27942), .Y(n28474) );
  AOI21XL U15487 ( .A0(OP2_done0), .A1(Q3[29]), .B0(n27939), .Y(n28464) );
  OAI2BB1XL U15488 ( .A0N(n27976), .A1N(Q0[29]), .B0(n27938), .Y(n28467) );
  AOI21XL U15489 ( .A0(OP2_done0), .A1(Q3[28]), .B0(n27935), .Y(n28457) );
  OAI2BB1XL U15490 ( .A0N(n27976), .A1N(Q0[28]), .B0(n27934), .Y(n28460) );
  OAI21XL U15491 ( .A0(Q2[25]), .A1(n27931), .B0(n27930), .Y(n28449) );
  OAI2BB1XL U15492 ( .A0N(Q0[25]), .A1N(OP2_done0), .B0(n27929), .Y(n28453) );
  OAI21XL U15493 ( .A0(Q1[25]), .A1(n27931), .B0(n27930), .Y(n28455) );
  OAI21XL U15494 ( .A0(Q1[24]), .A1(n27926), .B0(n27925), .Y(n28443) );
  OAI2BB1XL U15495 ( .A0N(Q0[24]), .A1N(OP2_done0), .B0(n27924), .Y(n28446) );
  OAI21XL U15496 ( .A0(Q2[24]), .A1(n27926), .B0(n27925), .Y(n28448) );
  OAI21XL U15497 ( .A0(Q1[23]), .A1(n27921), .B0(n27920), .Y(n28437) );
  OAI2BB1XL U15498 ( .A0N(Q0[23]), .A1N(OP2_done0), .B0(n27919), .Y(n28440) );
  OAI21XL U15499 ( .A0(Q2[23]), .A1(n27921), .B0(n27920), .Y(n28442) );
  OAI21XL U15500 ( .A0(Q2[22]), .A1(n27916), .B0(n27915), .Y(n28436) );
  OAI21XL U15501 ( .A0(Q1[22]), .A1(n27916), .B0(n27915), .Y(n28431) );
  OAI2BB1XL U15502 ( .A0N(Q0[22]), .A1N(OP2_done0), .B0(n27914), .Y(n28434) );
  OAI21XL U15503 ( .A0(Q2[21]), .A1(n27911), .B0(n27910), .Y(n28425) );
  OAI2BB1XL U15504 ( .A0N(Q0[21]), .A1N(n27976), .B0(n27909), .Y(n28428) );
  OAI21XL U15505 ( .A0(Q1[21]), .A1(n27911), .B0(n27910), .Y(n28430) );
  OAI21XL U15506 ( .A0(Q2[20]), .A1(n27906), .B0(n27905), .Y(n28419) );
  OAI2BB1XL U15507 ( .A0N(Q0[20]), .A1N(n27976), .B0(n27904), .Y(n28422) );
  OAI21XL U15508 ( .A0(Q1[20]), .A1(n27906), .B0(n27905), .Y(n28424) );
  OAI2BB1XL U15509 ( .A0N(n27976), .A1N(Q0[1]), .B0(n27819), .Y(n28292) );
  OAI21XL U15510 ( .A0(Q1[19]), .A1(n27901), .B0(n27900), .Y(n28418) );
  OAI2BB1XL U15511 ( .A0N(Q0[19]), .A1N(n27976), .B0(n27899), .Y(n28416) );
  OAI21XL U15512 ( .A0(Q2[19]), .A1(n27901), .B0(n27900), .Y(n28413) );
  OAI21XL U15513 ( .A0(Q2[18]), .A1(n27896), .B0(n27895), .Y(n28412) );
  OAI2BB1XL U15514 ( .A0N(Q0[18]), .A1N(OP2_done0), .B0(n27894), .Y(n28410) );
  OAI21XL U15515 ( .A0(Q1[18]), .A1(n27896), .B0(n27895), .Y(n28407) );
  OAI21XL U15516 ( .A0(Q1[17]), .A1(n27891), .B0(n27890), .Y(n28401) );
  OAI2BB1XL U15517 ( .A0N(Q0[17]), .A1N(OP2_done0), .B0(n27889), .Y(n28404) );
  OAI21XL U15518 ( .A0(Q2[17]), .A1(n27891), .B0(n27890), .Y(n28406) );
  OAI21XL U15519 ( .A0(Q2[16]), .A1(n27886), .B0(n27885), .Y(n28400) );
  OAI2BB1XL U15520 ( .A0N(Q0[16]), .A1N(OP2_done0), .B0(n27884), .Y(n28398) );
  OAI21XL U15521 ( .A0(Q1[16]), .A1(n27886), .B0(n27885), .Y(n28395) );
  OAI21XL U15522 ( .A0(Q2[15]), .A1(n27881), .B0(n27880), .Y(n28389) );
  OAI2BB1XL U15523 ( .A0N(Q0[15]), .A1N(n27976), .B0(n27879), .Y(n28392) );
  OAI21XL U15524 ( .A0(Q1[14]), .A1(n27876), .B0(n27875), .Y(n28388) );
  OAI2BB1XL U15525 ( .A0N(Q0[14]), .A1N(OP2_done0), .B0(n27874), .Y(n28386) );
  OAI21XL U15526 ( .A0(Q2[14]), .A1(n27876), .B0(n27875), .Y(n28382) );
  OAI21XL U15527 ( .A0(Q1[13]), .A1(n27871), .B0(n27870), .Y(n28381) );
  OAI2BB1XL U15528 ( .A0N(Q0[13]), .A1N(OP2_done0), .B0(n27869), .Y(n28379) );
  OAI21XL U15529 ( .A0(Q2[13]), .A1(n27871), .B0(n27870), .Y(n28375) );
  OAI21XL U15530 ( .A0(Q2[12]), .A1(n27866), .B0(n27865), .Y(n28368) );
  OAI2BB1XL U15531 ( .A0N(Q0[12]), .A1N(OP2_done0), .B0(n27864), .Y(n28372) );
  OAI21XL U15532 ( .A0(Q1[12]), .A1(n27866), .B0(n27865), .Y(n28374) );
  OAI21XL U15533 ( .A0(Q1[11]), .A1(n27861), .B0(n27860), .Y(n28367) );
  OAI2BB1XL U15534 ( .A0N(Q0[11]), .A1N(n27976), .B0(n27859), .Y(n28365) );
  OAI21XL U15535 ( .A0(Q2[11]), .A1(n27861), .B0(n27860), .Y(n28361) );
  AOI21XL U15536 ( .A0(OP2_done0), .A1(Q3[10]), .B0(n27856), .Y(n28355) );
  OAI2BB1XL U15537 ( .A0N(n27976), .A1N(Q0[10]), .B0(n27855), .Y(n28358) );
  AOI21XL U15538 ( .A0(OP2_done0), .A1(Q3[0]), .B0(n27816), .Y(n28282) );
  OAI2BB1XL U15539 ( .A0N(n27976), .A1N(Q0[0]), .B0(n27815), .Y(n28285) );
  NOR2BXL U15540 ( .AN(buffer[0]), .B(n27122), .Y(n28284) );
  AOI21XL U15541 ( .A0(n28640), .A1(n28641), .B0(n15027), .Y(n11910) );
  OR2X2 U15542 ( .A(n11907), .B(n28679), .Y(n7298) );
  NAND3X1 U15543 ( .A(n29110), .B(n29111), .C(cs[2]), .Y(n11913) );
  OAI21XL U15544 ( .A0(n7300), .A1(n28680), .B0(n7299), .Y(n28639) );
  AOI22XL U15545 ( .A0(n7305), .A1(n28703), .B0(n11879), .B1(n11633), .Y(
        n28637) );
  NAND2XL U15546 ( .A(n11611), .B(n11610), .Y(n11609) );
  AOI22X1 U15547 ( .A0(cnt[6]), .A1(n28680), .B0(n28704), .B1(cnt[4]), .Y(
        n7256) );
  INVX4 U15548 ( .A(n11913), .Y(n15027) );
  NOR2XL U15549 ( .A(n28758), .B(n27122), .Y(n15038) );
  NOR2XL U15550 ( .A(n28706), .B(n27122), .Y(n15031) );
  AOI22XL U15551 ( .A0(n11960), .A1(n28630), .B0(cnt[7]), .B1(n11968), .Y(
        n5672) );
  AOI22XL U15552 ( .A0(n11970), .A1(n11969), .B0(cnt[4]), .B1(n11968), .Y(
        n5675) );
  INVXL U15553 ( .A(n12337), .Y(n7752) );
  NOR2X1 U15554 ( .A(n7458), .B(n7384), .Y(n14973) );
  OAI21XL U15555 ( .A0(n7937), .A1(n16782), .B0(n7047), .Y(n7458) );
  NOR3X1 U15556 ( .A(n16785), .B(n7937), .C(n16781), .Y(n7384) );
  OAI2BB1XL U15557 ( .A0N(n5812), .A1N(n14498), .B0(n7237), .Y(n4693) );
  OAI22X1 U15558 ( .A0(n7598), .A1(n7596), .B0(n7707), .B1(U2_A_r_d[25]), .Y(
        n25526) );
  NOR2X1 U15559 ( .A(n25528), .B(n29010), .Y(n7596) );
  OAI21XL U15560 ( .A0(n14897), .A1(U1_A_r_d0[25]), .B0(n7674), .Y(n9723) );
  AOI21X1 U15561 ( .A0(n7645), .A1(n7631), .B0(n7630), .Y(n9549) );
  NOR2XL U15562 ( .A(n7653), .B(n7652), .Y(n7645) );
  AOI211XL U15563 ( .A0(n28673), .A1(n11969), .B0(n11640), .C0(n11966), .Y(
        n11639) );
  NAND2XL U15564 ( .A(n11965), .B(n11964), .Y(n5676) );
  AOI22XL U15565 ( .A0(n28630), .A1(n11967), .B0(cnt[3]), .B1(n11968), .Y(
        n11962) );
  INVX1 U15566 ( .A(n10446), .Y(n10438) );
  NOR2X2 U15567 ( .A(n8202), .B(AOPB[37]), .Y(n10456) );
  NOR2X1 U15568 ( .A(n10474), .B(n10469), .Y(n10461) );
  NOR2X2 U15569 ( .A(n10452), .B(n10456), .Y(n8218) );
  INVXL U15570 ( .A(n10465), .Y(n10453) );
  NAND2XL U15571 ( .A(n10461), .B(n10466), .Y(n10455) );
  NAND2X1 U15572 ( .A(n8202), .B(AOPB[37]), .Y(n10457) );
  INVXL U15573 ( .A(n10456), .Y(n10458) );
  INVXL U15574 ( .A(n10452), .Y(n10466) );
  INVXL U15575 ( .A(n10461), .Y(n10464) );
  AOI21XL U15576 ( .A0(n10438), .A1(n10449), .B0(n10437), .Y(n10439) );
  INVXL U15577 ( .A(n10448), .Y(n10437) );
  NAND2XL U15578 ( .A(n10418), .B(n10436), .Y(n10420) );
  AOI21XL U15579 ( .A0(n10438), .A1(n10427), .B0(n10426), .Y(n10428) );
  INVXL U15580 ( .A(n10492), .Y(n10494) );
  NOR2X2 U15581 ( .A(n10841), .B(n10861), .Y(n8250) );
  INVX1 U15582 ( .A(BOPC[7]), .Y(n8282) );
  INVXL U15583 ( .A(n11156), .Y(n11157) );
  AOI21XL U15584 ( .A0(n11160), .A1(n11156), .B0(n11147), .Y(n11148) );
  INVX1 U15585 ( .A(n11139), .Y(n11131) );
  AOI21X1 U15586 ( .A0(n11131), .A1(n11143), .B0(n11130), .Y(n11132) );
  INVXL U15587 ( .A(n11142), .Y(n11130) );
  NAND2X1 U15588 ( .A(n7060), .B(BOPC[39]), .Y(n11135) );
  AOI21XL U15589 ( .A0(n11131), .A1(n11120), .B0(n11119), .Y(n11121) );
  NAND2X2 U15590 ( .A(n8120), .B(BOPC[34]), .Y(n11169) );
  NAND2X1 U15591 ( .A(n8124), .B(BOPC[32]), .Y(n11182) );
  INVXL U15592 ( .A(n11176), .Y(n11178) );
  NOR2X2 U15593 ( .A(n10654), .B(n10656), .Y(n10646) );
  AOI21XL U15594 ( .A0(n10608), .A1(n10619), .B0(n10607), .Y(n10609) );
  INVXL U15595 ( .A(n10618), .Y(n10607) );
  AOI21XL U15596 ( .A0(n10608), .A1(n10597), .B0(n10596), .Y(n10598) );
  AOI21XL U15597 ( .A0(n10608), .A1(n8276), .B0(n8275), .Y(n8277) );
  NAND2XL U15598 ( .A(n8276), .B(n10606), .Y(n8278) );
  NOR2X1 U15599 ( .A(n8132), .B(BOPB[30]), .Y(n10654) );
  NOR2X1 U15600 ( .A(n10994), .B(n10989), .Y(n10979) );
  NOR2X1 U15601 ( .A(n11003), .B(n11005), .Y(n8316) );
  INVXL U15602 ( .A(n11323), .Y(n11312) );
  INVXL U15603 ( .A(n11340), .Y(n11328) );
  INVXL U15604 ( .A(n11331), .Y(n11333) );
  INVXL U15605 ( .A(n11327), .Y(n11341) );
  NOR2XL U15606 ( .A(n8074), .B(AOPC[30]), .Y(n11362) );
  NOR2X1 U15607 ( .A(n8062), .B(AOPC[34]), .Y(n11344) );
  NAND2X1 U15608 ( .A(n8067), .B(AOPC[32]), .Y(n11358) );
  NOR2X2 U15609 ( .A(n7951), .B(W0[26]), .Y(n10131) );
  NOR2X1 U15610 ( .A(W1[24]), .B(W1[8]), .Y(n9961) );
  NOR2X2 U15611 ( .A(W1[25]), .B(W1[9]), .Y(n9963) );
  NAND2X1 U15612 ( .A(W0[3]), .B(W0[19]), .Y(n9847) );
  NOR2X2 U15613 ( .A(W0[4]), .B(W0[20]), .Y(n9837) );
  INVXL U15614 ( .A(n12011), .Y(n12014) );
  NOR2XL U15615 ( .A(U0_U2_y2[3]), .B(U0_U2_y0[3]), .Y(n12011) );
  INVXL U15616 ( .A(n12018), .Y(n12026) );
  NOR2XL U15617 ( .A(U0_U2_y2[5]), .B(U0_U2_y0[5]), .Y(n12018) );
  NAND2X1 U15618 ( .A(n10461), .B(n8218), .Y(n10447) );
  NAND2X1 U15619 ( .A(n10480), .B(n8214), .Y(n8216) );
  NOR2X2 U15620 ( .A(n10485), .B(n10481), .Y(n8214) );
  NOR2X1 U15621 ( .A(n8108), .B(AOPB[45]), .Y(n10391) );
  NAND2XL U15622 ( .A(n10396), .B(n10401), .Y(n10390) );
  INVXL U15623 ( .A(n10404), .Y(n10406) );
  INVXL U15624 ( .A(n10396), .Y(n10399) );
  NAND2XL U15625 ( .A(n10371), .B(n10355), .Y(n8228) );
  NOR2X1 U15626 ( .A(n8098), .B(AOPB[47]), .Y(n10376) );
  INVXL U15627 ( .A(n10383), .Y(n10372) );
  NOR2X1 U15628 ( .A(n8085), .B(AOPB[28]), .Y(n10507) );
  INVX1 U15629 ( .A(U2_B_i[14]), .Y(n11438) );
  NAND2X1 U15630 ( .A(n7297), .B(n8314), .Y(n7760) );
  NOR2X1 U15631 ( .A(n8186), .B(BOPD[38]), .Y(n10779) );
  NOR2X1 U15632 ( .A(BOPD[14]), .B(n7053), .Y(n7387) );
  INVXL U15633 ( .A(n10849), .Y(n10698) );
  AOI21XL U15634 ( .A0(n10747), .A1(n10751), .B0(n10738), .Y(n10739) );
  INVXL U15635 ( .A(n10750), .Y(n10738) );
  NAND2XL U15636 ( .A(n10746), .B(n10751), .Y(n10740) );
  OAI21XL U15637 ( .A0(n10741), .A1(n10750), .B0(n10742), .Y(n8257) );
  INVXL U15638 ( .A(n10691), .Y(n10734) );
  NOR2XL U15639 ( .A(n8178), .B(BOPD[42]), .Y(n10755) );
  INVXL U15640 ( .A(n10756), .Y(n10758) );
  NAND2XL U15641 ( .A(n8172), .B(BOPD[44]), .Y(n10750) );
  INVXL U15642 ( .A(n10746), .Y(n10749) );
  NOR2X1 U15643 ( .A(n8182), .B(BOPD[39]), .Y(n10785) );
  INVXL U15644 ( .A(n10791), .Y(n10781) );
  NAND2X1 U15645 ( .A(n8182), .B(BOPD[39]), .Y(n10786) );
  NAND2X1 U15646 ( .A(n8186), .B(BOPD[38]), .Y(n10791) );
  NAND2X1 U15647 ( .A(n8192), .B(BOPD[36]), .Y(n10805) );
  INVXL U15648 ( .A(n10798), .Y(n10800) );
  INVXL U15649 ( .A(n10768), .Y(n7386) );
  INVXL U15650 ( .A(n7387), .Y(n10777) );
  OAI21X2 U15651 ( .A0(n10785), .A1(n10791), .B0(n10786), .Y(n10772) );
  NOR2X1 U15652 ( .A(n8121), .B(BOPD[34]), .Y(n10813) );
  INVXL U15653 ( .A(n10830), .Y(n10837) );
  NOR2X2 U15654 ( .A(n11185), .B(n11187), .Y(n11175) );
  NOR2X2 U15655 ( .A(n8282), .B(BOPC[33]), .Y(n11176) );
  OAI21X2 U15656 ( .A0(n11182), .A1(n11176), .B0(n11177), .Y(n7286) );
  INVXL U15657 ( .A(n11096), .Y(n11084) );
  NAND2XL U15658 ( .A(n11092), .B(n11097), .Y(n11086) );
  INVXL U15659 ( .A(n11100), .Y(n11102) );
  INVXL U15660 ( .A(n11092), .Y(n11095) );
  INVXL U15661 ( .A(n11093), .Y(n11094) );
  NAND2XL U15662 ( .A(n8158), .B(BOPC[48]), .Y(n11065) );
  INVXL U15663 ( .A(n11081), .Y(n11071) );
  INVXL U15664 ( .A(n11075), .Y(n11077) );
  INVXL U15665 ( .A(n11187), .Y(n11189) );
  INVXL U15666 ( .A(n10673), .Y(n10529) );
  AOI21XL U15667 ( .A0(n10580), .A1(n10584), .B0(n10571), .Y(n10572) );
  INVXL U15668 ( .A(n10583), .Y(n10571) );
  NAND2XL U15669 ( .A(n10579), .B(n10584), .Y(n10573) );
  NAND2X1 U15670 ( .A(n8126), .B(BOPB[31]), .Y(n10657) );
  INVXL U15671 ( .A(n10656), .Y(n10658) );
  AND2XL U15672 ( .A(n10627), .B(n10631), .Y(n7048) );
  NAND2X1 U15673 ( .A(n8187), .B(BOPB[37]), .Y(n10625) );
  INVXL U15674 ( .A(n10605), .Y(n10619) );
  INVX1 U15675 ( .A(n10616), .Y(n10608) );
  INVXL U15676 ( .A(n10617), .Y(n10606) );
  NAND2X2 U15677 ( .A(n8123), .B(BOPB[32]), .Y(n10651) );
  NAND2X2 U15678 ( .A(n8119), .B(BOPB[34]), .Y(n10640) );
  INVXL U15679 ( .A(n10579), .Y(n10582) );
  INVXL U15680 ( .A(n10570), .Y(n10584) );
  INVXL U15681 ( .A(n10566), .Y(n10555) );
  INVX1 U15682 ( .A(n10664), .Y(n10690) );
  INVXL U15683 ( .A(n10967), .Y(n10956) );
  NOR2X2 U15684 ( .A(n8068), .B(AOPD[32]), .Y(n10998) );
  NAND2XL U15685 ( .A(n10979), .B(n10984), .Y(n10973) );
  INVXL U15686 ( .A(n10974), .Y(n10976) );
  NAND2X1 U15687 ( .A(n8071), .B(AOPD[31]), .Y(n11006) );
  INVXL U15688 ( .A(n10979), .Y(n10982) );
  AOI21XL U15689 ( .A0(n10921), .A1(n10925), .B0(n10912), .Y(n10913) );
  INVXL U15690 ( .A(n10924), .Y(n10912) );
  NAND2XL U15691 ( .A(n10920), .B(n10925), .Y(n10914) );
  INVXL U15692 ( .A(n10920), .Y(n10923) );
  INVXL U15693 ( .A(n10911), .Y(n10925) );
  INVXL U15694 ( .A(n10907), .Y(n8329) );
  INVXL U15695 ( .A(n11015), .Y(n11017) );
  NOR2X2 U15696 ( .A(n5777), .B(AOPD[28]), .Y(n11037) );
  NOR2X1 U15697 ( .A(n8106), .B(AOPC[45]), .Y(n11271) );
  AOI21XL U15698 ( .A0(n11277), .A1(n11281), .B0(n11268), .Y(n11269) );
  INVXL U15699 ( .A(n11280), .Y(n11268) );
  NAND2XL U15700 ( .A(n11276), .B(n11281), .Y(n11270) );
  INVXL U15701 ( .A(n11222), .Y(n11264) );
  INVXL U15702 ( .A(n11276), .Y(n11279) );
  INVXL U15703 ( .A(n11267), .Y(n11281) );
  AOI21XL U15704 ( .A0(n11253), .A1(n11264), .B0(n8346), .Y(n8347) );
  INVXL U15705 ( .A(n11263), .Y(n8346) );
  NOR2X2 U15706 ( .A(n8084), .B(AOPC[28]), .Y(n11391) );
  XOR2X1 U15707 ( .A(n11348), .B(n11347), .Y(U0_U1_z0[8]) );
  NAND2XL U15708 ( .A(n11346), .B(n11345), .Y(n11347) );
  INVXL U15709 ( .A(n11344), .Y(n11346) );
  AND2XL U15710 ( .A(BOPA[38]), .B(BOPA[39]), .Y(n7032) );
  NAND3X1 U15711 ( .A(n7742), .B(n28681), .C(n28713), .Y(n7744) );
  NAND2X1 U15712 ( .A(n9619), .B(BOPA[39]), .Y(n7262) );
  NOR2XL U15713 ( .A(W3[8]), .B(W3[24]), .Y(n9784) );
  NAND2XL U15714 ( .A(n8045), .B(W3[25]), .Y(n10022) );
  NAND2XL U15715 ( .A(n8023), .B(W3[24]), .Y(n10052) );
  INVXL U15716 ( .A(n10051), .Y(n10054) );
  OR2X2 U15717 ( .A(n9837), .B(n9839), .Y(n7556) );
  INVXL U15718 ( .A(n10164), .Y(n10165) );
  INVX1 U15719 ( .A(n10153), .Y(n10193) );
  NAND2XL U15720 ( .A(n9848), .B(n9847), .Y(n10156) );
  INVXL U15721 ( .A(n9846), .Y(n9848) );
  NAND2X2 U15722 ( .A(n8014), .B(W0[20]), .Y(n10147) );
  NAND2X1 U15723 ( .A(W2[10]), .B(W2[26]), .Y(n9939) );
  INVXL U15724 ( .A(n9915), .Y(n9917) );
  NOR2X1 U15725 ( .A(W2[13]), .B(W2[29]), .Y(n9881) );
  NAND2X2 U15726 ( .A(n7946), .B(W2[22]), .Y(n10312) );
  INVXL U15727 ( .A(n9901), .Y(n9903) );
  INVXL U15728 ( .A(n10316), .Y(n10317) );
  NOR2X1 U15729 ( .A(n9963), .B(n9961), .Y(n9957) );
  OAI21X1 U15730 ( .A0(n9968), .A1(n9983), .B0(n9969), .Y(n7392) );
  NAND2XL U15731 ( .A(n8004), .B(W1[30]), .Y(n10251) );
  NAND2X1 U15732 ( .A(n8017), .B(W1[24]), .Y(n10224) );
  NAND2XL U15733 ( .A(n10008), .B(n10007), .Y(n10264) );
  INVXL U15734 ( .A(n10006), .Y(n10008) );
  INVXL U15735 ( .A(n9850), .Y(n9852) );
  NOR2XL U15736 ( .A(n14312), .B(n14317), .Y(n14179) );
  AND2XL U15737 ( .A(U0_U2_y2[10]), .B(U0_U2_y0[10]), .Y(n12045) );
  AND2XL U15738 ( .A(U0_U2_y2[11]), .B(U0_U2_y0[11]), .Y(n12044) );
  AND2XL U15739 ( .A(U0_U2_y2[9]), .B(U0_U2_y0[9]), .Y(n12041) );
  AOI21XL U15740 ( .A0(n12014), .A1(n7994), .B0(n12013), .Y(n12015) );
  AND2XL U15741 ( .A(U0_U2_y2[2]), .B(U0_U2_y0[2]), .Y(n7994) );
  AOI21XL U15742 ( .A0(n12009), .A1(n12008), .B0(n12007), .Y(n12017) );
  AND2XL U15743 ( .A(U0_U2_y2[1]), .B(U0_U2_y0[1]), .Y(n12007) );
  AND2XL U15744 ( .A(U0_U2_y2[6]), .B(U0_U2_y0[6]), .Y(n12028) );
  AOI21XL U15745 ( .A0(n12026), .A1(n12025), .B0(n12024), .Y(n12032) );
  AND2XL U15746 ( .A(U0_U2_y2[4]), .B(U0_U2_y0[4]), .Y(n12025) );
  NAND2XL U15747 ( .A(n12022), .B(n12029), .Y(n12031) );
  INVXL U15748 ( .A(n12020), .Y(n12022) );
  NOR2XL U15749 ( .A(U0_U2_y2[6]), .B(U0_U2_y0[6]), .Y(n12020) );
  NAND2XL U15750 ( .A(n12019), .B(n12026), .Y(n12023) );
  OR2XL U15751 ( .A(U0_U2_y2[4]), .B(U0_U2_y0[4]), .Y(n12019) );
  OAI21XL U15752 ( .A0(n8967), .A1(n8965), .B0(n8968), .Y(n7739) );
  AND2XL U15753 ( .A(U0_U1_y2[9]), .B(U0_U1_y0[9]), .Y(n12437) );
  AND2XL U15754 ( .A(U0_U1_y2[8]), .B(U0_U1_y0[8]), .Y(n12438) );
  AND2XL U15755 ( .A(U0_U1_y2[10]), .B(U0_U1_y0[10]), .Y(n12441) );
  AND2XL U15756 ( .A(U0_U1_y2[5]), .B(U0_U1_y0[5]), .Y(n12421) );
  AND2XL U15757 ( .A(U0_U1_y2[4]), .B(U0_U1_y0[4]), .Y(n12422) );
  AND2XL U15758 ( .A(U0_U1_y2[6]), .B(U0_U1_y0[6]), .Y(n12425) );
  AND2XL U15759 ( .A(U0_U1_y2[3]), .B(U0_U1_y0[3]), .Y(n12412) );
  OR2XL U15760 ( .A(U0_U1_y2[2]), .B(U0_U1_y0[2]), .Y(n12411) );
  AND2XL U15761 ( .A(U0_U1_y2[1]), .B(U0_U1_y0[1]), .Y(n12408) );
  NAND2XL U15762 ( .A(n12418), .B(n12423), .Y(n12420) );
  OR2XL U15763 ( .A(U0_U1_y2[4]), .B(U0_U1_y0[4]), .Y(n12418) );
  NAND2XL U15764 ( .A(n12419), .B(n12426), .Y(n12428) );
  AND2XL U15765 ( .A(U0_U0_y1[2]), .B(U0_U0_y0[2]), .Y(n13199) );
  AND2XL U15766 ( .A(U0_U0_y1[1]), .B(U0_U0_y0[1]), .Y(n13195) );
  OR2XL U15767 ( .A(U0_U0_y1[2]), .B(U0_U0_y0[2]), .Y(n13197) );
  AND2XL U15768 ( .A(U0_U0_y1[7]), .B(U0_U0_y0[7]), .Y(n13211) );
  AND2XL U15769 ( .A(U0_U0_y1[6]), .B(U0_U0_y0[6]), .Y(n13212) );
  AND2XL U15770 ( .A(U0_U0_y1[4]), .B(U0_U0_y0[4]), .Y(n13209) );
  INVXL U15771 ( .A(n13205), .Y(n13206) );
  NOR2XL U15772 ( .A(U0_U0_y1[6]), .B(U0_U0_y0[6]), .Y(n13205) );
  OR2XL U15773 ( .A(U0_U0_y1[4]), .B(U0_U0_y0[4]), .Y(n13204) );
  AOI21XL U15774 ( .A0(n12246), .A1(n7247), .B0(n7246), .Y(n7245) );
  OAI21X1 U15775 ( .A0(n9046), .A1(n9045), .B0(n9044), .Y(n9047) );
  INVXL U15776 ( .A(U0_U1_y1[13]), .Y(n8791) );
  INVX1 U15777 ( .A(U1_U0_y0[27]), .Y(n7632) );
  AND2XL U15778 ( .A(U1_U1_y2[5]), .B(U1_U1_y0[5]), .Y(n12669) );
  AND2XL U15779 ( .A(U1_U1_y2[4]), .B(U1_U1_y0[4]), .Y(n7021) );
  AND2XL U15780 ( .A(U1_U1_y2[6]), .B(U1_U1_y0[6]), .Y(n7017) );
  INVXL U15781 ( .A(n12654), .Y(n12656) );
  NOR2XL U15782 ( .A(U1_U1_y2[2]), .B(U1_U1_y0[2]), .Y(n12654) );
  AND2XL U15783 ( .A(U1_U1_y2[1]), .B(U1_U1_y0[1]), .Y(n12651) );
  AND2XL U15784 ( .A(U1_U1_y2[3]), .B(U1_U1_y0[3]), .Y(n12657) );
  AND2XL U15785 ( .A(U1_U1_y2[2]), .B(U1_U1_y0[2]), .Y(n7020) );
  INVXL U15786 ( .A(n12665), .Y(n12667) );
  NOR2XL U15787 ( .A(U1_U1_y2[6]), .B(U1_U1_y0[6]), .Y(n12665) );
  INVXL U15788 ( .A(n12662), .Y(n12664) );
  NOR2XL U15789 ( .A(U1_U1_y2[4]), .B(U1_U1_y0[4]), .Y(n12662) );
  AND2XL U15790 ( .A(U1_U1_y2[9]), .B(U1_U1_y0[9]), .Y(n12684) );
  AND2XL U15791 ( .A(U1_U1_y2[8]), .B(U1_U1_y0[8]), .Y(n7022) );
  AND2XL U15792 ( .A(U1_U1_y2[10]), .B(U1_U1_y0[10]), .Y(n7013) );
  NOR2X1 U15793 ( .A(n9372), .B(n9370), .Y(n9299) );
  NOR2X2 U15794 ( .A(n9433), .B(n9431), .Y(n7741) );
  NOR2X1 U15795 ( .A(n9357), .B(n9353), .Y(n9361) );
  AND2XL U15796 ( .A(U1_U1_y1[3]), .B(U1_U1_y0[3]), .Y(n14590) );
  AND2XL U15797 ( .A(U1_U1_y1[2]), .B(U1_U1_y0[2]), .Y(n14591) );
  INVXL U15798 ( .A(n14587), .Y(n14589) );
  NOR2XL U15799 ( .A(U1_U1_y1[2]), .B(U1_U1_y0[2]), .Y(n14587) );
  AND2XL U15800 ( .A(U1_U1_y1[4]), .B(U1_U1_y0[4]), .Y(n14602) );
  AOI21XL U15801 ( .A0(n14606), .A1(n14605), .B0(n14604), .Y(n14607) );
  NAND2XL U15802 ( .A(n14599), .B(n14606), .Y(n14608) );
  INVXL U15803 ( .A(n14598), .Y(n14599) );
  NOR2XL U15804 ( .A(U1_U1_y1[6]), .B(U1_U1_y0[6]), .Y(n14598) );
  NAND2XL U15805 ( .A(n14597), .B(n14603), .Y(n14600) );
  INVXL U15806 ( .A(n14596), .Y(n14597) );
  NOR2XL U15807 ( .A(U1_U1_y1[4]), .B(U1_U1_y0[4]), .Y(n14596) );
  AND2XL U15808 ( .A(U1_U1_y1[10]), .B(U1_U1_y0[10]), .Y(n14622) );
  AND2XL U15809 ( .A(U1_U1_y1[11]), .B(U1_U1_y0[11]), .Y(n14621) );
  AND2XL U15810 ( .A(U1_U1_y1[9]), .B(U1_U1_y0[9]), .Y(n14618) );
  INVX1 U15811 ( .A(n13600), .Y(n7277) );
  OAI21XL U15812 ( .A0(n10376), .A1(n10383), .B0(n10377), .Y(n10357) );
  NAND2XL U15813 ( .A(n10352), .B(n10514), .Y(n10353) );
  OAI21X1 U15814 ( .A0(n10522), .A1(n10351), .B0(n10350), .Y(n10354) );
  INVXL U15815 ( .A(n10516), .Y(n10352) );
  NAND2X1 U15816 ( .A(n7758), .B(n7756), .Y(n11549) );
  INVXL U15817 ( .A(n8245), .Y(n7757) );
  INVXL U15818 ( .A(U2_B_r[11]), .Y(n7759) );
  NOR2X1 U15819 ( .A(n9635), .B(U2_B_r[10]), .Y(n11548) );
  NAND2X2 U15820 ( .A(U2_B_i[11]), .B(n7759), .Y(n8147) );
  INVX1 U15821 ( .A(n11548), .Y(n11553) );
  INVX1 U15822 ( .A(U2_B_r[1]), .Y(n7550) );
  NAND2XL U15823 ( .A(BOPD[25]), .B(n8131), .Y(n10848) );
  NOR2X2 U15824 ( .A(n10779), .B(n10785), .Y(n10773) );
  NAND2X2 U15825 ( .A(n8168), .B(BOPD[27]), .Y(n10858) );
  NAND2XL U15826 ( .A(n8154), .B(BOPC[49]), .Y(n11056) );
  INVXL U15827 ( .A(n11210), .Y(n11042) );
  INVXL U15828 ( .A(n11207), .Y(n11043) );
  NOR2XL U15829 ( .A(n8150), .B(BOPB[50]), .Y(n10670) );
  NAND2XL U15830 ( .A(BOPB[25]), .B(n8129), .Y(n10672) );
  NAND2XL U15831 ( .A(n8150), .B(BOPB[50]), .Y(n10673) );
  INVXL U15832 ( .A(n10671), .Y(n9567) );
  NAND2XL U15833 ( .A(AOPD[25]), .B(n8056), .Y(n11022) );
  NAND2XL U15834 ( .A(n11427), .B(BOPA[22]), .Y(n9608) );
  NOR2X2 U15835 ( .A(n9619), .B(n7043), .Y(n7781) );
  NAND2XL U15836 ( .A(n11427), .B(BOPA[13]), .Y(n8690) );
  NOR2XL U15837 ( .A(n11427), .B(n7032), .Y(n7743) );
  INVXL U15838 ( .A(n9784), .Y(n9798) );
  NAND2XL U15839 ( .A(BOPA[20]), .B(n11428), .Y(n11420) );
  OAI21XL U15840 ( .A0(n28685), .A1(n11428), .B0(n11414), .Y(U2_B_r[21]) );
  NAND2XL U15841 ( .A(BOPA[21]), .B(n11430), .Y(n11414) );
  NAND2XL U15842 ( .A(BOPA[19]), .B(n11428), .Y(n9725) );
  NAND2XL U15843 ( .A(BOPA[14]), .B(n11430), .Y(n11409) );
  OAI21XL U15844 ( .A0(n28681), .A1(n11428), .B0(n9622), .Y(U2_B_r[13]) );
  NAND2XL U15845 ( .A(BOPA[13]), .B(n11428), .Y(n9622) );
  NAND2XL U15846 ( .A(BOPA[16]), .B(n11428), .Y(n11406) );
  NAND2X1 U15847 ( .A(n8036), .B(W3[18]), .Y(n10071) );
  NAND2XL U15848 ( .A(n9766), .B(n9765), .Y(n10073) );
  OAI21XL U15849 ( .A0(n28746), .A1(n11430), .B0(n11408), .Y(U2_B_r[15]) );
  NAND2XL U15850 ( .A(BOPA[15]), .B(n11428), .Y(n11408) );
  OAI21X1 U15851 ( .A0(n28750), .A1(n11430), .B0(n9612), .Y(U2_B_r[6]) );
  NAND2XL U15852 ( .A(BOPA[12]), .B(n11430), .Y(n9621) );
  NAND2XL U15853 ( .A(n9782), .B(n9781), .Y(n10062) );
  INVXL U15854 ( .A(n9803), .Y(n9805) );
  AOI21XL U15855 ( .A0(n10103), .A1(n10099), .B0(n10098), .Y(n10100) );
  XNOR2X1 U15856 ( .A(n10089), .B(n10088), .Y(U2_U0_z1[4]) );
  INVXL U15857 ( .A(n10087), .Y(n10088) );
  INVXL U15858 ( .A(n9977), .Y(n9978) );
  INVXL U15859 ( .A(n10238), .Y(n10239) );
  XNOR2XL U15860 ( .A(n10190), .B(n10189), .Y(U0_U0_z1[4]) );
  INVXL U15861 ( .A(n10188), .Y(n10189) );
  INVXL U15862 ( .A(n10166), .Y(n10167) );
  NAND2X1 U15863 ( .A(W2[7]), .B(W2[23]), .Y(n9898) );
  NOR2X2 U15864 ( .A(W2[6]), .B(W2[22]), .Y(n9901) );
  NAND2XL U15865 ( .A(n9943), .B(n9942), .Y(n10334) );
  INVXL U15866 ( .A(n10304), .Y(n10305) );
  INVXL U15867 ( .A(n10332), .Y(n10333) );
  INVXL U15868 ( .A(n10337), .Y(n10338) );
  INVXL U15869 ( .A(n10322), .Y(n10323) );
  NOR2XL U15870 ( .A(n10211), .B(n10208), .Y(n10210) );
  OAI21XL U15871 ( .A0(n10212), .A1(n10208), .B0(n10207), .Y(n10209) );
  INVXL U15872 ( .A(n10244), .Y(n10245) );
  NOR2XL U15873 ( .A(n9072), .B(n9162), .Y(n7776) );
  NAND2XL U15874 ( .A(n24758), .B(n24762), .Y(n24659) );
  NAND3BX2 U15875 ( .AN(n14421), .B(n7594), .C(n7593), .Y(n7592) );
  NOR2X1 U15876 ( .A(n14249), .B(n14248), .Y(n14438) );
  CMPR22X1 U15877 ( .A(U0_U0_y2[28]), .B(U0_U0_y0[28]), .CO(n14242), .S(n14239) );
  CMPR22X1 U15878 ( .A(U0_U0_y2[27]), .B(U0_U0_y0[27]), .CO(n14240), .S(n14237) );
  CMPR22X1 U15879 ( .A(U0_U0_y2[25]), .B(U0_U0_y0[25]), .CO(n14234), .S(n14231) );
  NOR2XL U15880 ( .A(n14178), .B(n14177), .Y(n14309) );
  NAND2XL U15881 ( .A(n14176), .B(n14175), .Y(n14178) );
  AOI21XL U15882 ( .A0(n14167), .A1(n14166), .B0(n14165), .Y(n14168) );
  AOI21XL U15883 ( .A0(n14175), .A1(n14163), .B0(n14162), .Y(n14169) );
  AND2XL U15884 ( .A(U0_U0_y2[11]), .B(U0_U0_y0[11]), .Y(n14165) );
  NOR2XL U15885 ( .A(n14193), .B(n14201), .Y(n14204) );
  CMPR22X1 U15886 ( .A(U0_U1_y2[36]), .B(U0_U1_y0[36]), .CO(n13163), .S(n13156) );
  INVXL U15887 ( .A(n14355), .Y(n14350) );
  NAND2XL U15888 ( .A(n14221), .B(n14220), .Y(n14278) );
  NOR2X1 U15889 ( .A(n14133), .B(U2_A_i_d[20]), .Y(n14129) );
  INVX1 U15890 ( .A(n13447), .Y(n7288) );
  NAND2XL U15891 ( .A(n14086), .B(n7079), .Y(n14094) );
  NOR2X1 U15892 ( .A(n9166), .B(n9162), .Y(n9168) );
  CMPR22X1 U15893 ( .A(U0_U2_y2[16]), .B(U0_U2_y0[16]), .CO(n12063), .S(n12060) );
  AND2XL U15894 ( .A(n12050), .B(U0_U2_y0[13]), .Y(n7961) );
  CMPR22X1 U15895 ( .A(U0_U2_y1[33]), .B(U0_U2_y0[33]), .CO(n9039), .S(n9035)
         );
  CMPR22X1 U15896 ( .A(U0_U2_y1[32]), .B(U0_U2_y0[32]), .CO(n9036), .S(n9031)
         );
  CMPR22X1 U15897 ( .A(U0_U2_y1[31]), .B(U0_U2_y0[31]), .CO(n9032), .S(n9029)
         );
  CMPR22X1 U15898 ( .A(U0_U1_y2[29]), .B(U0_U1_y0[29]), .CO(n12598), .S(n12592) );
  CMPR22X1 U15899 ( .A(U0_U1_y2[28]), .B(U0_U1_y0[28]), .CO(n12593), .S(n12590) );
  CMPR22X1 U15900 ( .A(U0_U2_y1[28]), .B(U0_U2_y0[28]), .CO(n9023), .S(n9020)
         );
  CMPR22X1 U15901 ( .A(U0_U1_y2[27]), .B(U0_U1_y0[27]), .CO(n12591), .S(n12588) );
  CMPR22X1 U15902 ( .A(U0_U2_y1[26]), .B(U0_U2_y0[26]), .CO(n9019), .S(n8995)
         );
  CMPR22X1 U15903 ( .A(U0_U2_y1[22]), .B(U0_U2_y0[22]), .CO(n8955), .S(n8949)
         );
  CMPR22X1 U15904 ( .A(U0_U1_y2[22]), .B(U0_U1_y0[22]), .CO(n12544), .S(n12533) );
  CMPR22X1 U15905 ( .A(U0_U1_y2[23]), .B(U0_U1_y0[23]), .CO(n12546), .S(n12543) );
  AOI21X2 U15906 ( .A0(n12542), .A1(n12541), .B0(n12540), .Y(n13154) );
  NOR2X1 U15907 ( .A(n12531), .B(n12538), .Y(n12542) );
  NAND2X1 U15908 ( .A(n12530), .B(n12536), .Y(n12538) );
  OAI21X1 U15909 ( .A0(n8824), .A1(n8823), .B0(n8822), .Y(n8951) );
  NOR2X1 U15910 ( .A(n8824), .B(n8821), .Y(n8947) );
  AOI21XL U15911 ( .A0(n12448), .A1(n12447), .B0(n7962), .Y(n12498) );
  AND2X1 U15912 ( .A(n12446), .B(U0_U1_y0[13]), .Y(n7962) );
  NOR2XL U15913 ( .A(n8722), .B(n8730), .Y(n8861) );
  NAND2XL U15914 ( .A(n8720), .B(n8725), .Y(n8722) );
  AOI21XL U15915 ( .A0(n8728), .A1(n8727), .B0(n8726), .Y(n8729) );
  AOI21XL U15916 ( .A0(n8725), .A1(n8724), .B0(n8723), .Y(n8731) );
  AND2XL U15917 ( .A(U0_U2_y1[11]), .B(U0_U2_y0[11]), .Y(n8726) );
  AOI21XL U15918 ( .A0(n8718), .A1(n8717), .B0(n8716), .Y(n8859) );
  NOR2X2 U15919 ( .A(n13416), .B(n13421), .Y(n13404) );
  CMPR22X1 U15920 ( .A(U0_U0_y1[27]), .B(U0_U0_y0[27]), .CO(n13268), .S(n13265) );
  CMPR22X1 U15921 ( .A(U0_U0_y1[26]), .B(U0_U0_y0[26]), .CO(n13266), .S(n13263) );
  CMPR22X1 U15922 ( .A(U0_U0_y1[25]), .B(U0_U0_y0[25]), .CO(n13264), .S(n13262) );
  NAND2XL U15923 ( .A(n13388), .B(n13389), .Y(n7607) );
  NAND2XL U15924 ( .A(n13387), .B(n13389), .Y(n7340) );
  XOR2X1 U15925 ( .A(U0_U0_y1[23]), .B(U0_U0_y0[23]), .Y(n13259) );
  NOR2X2 U15926 ( .A(n7569), .B(n13261), .Y(n13366) );
  NAND2X1 U15927 ( .A(n13261), .B(n7569), .Y(n13367) );
  NOR2XL U15928 ( .A(n13227), .B(n13233), .Y(n13334) );
  NAND2XL U15929 ( .A(n13222), .B(n13229), .Y(n13227) );
  AOI21XL U15930 ( .A0(n13229), .A1(n8046), .B0(n13228), .Y(n13234) );
  AOI21XL U15931 ( .A0(n13231), .A1(n7977), .B0(n13230), .Y(n13232) );
  AND2XL U15932 ( .A(U0_U0_y1[8]), .B(U0_U0_y0[8]), .Y(n8046) );
  NAND2X1 U15933 ( .A(n13238), .B(n13221), .Y(n13337) );
  NAND2X1 U15934 ( .A(n12216), .B(n12215), .Y(n12226) );
  OAI21X2 U15935 ( .A0(n9119), .A1(n9128), .B0(n9120), .Y(n9095) );
  CMPR22X1 U15936 ( .A(U0_U1_y1[25]), .B(U0_U1_y0[25]), .CO(n8986), .S(n8983)
         );
  NOR2X1 U15937 ( .A(n8982), .B(n8979), .Y(n9043) );
  CMPR22X1 U15938 ( .A(U0_U1_y1[23]), .B(U0_U1_y0[23]), .CO(n8943), .S(n8939)
         );
  NOR2BX1 U15939 ( .AN(U0_U1_y1[19]), .B(n7772), .Y(n8813) );
  CMPR22X1 U15940 ( .A(U0_U1_y1[17]), .B(U0_U1_y0[17]), .CO(n8807), .S(n8804)
         );
  NOR2XL U15941 ( .A(n8782), .B(n8789), .Y(n8876) );
  NAND2XL U15942 ( .A(n8780), .B(n8785), .Y(n8782) );
  AOI21XL U15943 ( .A0(n8785), .A1(n8784), .B0(n8783), .Y(n8790) );
  AND2XL U15944 ( .A(U0_U1_y1[8]), .B(U0_U1_y0[8]), .Y(n8784) );
  NOR2XL U15945 ( .A(n8765), .B(n8773), .Y(n8776) );
  AND2X1 U15946 ( .A(n8791), .B(U0_U1_y0[13]), .Y(n8792) );
  NOR2X1 U15947 ( .A(n7705), .B(n14429), .Y(n7704) );
  OR2X2 U15948 ( .A(n7592), .B(n14438), .Y(n7591) );
  NAND2XL U15949 ( .A(n14422), .B(n14433), .Y(n7590) );
  AND2X2 U15950 ( .A(U1_U0_y0[28]), .B(U1_U0_y1[28]), .Y(n9321) );
  AOI21XL U15951 ( .A0(n9268), .A1(n9267), .B0(n9266), .Y(n9380) );
  NOR2XL U15952 ( .A(n9256), .B(n9264), .Y(n9267) );
  NOR2XL U15953 ( .A(n9275), .B(n9283), .Y(n9382) );
  NAND2XL U15954 ( .A(n9271), .B(n9278), .Y(n9275) );
  AOI21XL U15955 ( .A0(n9278), .A1(n9277), .B0(n9276), .Y(n9284) );
  AND2XL U15956 ( .A(U1_U0_y1[8]), .B(U1_U0_y0[8]), .Y(n9277) );
  NAND2X1 U15957 ( .A(n7301), .B(n7081), .Y(n8676) );
  CMPR22X1 U15958 ( .A(U1_U1_y2[26]), .B(U1_U1_y0[26]), .CO(n12983), .S(n12942) );
  OAI21X2 U15959 ( .A0(n13016), .A1(n13027), .B0(n13017), .Y(n13062) );
  INVX1 U15960 ( .A(n13057), .Y(n7524) );
  NAND2X1 U15961 ( .A(n6900), .B(n16813), .Y(n7457) );
  NOR2X1 U15962 ( .A(n9292), .B(n9293), .Y(n9404) );
  NAND2X1 U15963 ( .A(n9291), .B(n9290), .Y(n9401) );
  NAND2X1 U15964 ( .A(n9438), .B(n9315), .Y(n9462) );
  INVX1 U15965 ( .A(n9477), .Y(n7698) );
  NAND2X1 U15966 ( .A(n9318), .B(n9319), .Y(n9474) );
  INVXL U15967 ( .A(n9687), .Y(n9697) );
  NOR2XL U15968 ( .A(n9694), .B(U1_A_r_d0[16]), .Y(n9687) );
  NAND2XL U15969 ( .A(n9697), .B(n9688), .Y(n9699) );
  INVXL U15970 ( .A(n19132), .Y(n9688) );
  NOR2XL U15971 ( .A(n8373), .B(n8380), .Y(n8383) );
  NOR2XL U15972 ( .A(n8388), .B(n8396), .Y(n8495) );
  NAND2XL U15973 ( .A(n8386), .B(n8391), .Y(n8388) );
  AOI21XL U15974 ( .A0(n8391), .A1(n8390), .B0(n8389), .Y(n8397) );
  AOI21XL U15975 ( .A0(n8394), .A1(n8393), .B0(n8392), .Y(n8395) );
  NOR2X2 U15976 ( .A(n8596), .B(n8601), .Y(n8588) );
  NOR2XL U15977 ( .A(n13747), .B(n13754), .Y(n13757) );
  NOR2XL U15978 ( .A(n13764), .B(n13769), .Y(n13819) );
  NAND2XL U15979 ( .A(n13761), .B(n13760), .Y(n13764) );
  AOI21XL U15980 ( .A0(n13760), .A1(n13766), .B0(n13765), .Y(n13770) );
  OAI21XL U15981 ( .A0(n12864), .A1(n12866), .B0(n12867), .Y(n12797) );
  NAND2X1 U15982 ( .A(n9366), .B(n9299), .Y(n9352) );
  AOI21XL U15983 ( .A0(n9299), .A1(n9367), .B0(n9298), .Y(n9351) );
  OAI21XL U15984 ( .A0(n9372), .A1(n9376), .B0(n9373), .Y(n9298) );
  NOR2X1 U15985 ( .A(n9300), .B(n9301), .Y(n9357) );
  NOR2X2 U15986 ( .A(n9304), .B(n9305), .Y(n9431) );
  AOI21X1 U15987 ( .A0(n9362), .A1(n9361), .B0(n9360), .Y(n9432) );
  INVX1 U15988 ( .A(n9434), .Y(n7656) );
  NAND3X2 U15989 ( .A(n7658), .B(n9361), .C(n7741), .Y(n7657) );
  NAND2X1 U15990 ( .A(n7659), .B(n9351), .Y(n7658) );
  INVX1 U15991 ( .A(U1_U0_y0[25]), .Y(n7623) );
  CMPR22X1 U15992 ( .A(U1_U0_y1[24]), .B(U1_U0_y0[24]), .CO(n9313), .S(n9310)
         );
  NOR2X2 U15993 ( .A(n9314), .B(n5764), .Y(n9439) );
  NAND2X1 U15994 ( .A(n9472), .B(n7692), .Y(n7691) );
  NOR2XL U15995 ( .A(n7693), .B(n9468), .Y(n7692) );
  AOI21XL U15996 ( .A0(n9463), .A1(n9470), .B0(n7690), .Y(n7689) );
  NAND2X1 U15997 ( .A(n9322), .B(n7029), .Y(n9465) );
  CLKINVX3 U15998 ( .A(n9491), .Y(n9520) );
  NAND2X1 U15999 ( .A(n9327), .B(n9326), .Y(n9493) );
  NOR2X1 U16000 ( .A(n9482), .B(n9481), .Y(n7641) );
  NAND3X1 U16001 ( .A(n5870), .B(n7642), .C(n7680), .Y(n7341) );
  NOR2XL U16002 ( .A(n12720), .B(n12728), .Y(n12731) );
  NAND2XL U16003 ( .A(n12734), .B(n12739), .Y(n12736) );
  AND2XL U16004 ( .A(n12746), .B(U1_U2_y0[13]), .Y(n12747) );
  AND2XL U16005 ( .A(n14627), .B(U1_U1_y0[13]), .Y(n14628) );
  CMPR22X1 U16006 ( .A(U1_U2_y1[16]), .B(U1_U2_y0[16]), .CO(n12760), .S(n12757) );
  OAI21XL U16007 ( .A0(n12871), .A1(n12874), .B0(n12875), .Y(n12808) );
  CMPR22X1 U16008 ( .A(U1_U2_y1[19]), .B(U1_U2_y0[19]), .CO(n12767), .S(n12764) );
  NOR2XL U16009 ( .A(n12908), .B(n12907), .Y(n12946) );
  CMPR22X1 U16010 ( .A(U1_U2_y1[24]), .B(U1_U2_y0[24]), .CO(n12951), .S(n12910) );
  CMPR22X1 U16011 ( .A(U1_U2_y1[26]), .B(U1_U2_y0[26]), .CO(n13001), .S(n12952) );
  NOR2X2 U16012 ( .A(n13020), .B(n13031), .Y(n13040) );
  INVX1 U16013 ( .A(n14805), .Y(n7897) );
  NOR2X1 U16014 ( .A(n7888), .B(n6130), .Y(n7807) );
  NOR2X1 U16015 ( .A(n14840), .B(n14841), .Y(n7258) );
  NOR2XL U16016 ( .A(n9404), .B(n9402), .Y(n9366) );
  OAI21XL U16017 ( .A0(n9404), .A1(n9401), .B0(n9405), .Y(n9367) );
  OAI21XL U16018 ( .A0(n11483), .A1(n11491), .B0(n11484), .Y(n11454) );
  OAI21XL U16019 ( .A0(n11504), .A1(n11514), .B0(n11515), .Y(n11505) );
  NOR2XL U16020 ( .A(n10850), .B(n10846), .Y(n10852) );
  NOR2X2 U16021 ( .A(n8288), .B(n11140), .Y(n7564) );
  NOR2XL U16022 ( .A(n11024), .B(n11020), .Y(n11026) );
  OAI21XL U16023 ( .A0(n10905), .A1(n10872), .B0(n10871), .Y(n11027) );
  AOI21XL U16024 ( .A0(n10870), .A1(n10895), .B0(n10869), .Y(n10871) );
  NOR2XL U16025 ( .A(n11383), .B(n11379), .Y(n11385) );
  OAI21XL U16026 ( .A0(n11261), .A1(n11228), .B0(n11227), .Y(n11386) );
  AOI21XL U16027 ( .A0(n11226), .A1(n11251), .B0(n11225), .Y(n11227) );
  XOR2X1 U16028 ( .A(n7769), .B(BOPA[51]), .Y(n7768) );
  NAND2XL U16029 ( .A(n11427), .B(BOPA[23]), .Y(n11411) );
  NOR2XL U16030 ( .A(n9752), .B(n9757), .Y(n9760) );
  INVXL U16031 ( .A(n9751), .Y(n9739) );
  XOR2XL U16032 ( .A(n9796), .B(n10084), .Y(U2_U0_z2[2]) );
  NAND2XL U16033 ( .A(BOPA[22]), .B(n11430), .Y(n9609) );
  NAND2XL U16034 ( .A(BOPA[25]), .B(n11428), .Y(n11429) );
  NAND2XL U16035 ( .A(BOPA[23]), .B(n11430), .Y(n11412) );
  XNOR2X1 U16036 ( .A(n10103), .B(n10102), .Y(U2_U0_z1[8]) );
  INVXL U16037 ( .A(n10067), .Y(n10068) );
  OAI21XL U16038 ( .A0(n10083), .A1(n10066), .B0(n10065), .Y(n10069) );
  INVXL U16039 ( .A(n10034), .Y(n10035) );
  INVXL U16040 ( .A(n10094), .Y(n10032) );
  NOR2X1 U16041 ( .A(n19248), .B(n14852), .Y(n14854) );
  NOR2X1 U16042 ( .A(n24680), .B(n24681), .Y(n24683) );
  NAND2X1 U16043 ( .A(n7696), .B(n7081), .Y(n9513) );
  NAND2X1 U16044 ( .A(n9471), .B(n9507), .Y(n9509) );
  AOI21XL U16045 ( .A0(n26492), .A1(n26491), .B0(n26490), .Y(n26493) );
  AOI21XL U16046 ( .A0(n23818), .A1(n23817), .B0(n23816), .Y(n23819) );
  NOR2XL U16047 ( .A(n23582), .B(n23586), .Y(n23589) );
  AOI21XL U16048 ( .A0(n26579), .A1(n26578), .B0(n26577), .Y(n26580) );
  AOI21XL U16049 ( .A0(n23837), .A1(n23836), .B0(n23835), .Y(n23838) );
  NOR2XL U16050 ( .A(n23595), .B(n23599), .Y(n23602) );
  AOI21XL U16051 ( .A0(n23886), .A1(n23885), .B0(n23884), .Y(n23887) );
  AOI21XL U16052 ( .A0(n26531), .A1(n26530), .B0(n26529), .Y(n26532) );
  AOI21XL U16053 ( .A0(n23856), .A1(n23855), .B0(n23854), .Y(n23857) );
  AOI21XL U16054 ( .A0(n26551), .A1(n26550), .B0(n26549), .Y(n26552) );
  AOI21XL U16055 ( .A0(n21224), .A1(n21223), .B0(n21222), .Y(n21225) );
  NOR2XL U16056 ( .A(n18231), .B(n18235), .Y(n18238) );
  AOI21XL U16057 ( .A0(n18432), .A1(n18431), .B0(n18430), .Y(n18433) );
  AOI21XL U16058 ( .A0(n21204), .A1(n21203), .B0(n21202), .Y(n21205) );
  AOI21XL U16059 ( .A0(n18508), .A1(n18507), .B0(n18506), .Y(n18509) );
  AOI21XL U16060 ( .A0(n18451), .A1(n18450), .B0(n18449), .Y(n18452) );
  AOI21XL U16061 ( .A0(n21252), .A1(n21251), .B0(n21250), .Y(n21253) );
  AOI21XL U16062 ( .A0(n21155), .A1(n21154), .B0(n21153), .Y(n21156) );
  XOR2X1 U16063 ( .A(U2_U0_y1[20]), .B(U2_U0_y0[20]), .Y(n26081) );
  AND2X2 U16064 ( .A(U2_U0_y0[20]), .B(U2_U0_y1[20]), .Y(n26153) );
  CMPR22X1 U16065 ( .A(U2_U0_y1[21]), .B(U2_U0_y0[21]), .CO(n26188), .S(n26154) );
  XOR2X2 U16066 ( .A(U2_U0_y1[28]), .B(U2_U0_y0[28]), .Y(n26516) );
  NOR2X1 U16067 ( .A(n21413), .B(n21417), .Y(n21420) );
  INVXL U16068 ( .A(n23132), .Y(n17753) );
  CMPR22X1 U16069 ( .A(U2_U0_y2[18]), .B(U2_U0_y0[18]), .CO(n23365), .S(n23322) );
  NOR2XL U16070 ( .A(n18700), .B(n18704), .Y(n18707) );
  NOR2XL U16071 ( .A(U2_U0_y0[11]), .B(U2_U0_y1[11]), .Y(n19051) );
  NOR2XL U16072 ( .A(U2_U0_y0[9]), .B(U2_U0_y1[9]), .Y(n19048) );
  NOR2XL U16073 ( .A(n19042), .B(n19051), .Y(n19054) );
  NOR2XL U16074 ( .A(U2_U0_y0[10]), .B(U2_U0_y1[10]), .Y(n19042) );
  INVX1 U16075 ( .A(n24644), .Y(n24655) );
  INVXL U16076 ( .A(n8921), .Y(n8911) );
  INVXL U16077 ( .A(n12098), .Y(n12093) );
  NAND2XL U16078 ( .A(n22116), .B(n22242), .Y(n22120) );
  NOR2XL U16079 ( .A(n22108), .B(n22110), .Y(n22119) );
  OAI21XL U16080 ( .A0(n24669), .A1(n24731), .B0(n24668), .Y(n24670) );
  AOI21XL U16081 ( .A0(n24735), .A1(n24733), .B0(n24667), .Y(n24668) );
  AOI21XL U16082 ( .A0(n7999), .A1(n24778), .B0(n24635), .Y(n24636) );
  AND2X2 U16083 ( .A(n24634), .B(n24633), .Y(n24635) );
  INVXL U16084 ( .A(n24615), .Y(n24625) );
  INVXL U16085 ( .A(n8917), .Y(n8899) );
  NOR2XL U16086 ( .A(n14147), .B(U2_A_r_d[22]), .Y(n7720) );
  INVXL U16087 ( .A(n13445), .Y(n13459) );
  NOR2XL U16088 ( .A(n14100), .B(U2_A_r_d[18]), .Y(n13445) );
  AOI21XL U16089 ( .A0(n8035), .A1(n9142), .B0(n8034), .Y(n9143) );
  NOR2X1 U16090 ( .A(n14258), .B(n14257), .Y(n14465) );
  NAND2X1 U16091 ( .A(n6948), .B(n25488), .Y(n25508) );
  AOI21XL U16092 ( .A0(n6948), .A1(n25506), .B0(n25505), .Y(n25507) );
  AOI21X1 U16093 ( .A0(n14409), .A1(n14396), .B0(n14395), .Y(n14407) );
  INVXL U16094 ( .A(n14313), .Y(n14314) );
  INVXL U16095 ( .A(n14312), .Y(n14315) );
  INVX1 U16096 ( .A(n13167), .Y(n14572) );
  AND2X1 U16097 ( .A(n14564), .B(n22930), .Y(n14565) );
  AOI21XL U16098 ( .A0(n7016), .A1(n14557), .B0(n14556), .Y(n14558) );
  NAND2X1 U16099 ( .A(n14532), .B(n22926), .Y(n14542) );
  NAND2XL U16100 ( .A(n12461), .B(n12460), .Y(n12519) );
  NOR2XL U16101 ( .A(n21760), .B(n21896), .Y(n21763) );
  NOR2XL U16102 ( .A(n22044), .B(n22050), .Y(n13117) );
  NOR2XL U16103 ( .A(n14382), .B(n25222), .Y(n14385) );
  NAND2XL U16104 ( .A(n14363), .B(n14362), .Y(n14364) );
  INVXL U16105 ( .A(n14361), .Y(n14363) );
  NAND2XL U16106 ( .A(n14300), .B(n14299), .Y(n14301) );
  NAND2XL U16107 ( .A(n14333), .B(n14332), .Y(n14334) );
  XOR2X1 U16108 ( .A(n14330), .B(n14323), .Y(n25281) );
  NAND2XL U16109 ( .A(n14322), .B(n14328), .Y(n14323) );
  INVXL U16110 ( .A(n14329), .Y(n14322) );
  INVXL U16111 ( .A(n9187), .Y(n9156) );
  XNOR2X1 U16112 ( .A(n13161), .B(n13158), .Y(n22958) );
  AOI21XL U16113 ( .A0(n23056), .A1(n23054), .B0(n22927), .Y(n22928) );
  NOR2XL U16114 ( .A(n14100), .B(U2_A_i_d[18]), .Y(n14097) );
  NOR2XL U16115 ( .A(n14078), .B(n22822), .Y(n14081) );
  INVXL U16116 ( .A(n12272), .Y(n12267) );
  XOR2X2 U16117 ( .A(n12264), .B(n6926), .Y(n13167) );
  NAND2X1 U16118 ( .A(n12218), .B(n12217), .Y(n12244) );
  INVXL U16119 ( .A(n9162), .Y(n9075) );
  NOR2X2 U16120 ( .A(n12213), .B(n12214), .Y(n12229) );
  AOI21X1 U16121 ( .A0(n25728), .A1(n25726), .B0(n12171), .Y(n12172) );
  CLKINVX3 U16122 ( .A(n12194), .Y(n12203) );
  NOR2XL U16123 ( .A(n25741), .B(n25739), .Y(n12170) );
  NOR2X1 U16124 ( .A(n12053), .B(U0_U2_y2[13]), .Y(n12111) );
  INVXL U16125 ( .A(n12106), .Y(n12110) );
  INVXL U16126 ( .A(n12102), .Y(n12105) );
  INVXL U16127 ( .A(n12107), .Y(n12108) );
  NAND2XL U16128 ( .A(n14117), .B(n22617), .Y(n14120) );
  NAND3BX1 U16129 ( .AN(n9034), .B(n5821), .C(n9184), .Y(n7335) );
  INVXL U16130 ( .A(n9088), .Y(n9079) );
  NAND2XL U16131 ( .A(n22643), .B(n22638), .Y(n12617) );
  NAND2X2 U16132 ( .A(n5881), .B(n7737), .Y(n7738) );
  NAND2X1 U16133 ( .A(n9184), .B(n5821), .Y(n7737) );
  NAND2X1 U16134 ( .A(n9020), .B(n9021), .Y(n9125) );
  AOI21XL U16135 ( .A0(n6997), .A1(n22660), .B0(n12576), .Y(n12577) );
  NAND2XL U16136 ( .A(n12567), .B(n12566), .Y(n12583) );
  NAND2X1 U16137 ( .A(n8994), .B(n7559), .Y(n9015) );
  INVXL U16138 ( .A(n8992), .Y(n8956) );
  INVX1 U16139 ( .A(n13154), .Y(n12551) );
  INVXL U16140 ( .A(n12559), .Y(n12549) );
  INVXL U16141 ( .A(n8967), .Y(n8969) );
  OAI2BB1X1 U16142 ( .A0N(n8947), .A1N(n8825), .B0(n7222), .Y(n7221) );
  OAI21XL U16143 ( .A0(n8897), .A1(n8896), .B0(n8895), .Y(n8920) );
  XNOR2X1 U16144 ( .A(n12486), .B(n12485), .Y(n22897) );
  NAND2XL U16145 ( .A(n12484), .B(n12483), .Y(n12485) );
  NAND2XL U16146 ( .A(n8842), .B(n8841), .Y(n8843) );
  INVXL U16147 ( .A(n8840), .Y(n8842) );
  INVXL U16148 ( .A(n12496), .Y(n12501) );
  INVXL U16149 ( .A(n12492), .Y(n12495) );
  INVXL U16150 ( .A(n12498), .Y(n12499) );
  INVXL U16151 ( .A(n8864), .Y(n8867) );
  INVXL U16152 ( .A(n8865), .Y(n8866) );
  NAND2XL U16153 ( .A(n8735), .B(U0_U2_y1[13]), .Y(n8870) );
  INVXL U16154 ( .A(n13477), .Y(n13479) );
  NAND2X2 U16155 ( .A(n13269), .B(n13270), .Y(n13410) );
  NAND2X1 U16156 ( .A(n13266), .B(n13265), .Y(n13422) );
  XNOR2X1 U16157 ( .A(n13380), .B(n13379), .Y(n14030) );
  NAND2XL U16158 ( .A(n13378), .B(n13377), .Y(n13379) );
  NAND2X1 U16159 ( .A(n13250), .B(n13251), .Y(n13324) );
  NAND2X1 U16160 ( .A(n13248), .B(n13249), .Y(n13328) );
  INVXL U16161 ( .A(n13317), .Y(n13320) );
  INVXL U16162 ( .A(n13321), .Y(n13329) );
  NOR2X1 U16163 ( .A(n13239), .B(U0_U0_y1[13]), .Y(n13342) );
  INVXL U16164 ( .A(n13336), .Y(n13341) );
  AOI21XL U16165 ( .A0(n13335), .A1(n13334), .B0(n13333), .Y(n13336) );
  INVXL U16166 ( .A(n13332), .Y(n13335) );
  INVXL U16167 ( .A(n13338), .Y(n13339) );
  INVXL U16168 ( .A(n13337), .Y(n13340) );
  INVXL U16169 ( .A(n13353), .Y(n13347) );
  NAND2XL U16170 ( .A(n9217), .B(n9216), .Y(n9225) );
  NAND2X2 U16171 ( .A(n9055), .B(n9054), .Y(n9105) );
  NAND2X1 U16172 ( .A(n9053), .B(n9052), .Y(n9120) );
  NOR2XL U16173 ( .A(n25389), .B(n25387), .Y(n12377) );
  INVXL U16174 ( .A(n8981), .Y(n8941) );
  INVXL U16175 ( .A(n8979), .Y(n8961) );
  INVXL U16176 ( .A(n8974), .Y(n8976) );
  XNOR2X1 U16177 ( .A(n12155), .B(n12154), .Y(n13113) );
  NOR2X1 U16178 ( .A(n8836), .B(n8835), .Y(n8972) );
  NOR2X1 U16179 ( .A(n8812), .B(n8813), .Y(n8833) );
  INVXL U16180 ( .A(n8910), .Y(n8922) );
  NAND2XL U16181 ( .A(n8847), .B(n8846), .Y(n8848) );
  INVXL U16182 ( .A(n8845), .Y(n8847) );
  NAND2XL U16183 ( .A(n12125), .B(n12124), .Y(n12126) );
  INVXL U16184 ( .A(n8880), .Y(n8881) );
  INVXL U16185 ( .A(n8879), .Y(n8882) );
  AND2X2 U16186 ( .A(n14266), .B(n14481), .Y(n7252) );
  XOR2X1 U16187 ( .A(n14495), .B(n14494), .Y(n25125) );
  NAND2XL U16188 ( .A(n14493), .B(n14492), .Y(n14494) );
  INVXL U16189 ( .A(n14491), .Y(n14493) );
  INVXL U16190 ( .A(n14434), .Y(n14436) );
  AND2XL U16191 ( .A(n21764), .B(U2_A_r_d[12]), .Y(n14387) );
  NAND2XL U16192 ( .A(n7542), .B(n7071), .Y(n19766) );
  NAND2X1 U16193 ( .A(n19769), .B(n19827), .Y(n19771) );
  AOI21XL U16194 ( .A0(n19769), .A1(n19826), .B0(n19768), .Y(n19770) );
  NOR2XL U16195 ( .A(n20121), .B(n20119), .Y(n19983) );
  INVXL U16196 ( .A(n14797), .Y(n7893) );
  NAND2XL U16197 ( .A(n7913), .B(n19998), .Y(n20012) );
  AOI21XL U16198 ( .A0(n20108), .A1(n20106), .B0(n19988), .Y(n19989) );
  NOR2XL U16199 ( .A(n17245), .B(n17243), .Y(n9580) );
  NAND2X1 U16200 ( .A(n17217), .B(n17221), .Y(n9590) );
  INVXL U16201 ( .A(n12818), .Y(n12801) );
  NAND2X1 U16202 ( .A(n17335), .B(n17330), .Y(n13562) );
  NAND2X1 U16203 ( .A(n14640), .B(n14641), .Y(n14710) );
  INVX1 U16204 ( .A(n14641), .Y(n7358) );
  NAND2X1 U16205 ( .A(n7839), .B(n13876), .Y(n13892) );
  NAND2X1 U16206 ( .A(n14664), .B(n14665), .Y(n14810) );
  NAND2X1 U16207 ( .A(n7025), .B(n20308), .Y(n20317) );
  AND2XL U16208 ( .A(n9668), .B(U1_A_i_d0[7]), .Y(n9417) );
  NAND2X1 U16209 ( .A(n9321), .B(n9320), .Y(n9469) );
  NAND2XL U16210 ( .A(n13699), .B(n8173), .Y(n9511) );
  INVXL U16211 ( .A(n12822), .Y(n12812) );
  NOR2X1 U16212 ( .A(n12910), .B(n12911), .Y(n12949) );
  NAND2X1 U16213 ( .A(n12910), .B(n12911), .Y(n12947) );
  NAND2XL U16214 ( .A(n12945), .B(n7819), .Y(n7818) );
  NAND2XL U16215 ( .A(n13082), .B(n13578), .Y(n7835) );
  INVXL U16216 ( .A(n7912), .Y(n7907) );
  AOI21XL U16217 ( .A0(n7911), .A1(n7880), .B0(n7909), .Y(n7908) );
  AND2XL U16218 ( .A(n19727), .B(U1_A_r_d0[7]), .Y(n19728) );
  INVXL U16219 ( .A(n9383), .Y(n9388) );
  AOI21XL U16220 ( .A0(n5919), .A1(n9382), .B0(n9381), .Y(n9383) );
  INVXL U16221 ( .A(n9385), .Y(n9386) );
  INVXL U16222 ( .A(n9384), .Y(n9387) );
  NAND2X1 U16223 ( .A(n13901), .B(n13900), .Y(n7184) );
  INVXL U16224 ( .A(n13922), .Y(n13904) );
  NOR2X2 U16225 ( .A(n13901), .B(n13900), .Y(n13918) );
  AOI21X1 U16226 ( .A0(n7837), .A1(n7462), .B0(n7461), .Y(n7460) );
  NAND2XL U16227 ( .A(n13918), .B(n7184), .Y(n7462) );
  NOR2X1 U16228 ( .A(n7837), .B(n7464), .Y(n7461) );
  OAI21XL U16229 ( .A0(n13581), .A1(n13580), .B0(n13579), .Y(n13582) );
  NOR2XL U16230 ( .A(n16718), .B(n8659), .Y(n7217) );
  NAND2XL U16231 ( .A(n16656), .B(n8680), .Y(n8681) );
  NAND2X1 U16232 ( .A(n8676), .B(n16660), .Y(n8678) );
  AOI22XL U16233 ( .A0(n16659), .A1(n8676), .B0(U1_A_i_d0[20]), .B1(n8675), 
        .Y(n8677) );
  NAND2BX1 U16234 ( .AN(n12980), .B(n7822), .Y(n7823) );
  OR2X2 U16235 ( .A(n7826), .B(n7824), .Y(n7832) );
  NAND2XL U16236 ( .A(n12970), .B(n14929), .Y(n14942) );
  INVX1 U16237 ( .A(n13063), .Y(n7514) );
  INVXL U16238 ( .A(n13061), .Y(n12990) );
  INVXL U16239 ( .A(n13934), .Y(n13936) );
  NOR2X1 U16240 ( .A(n16810), .B(n7457), .Y(n7433) );
  NOR2X1 U16241 ( .A(n7457), .B(n16811), .Y(n7455) );
  NAND2XL U16242 ( .A(n9394), .B(n9401), .Y(n9395) );
  INVXL U16243 ( .A(n9402), .Y(n9394) );
  NAND2XL U16244 ( .A(n9406), .B(n9405), .Y(n9407) );
  OAI21XL U16245 ( .A0(n9403), .A1(n9402), .B0(n9401), .Y(n9408) );
  INVXL U16246 ( .A(n9404), .Y(n9406) );
  INVX1 U16247 ( .A(n13669), .Y(n9655) );
  AOI21XL U16248 ( .A0(n6953), .A1(n19155), .B0(n9682), .Y(n9683) );
  NOR2XL U16249 ( .A(n9699), .B(n19127), .Y(n19103) );
  NAND2X1 U16250 ( .A(n5882), .B(n7886), .Y(n7161) );
  INVXL U16251 ( .A(n8499), .Y(n8500) );
  NAND2XL U16252 ( .A(n8508), .B(n8512), .Y(n8509) );
  INVXL U16253 ( .A(n8513), .Y(n8508) );
  NAND2XL U16254 ( .A(n8517), .B(n8516), .Y(n8518) );
  XOR2X1 U16255 ( .A(n8488), .B(n8487), .Y(n12292) );
  NAND2XL U16256 ( .A(n8486), .B(n8485), .Y(n8487) );
  INVXL U16257 ( .A(n8534), .Y(n8476) );
  NOR2XL U16258 ( .A(n16722), .B(n16728), .Y(n8556) );
  INVX1 U16259 ( .A(n7543), .Y(n7542) );
  INVXL U16260 ( .A(n13821), .Y(n13825) );
  AOI21XL U16261 ( .A0(n13820), .A1(n13819), .B0(n13818), .Y(n13821) );
  INVXL U16262 ( .A(n13817), .Y(n13820) );
  INVXL U16263 ( .A(n13823), .Y(n13824) );
  INVXL U16264 ( .A(n12830), .Y(n12835) );
  AOI21XL U16265 ( .A0(n12829), .A1(n12828), .B0(n12827), .Y(n12830) );
  INVXL U16266 ( .A(n12826), .Y(n12829) );
  INVXL U16267 ( .A(n12832), .Y(n12833) );
  INVXL U16268 ( .A(n12831), .Y(n12834) );
  NOR2X1 U16269 ( .A(n12692), .B(U1_U1_y2[13]), .Y(n12836) );
  NAND2XL U16270 ( .A(n13839), .B(n13838), .Y(n13840) );
  INVXL U16271 ( .A(n12922), .Y(n12924) );
  INVXL U16272 ( .A(n13865), .Y(n13867) );
  OAI21X1 U16273 ( .A0(n9403), .A1(n9352), .B0(n9351), .Y(n9362) );
  NAND4X1 U16274 ( .A(n7655), .B(n7660), .C(n7657), .D(n7614), .Y(n7613) );
  NOR2X2 U16275 ( .A(n9312), .B(n9313), .Y(n9444) );
  INVXL U16276 ( .A(n12845), .Y(n12850) );
  AOI21XL U16277 ( .A0(n12844), .A1(n12843), .B0(n12842), .Y(n12845) );
  INVXL U16278 ( .A(n12841), .Y(n12844) );
  INVXL U16279 ( .A(n12847), .Y(n12848) );
  NOR2X1 U16280 ( .A(n14631), .B(U1_U1_y1[13]), .Y(n14726) );
  INVXL U16281 ( .A(n14720), .Y(n14725) );
  INVXL U16282 ( .A(n14716), .Y(n14719) );
  XNOR2X1 U16283 ( .A(n14744), .B(n14743), .Y(n19956) );
  NAND2XL U16284 ( .A(n14742), .B(n14741), .Y(n14743) );
  NAND2XL U16285 ( .A(n14638), .B(n14639), .Y(n14713) );
  OAI21XL U16286 ( .A0(n14740), .A1(n14709), .B0(n14708), .Y(n14715) );
  OAI21XL U16287 ( .A0(n14738), .A1(n7793), .B0(n14741), .Y(n14707) );
  NAND2X1 U16288 ( .A(n12760), .B(n12759), .Y(n12822) );
  AOI21XL U16289 ( .A0(n12790), .A1(n12900), .B0(n12904), .Y(n12929) );
  NAND2XL U16290 ( .A(n12908), .B(n12907), .Y(n12948) );
  NAND3X2 U16291 ( .A(n7202), .B(n7448), .C(n12900), .Y(n7201) );
  INVXL U16292 ( .A(n14769), .Y(n14771) );
  NAND2X1 U16293 ( .A(n12951), .B(n12950), .Y(n12995) );
  NOR2X1 U16294 ( .A(n13001), .B(n13000), .Y(n13031) );
  NAND2X1 U16295 ( .A(n13002), .B(n13003), .Y(n13021) );
  NAND2X1 U16296 ( .A(n7802), .B(n7894), .Y(n7441) );
  NAND2XL U16297 ( .A(n13603), .B(n13565), .Y(n7500) );
  NAND2XL U16298 ( .A(n7912), .B(n13565), .Y(n7499) );
  NOR2X1 U16299 ( .A(n13567), .B(n13568), .Y(n7174) );
  NAND2XL U16300 ( .A(n27814), .B(n28922), .Y(n11985) );
  INVX2 U16301 ( .A(U2_B_i[0]), .Y(n11603) );
  OR2X2 U16302 ( .A(n7987), .B(n6897), .Y(n7765) );
  INVX1 U16303 ( .A(n7959), .Y(n7406) );
  XOR2X1 U16304 ( .A(n9200), .B(n9214), .Y(n24676) );
  NAND2XL U16305 ( .A(n9199), .B(n9212), .Y(n9200) );
  INVXL U16306 ( .A(n9213), .Y(n9199) );
  NAND2X1 U16307 ( .A(n20337), .B(n20336), .Y(n7872) );
  NAND2X1 U16308 ( .A(n7669), .B(n9535), .Y(n17462) );
  NOR2X1 U16309 ( .A(n9509), .B(n17502), .Y(n17478) );
  AOI2BB2X1 U16310 ( .B0(n9513), .B1(n17481), .A0N(n7696), .A1N(n7081), .Y(
        n9514) );
  NOR2X1 U16311 ( .A(n7751), .B(n7315), .Y(n7314) );
  INVXL U16312 ( .A(n7751), .Y(n7312) );
  NAND2BX1 U16313 ( .AN(n9344), .B(n7664), .Y(n7663) );
  INVXL U16314 ( .A(n9533), .Y(n9344) );
  NOR3XL U16315 ( .A(n28705), .B(n28679), .C(n11963), .Y(n11961) );
  NOR2XL U16316 ( .A(n26566), .B(n26565), .Y(n26629) );
  NOR2XL U16317 ( .A(n26500), .B(n26499), .Y(n26626) );
  NOR2XL U16318 ( .A(n26437), .B(n26436), .Y(n26489) );
  NOR2XL U16319 ( .A(n26388), .B(n26387), .Y(n26484) );
  AOI21XL U16320 ( .A0(n26263), .A1(n26262), .B0(n26261), .Y(n26495) );
  NAND2XL U16321 ( .A(n26257), .B(n26263), .Y(n26486) );
  NOR2XL U16322 ( .A(n26210), .B(n26209), .Y(n26260) );
  NOR2XL U16323 ( .A(n26173), .B(n26172), .Y(n26256) );
  AOI21XL U16324 ( .A0(n26318), .A1(n26317), .B0(n26316), .Y(n26554) );
  NAND2XL U16325 ( .A(n26312), .B(n26318), .Y(n26545) );
  NOR2XL U16326 ( .A(n26282), .B(n26281), .Y(n26315) );
  NOR2XL U16327 ( .A(n26232), .B(n26231), .Y(n26311) );
  NOR2XL U16328 ( .A(n25978), .B(n25977), .Y(n25996) );
  AOI21XL U16329 ( .A0(n25931), .A1(n25930), .B0(n25929), .Y(n26136) );
  NOR2XL U16330 ( .A(n25925), .B(n25928), .Y(n25931) );
  NOR2XL U16331 ( .A(n25933), .B(n25932), .Y(n25993) );
  NOR2XL U16332 ( .A(n23917), .B(n23916), .Y(n23972) );
  NOR2XL U16333 ( .A(n23826), .B(n23825), .Y(n23969) );
  NOR2XL U16334 ( .A(n23765), .B(n23764), .Y(n23815) );
  NOR2XL U16335 ( .A(n23736), .B(n23735), .Y(n23810) );
  NOR2XL U16336 ( .A(n23565), .B(n23564), .Y(n23586) );
  NOR2XL U16337 ( .A(n23521), .B(n23520), .Y(n23582) );
  NOR2XL U16338 ( .A(n26507), .B(n26506), .Y(n26576) );
  NOR2XL U16339 ( .A(n26430), .B(n26429), .Y(n26571) );
  AOI21XL U16340 ( .A0(n26340), .A1(n26339), .B0(n26338), .Y(n26582) );
  NAND2XL U16341 ( .A(n26334), .B(n26340), .Y(n26573) );
  NOR2XL U16342 ( .A(n26251), .B(n26250), .Y(n26337) );
  NOR2XL U16343 ( .A(n26203), .B(n26202), .Y(n26333) );
  NOR2XL U16344 ( .A(n25952), .B(n25951), .Y(n26023) );
  AOI21XL U16345 ( .A0(n25901), .A1(n25900), .B0(n25899), .Y(n26098) );
  NOR2XL U16346 ( .A(n25895), .B(n25898), .Y(n25901) );
  NOR2XL U16347 ( .A(n25903), .B(n25902), .Y(n26020) );
  NOR2XL U16348 ( .A(n23909), .B(n23908), .Y(n23962) );
  NOR2XL U16349 ( .A(n23845), .B(n23844), .Y(n23959) );
  NOR2XL U16350 ( .A(n23774), .B(n23773), .Y(n23834) );
  NOR2XL U16351 ( .A(n23725), .B(n23724), .Y(n23829) );
  NOR2XL U16352 ( .A(n23545), .B(n23544), .Y(n23599) );
  NOR2XL U16353 ( .A(n23505), .B(n23504), .Y(n23595) );
  NOR2XL U16354 ( .A(n23805), .B(n23804), .Y(n23883) );
  NOR2XL U16355 ( .A(n23758), .B(n23757), .Y(n23878) );
  AOI21XL U16356 ( .A0(n23648), .A1(n23647), .B0(n23646), .Y(n23889) );
  NAND2XL U16357 ( .A(n23642), .B(n23648), .Y(n23880) );
  NOR2XL U16358 ( .A(n23612), .B(n23611), .Y(n23645) );
  NOR2XL U16359 ( .A(n23557), .B(n23556), .Y(n23641) );
  NOR2XL U16360 ( .A(n23304), .B(n23303), .Y(n23346) );
  NOR2XL U16361 ( .A(n23249), .B(n23252), .Y(n23255) );
  NOR2XL U16362 ( .A(n23257), .B(n23256), .Y(n23343) );
  NOR2XL U16363 ( .A(n26470), .B(n26469), .Y(n26528) );
  NOR2XL U16364 ( .A(n26419), .B(n26418), .Y(n26523) );
  AOI21XL U16365 ( .A0(n26305), .A1(n26304), .B0(n26303), .Y(n26534) );
  NAND2XL U16366 ( .A(n26299), .B(n26305), .Y(n26525) );
  NOR2XL U16367 ( .A(n26273), .B(n26272), .Y(n26302) );
  NOR2XL U16368 ( .A(n26222), .B(n26221), .Y(n26298) );
  NOR2XL U16369 ( .A(n25970), .B(n25969), .Y(n26013) );
  AOI21XL U16370 ( .A0(n25920), .A1(n25919), .B0(n25918), .Y(n26120) );
  NOR2XL U16371 ( .A(n25914), .B(n25917), .Y(n25920) );
  NOR2XL U16372 ( .A(n25922), .B(n25921), .Y(n26010) );
  NOR2XL U16373 ( .A(n23901), .B(n23900), .Y(n23952) );
  NOR2XL U16374 ( .A(n23783), .B(n23782), .Y(n23853) );
  NOR2XL U16375 ( .A(n23714), .B(n23713), .Y(n23848) );
  AOI21XL U16376 ( .A0(n23624), .A1(n23623), .B0(n23622), .Y(n23859) );
  NAND2XL U16377 ( .A(n23618), .B(n23624), .Y(n23850) );
  NOR2XL U16378 ( .A(n23488), .B(n23491), .Y(n23618) );
  NOR2XL U16379 ( .A(n26479), .B(n26478), .Y(n26548) );
  NOR2XL U16380 ( .A(n26450), .B(n26449), .Y(n26543) );
  NOR2XL U16381 ( .A(n21115), .B(n21114), .Y(n21216) );
  NOR2XL U16382 ( .A(n21170), .B(n21169), .Y(n21221) );
  NOR2XL U16383 ( .A(n17805), .B(n17804), .Y(n17923) );
  NOR2XL U16384 ( .A(n17853), .B(n17852), .Y(n17926) );
  AOI21XL U16385 ( .A0(n17803), .A1(n17802), .B0(n17801), .Y(n17995) );
  NOR2XL U16386 ( .A(n17800), .B(n17797), .Y(n17803) );
  NOR2XL U16387 ( .A(n18107), .B(n18106), .Y(n18231) );
  NOR2XL U16388 ( .A(n18152), .B(n18151), .Y(n18235) );
  NOR2XL U16389 ( .A(n18327), .B(n18326), .Y(n18424) );
  NOR2XL U16390 ( .A(n18399), .B(n18398), .Y(n18429) );
  NOR2XL U16391 ( .A(n18523), .B(n18522), .Y(n18584) );
  NOR2XL U16392 ( .A(n18440), .B(n18439), .Y(n18581) );
  NOR2XL U16393 ( .A(n20587), .B(n20586), .Y(n20674) );
  NOR2XL U16394 ( .A(n20632), .B(n20631), .Y(n20677) );
  AOI21XL U16395 ( .A0(n20585), .A1(n20584), .B0(n20583), .Y(n20790) );
  NOR2XL U16396 ( .A(n20579), .B(n20582), .Y(n20585) );
  AOI21XL U16397 ( .A0(n20972), .A1(n20971), .B0(n20970), .Y(n21207) );
  NAND2XL U16398 ( .A(n20966), .B(n20972), .Y(n21198) );
  NOR2XL U16399 ( .A(n21084), .B(n21083), .Y(n21196) );
  NOR2XL U16400 ( .A(n21133), .B(n21132), .Y(n21201) );
  NOR2XL U16401 ( .A(n17874), .B(n17873), .Y(n17959) );
  NOR2XL U16402 ( .A(n17918), .B(n17917), .Y(n17962) );
  AOI21XL U16403 ( .A0(n17872), .A1(n17871), .B0(n17870), .Y(n18080) );
  NOR2XL U16404 ( .A(n17866), .B(n17869), .Y(n17872) );
  AOI21XL U16405 ( .A0(n18266), .A1(n18265), .B0(n18264), .Y(n18511) );
  NAND2XL U16406 ( .A(n18260), .B(n18266), .Y(n18502) );
  NOR2XL U16407 ( .A(n18374), .B(n18373), .Y(n18500) );
  NOR2XL U16408 ( .A(n18419), .B(n18418), .Y(n18505) );
  AOI21XL U16409 ( .A0(n18216), .A1(n18215), .B0(n18214), .Y(n18454) );
  NAND2XL U16410 ( .A(n18210), .B(n18216), .Y(n18445) );
  NOR2XL U16411 ( .A(n18219), .B(n18218), .Y(n18330) );
  NOR2XL U16412 ( .A(n18285), .B(n18284), .Y(n18333) );
  NOR2XL U16413 ( .A(n18330), .B(n18333), .Y(n18444) );
  NOR2XL U16414 ( .A(n18531), .B(n18530), .Y(n18574) );
  NOR2XL U16415 ( .A(n18459), .B(n18458), .Y(n18571) );
  NOR2XL U16416 ( .A(n20568), .B(n20567), .Y(n20684) );
  NOR2XL U16417 ( .A(n20640), .B(n20639), .Y(n20687) );
  AOI21XL U16418 ( .A0(n20566), .A1(n20565), .B0(n20564), .Y(n20768) );
  NOR2XL U16419 ( .A(n20560), .B(n20563), .Y(n20566) );
  AOI21XL U16420 ( .A0(n20985), .A1(n20984), .B0(n20983), .Y(n21255) );
  NAND2XL U16421 ( .A(n20979), .B(n20985), .Y(n21246) );
  NOR2XL U16422 ( .A(n21095), .B(n21094), .Y(n21244) );
  NOR2XL U16423 ( .A(n21142), .B(n21141), .Y(n21249) );
  NOR2XL U16424 ( .A(n17834), .B(n17833), .Y(n17895) );
  NOR2XL U16425 ( .A(n17880), .B(n17879), .Y(n17898) );
  NOR2XL U16426 ( .A(n18180), .B(n18179), .Y(n18200) );
  NOR2XL U16427 ( .A(n18478), .B(n18477), .Y(n18561) );
  INVXL U16428 ( .A(n18638), .Y(n18639) );
  NAND2XL U16429 ( .A(n18637), .B(n18565), .Y(n18667) );
  NOR2XL U16430 ( .A(n18644), .B(n18643), .Y(n18669) );
  AOI21XL U16431 ( .A0(n18476), .A1(n18475), .B0(n18474), .Y(n18734) );
  NOR2XL U16432 ( .A(n18464), .B(n18472), .Y(n18475) );
  NAND2XL U16433 ( .A(n18463), .B(n18470), .Y(n18472) );
  NOR2XL U16434 ( .A(n20598), .B(n20597), .Y(n20657) );
  NOR2XL U16435 ( .A(n20614), .B(n20613), .Y(n20660) );
  AOI21XL U16436 ( .A0(n20596), .A1(n20595), .B0(n20594), .Y(n20806) );
  NOR2XL U16437 ( .A(n20590), .B(n20593), .Y(n20596) );
  AOI21XL U16438 ( .A0(n21007), .A1(n21006), .B0(n21005), .Y(n21227) );
  NAND2XL U16439 ( .A(n21001), .B(n21007), .Y(n21218) );
  NOR2XL U16440 ( .A(n20574), .B(n20573), .Y(n20622) );
  AOI21XL U16441 ( .A0(n20926), .A1(n20925), .B0(n20924), .Y(n21158) );
  NAND2XL U16442 ( .A(n20920), .B(n20926), .Y(n21149) );
  NOR2XL U16443 ( .A(n21051), .B(n21050), .Y(n21147) );
  NOR2XL U16444 ( .A(n21102), .B(n21101), .Y(n21152) );
  NOR2XL U16445 ( .A(n21239), .B(n21238), .Y(n21290) );
  NOR2XL U16446 ( .A(n21163), .B(n21162), .Y(n21287) );
  AOI21XL U16447 ( .A0(n20528), .A1(n20527), .B0(n20526), .Y(n20720) );
  NOR2XL U16448 ( .A(n20525), .B(n20522), .Y(n20528) );
  NOR2XL U16449 ( .A(n20530), .B(n20529), .Y(n20619) );
  INVX1 U16450 ( .A(n26755), .Y(n7549) );
  NOR2X1 U16451 ( .A(n26754), .B(n26817), .Y(n7547) );
  INVX1 U16452 ( .A(n26906), .Y(n7540) );
  OAI21XL U16453 ( .A0(n23791), .A1(n23790), .B0(n23789), .Y(n23929) );
  XNOR2XL U16454 ( .A(n20469), .B(n20468), .Y(n19065) );
  INVXL U16455 ( .A(n25888), .Y(n20555) );
  NOR2XL U16456 ( .A(n20557), .B(n20556), .Y(n20645) );
  INVX1 U16457 ( .A(n26241), .Y(n20902) );
  NOR2X1 U16458 ( .A(n20905), .B(n20904), .Y(n20954) );
  INVX1 U16459 ( .A(n26403), .Y(n21070) );
  NOR2XL U16460 ( .A(n21063), .B(n21066), .Y(n21176) );
  INVXL U16461 ( .A(n16617), .Y(n16618) );
  NAND2XL U16462 ( .A(n17752), .B(U2_U0_y0[13]), .Y(n16614) );
  AOI21XL U16463 ( .A0(n16613), .A1(n16612), .B0(n16611), .Y(n16620) );
  NOR2XL U16464 ( .A(U2_U0_y0[12]), .B(U2_U0_y2[12]), .Y(n16603) );
  NAND2XL U16465 ( .A(n16602), .B(n16613), .Y(n16604) );
  NOR2XL U16466 ( .A(n16600), .B(n16607), .Y(n16602) );
  NOR2XL U16467 ( .A(U2_U0_y0[8]), .B(U2_U0_y2[8]), .Y(n16600) );
  AOI21XL U16468 ( .A0(n16596), .A1(n16595), .B0(n16594), .Y(n16597) );
  XNOR2XL U16469 ( .A(n17753), .B(n17752), .Y(n16624) );
  INVXL U16470 ( .A(n23225), .Y(n17845) );
  INVXL U16471 ( .A(n23224), .Y(n17844) );
  INVXL U16472 ( .A(n23275), .Y(n17887) );
  NOR2X1 U16473 ( .A(n17890), .B(n17889), .Y(n17936) );
  OAI21XL U16474 ( .A0(n18139), .A1(n18138), .B0(n18137), .Y(n18250) );
  INVX1 U16475 ( .A(n23795), .Y(n18407) );
  INVX1 U16476 ( .A(n23796), .Y(n18408) );
  ADDFX2 U16477 ( .A(n18907), .B(n18906), .CI(U2_A_i_d[22]), .CO(n18908), .S(
        n18867) );
  ADDFX2 U16478 ( .A(n25944), .B(n25943), .CI(U2_A_r_d[3]), .CO(n25945), .S(
        n25890) );
  ADDFX2 U16479 ( .A(n25986), .B(n25985), .CI(U2_A_r_d[4]), .CO(n25987), .S(
        n25946) );
  NOR2XL U16480 ( .A(n25946), .B(n25945), .Y(n26030) );
  INVXL U16481 ( .A(n19058), .Y(n19059) );
  NAND2XL U16482 ( .A(n20468), .B(U2_U0_y0[13]), .Y(n19055) );
  NOR2XL U16483 ( .A(U2_U0_y0[12]), .B(U2_U0_y1[12]), .Y(n19044) );
  NAND2XL U16484 ( .A(n19043), .B(n19054), .Y(n19045) );
  NOR2XL U16485 ( .A(n19041), .B(n19048), .Y(n19043) );
  NOR2XL U16486 ( .A(U2_U0_y0[8]), .B(U2_U0_y1[8]), .Y(n19041) );
  AOI21XL U16487 ( .A0(n19037), .A1(n19036), .B0(n19035), .Y(n19038) );
  AOI21X1 U16488 ( .A0(n25040), .A1(n25038), .B0(n9137), .Y(n25028) );
  NAND2XL U16489 ( .A(n24469), .B(n24473), .Y(n13998) );
  INVX1 U16490 ( .A(n24921), .Y(n7326) );
  NAND2XL U16491 ( .A(n24509), .B(n13507), .Y(n13513) );
  INVXL U16492 ( .A(n24946), .Y(n13503) );
  INVXL U16493 ( .A(n24767), .Y(n24651) );
  AOI21XL U16494 ( .A0(n24811), .A1(n24585), .B0(n24612), .Y(n24613) );
  INVXL U16495 ( .A(n24813), .Y(n24612) );
  AOI21XL U16496 ( .A0(n13459), .A1(n24466), .B0(n13458), .Y(n24452) );
  AND2X1 U16497 ( .A(n14100), .B(U2_A_r_d[18]), .Y(n13458) );
  NAND2XL U16498 ( .A(n13459), .B(n24467), .Y(n24453) );
  NAND2X1 U16499 ( .A(n24507), .B(n13399), .Y(n7603) );
  NAND2X1 U16500 ( .A(n7600), .B(n7037), .Y(n7599) );
  NAND2XL U16501 ( .A(n13398), .B(U2_A_r_d[12]), .Y(n7037) );
  NAND2XL U16502 ( .A(n13397), .B(n13396), .Y(n7586) );
  NAND2X1 U16503 ( .A(n7589), .B(n13363), .Y(n24503) );
  INVXL U16504 ( .A(n24540), .Y(n13362) );
  INVXL U16505 ( .A(n24930), .Y(n24533) );
  NOR2X1 U16506 ( .A(n24677), .B(n24687), .Y(n24704) );
  NAND2XL U16507 ( .A(n14356), .B(n14355), .Y(n14357) );
  NAND2XL U16508 ( .A(n14542), .B(n22028), .Y(n14544) );
  NAND2XL U16509 ( .A(n14541), .B(n14531), .Y(n22026) );
  INVXL U16510 ( .A(n22061), .Y(n14528) );
  OAI21XL U16511 ( .A0(n21755), .A1(n21910), .B0(n21754), .Y(n21881) );
  AOI21XL U16512 ( .A0(n21911), .A1(n21753), .B0(n21752), .Y(n21754) );
  INVXL U16513 ( .A(n22329), .Y(n13130) );
  NOR2XL U16514 ( .A(n22363), .B(n13120), .Y(n13121) );
  OAI21XL U16515 ( .A0(n14348), .A1(n25239), .B0(n14347), .Y(n25207) );
  AOI21XL U16516 ( .A0(n25240), .A1(n14346), .B0(n14345), .Y(n14347) );
  INVX1 U16517 ( .A(n25251), .Y(n21748) );
  INVXL U16518 ( .A(n25281), .Y(n21735) );
  NAND2XL U16519 ( .A(n23043), .B(n22937), .Y(n23026) );
  XOR2XL U16520 ( .A(n13298), .B(n13297), .Y(n13299) );
  AOI2BB1X1 U16521 ( .A0N(n14097), .A1N(n7292), .B0(n14101), .Y(n7296) );
  AND2X2 U16522 ( .A(n14100), .B(U2_A_i_d[18]), .Y(n14101) );
  NAND2BX1 U16523 ( .AN(n14097), .B(n14098), .Y(n14131) );
  NAND2XL U16524 ( .A(n22840), .B(n22842), .Y(n14070) );
  INVXL U16525 ( .A(n22841), .Y(n14068) );
  INVXL U16526 ( .A(n14018), .Y(n14057) );
  AOI21XL U16527 ( .A0(n25339), .A1(n12236), .B0(n12235), .Y(n25681) );
  NAND2XL U16528 ( .A(n25716), .B(n12204), .Y(n25699) );
  NAND2XL U16529 ( .A(n12075), .B(n12080), .Y(n12076) );
  INVXL U16530 ( .A(n12078), .Y(n12075) );
  AOI21X1 U16531 ( .A0(n6904), .A1(n12635), .B0(n12634), .Y(n14119) );
  NAND2BXL U16532 ( .AN(n12481), .B(n22689), .Y(n12529) );
  NAND2BXL U16533 ( .AN(n12481), .B(n22688), .Y(n7225) );
  XNOR2X1 U16534 ( .A(n12470), .B(n12469), .Y(n22885) );
  AOI21XL U16535 ( .A0(n22506), .A1(n14044), .B0(n14043), .Y(n14045) );
  OAI21XL U16536 ( .A0(n22522), .A1(n14037), .B0(n14036), .Y(n14038) );
  NAND2XL U16537 ( .A(n22526), .B(n14029), .Y(n14037) );
  NOR2X1 U16538 ( .A(n14031), .B(U2_A_i_d[10]), .Y(n22535) );
  OAI21XL U16539 ( .A0(n13312), .A1(n13308), .B0(n13309), .Y(n13307) );
  XOR2X1 U16540 ( .A(n13312), .B(n13311), .Y(n14024) );
  INVXL U16541 ( .A(n13308), .Y(n13310) );
  XOR2X1 U16542 ( .A(n8820), .B(n8819), .Y(n24583) );
  INVXL U16543 ( .A(n20139), .Y(n19971) );
  NOR2X1 U16544 ( .A(n19980), .B(n19979), .Y(n20121) );
  NAND2XL U16545 ( .A(n6991), .B(n9577), .Y(n9583) );
  AOI21XL U16546 ( .A0(n6991), .A1(n17235), .B0(n9581), .Y(n9582) );
  INVXL U16547 ( .A(n17262), .Y(n9574) );
  NAND2X1 U16548 ( .A(n17229), .B(n6996), .Y(n17211) );
  NAND2XL U16549 ( .A(n7001), .B(n17208), .Y(n13722) );
  AOI21XL U16550 ( .A0(n13728), .A1(n9594), .B0(n9593), .Y(n9595) );
  NOR2X1 U16551 ( .A(n9590), .B(n17211), .Y(n13721) );
  OAI21XL U16552 ( .A0(n13544), .A1(n17403), .B0(n13543), .Y(n17372) );
  NOR2XL U16553 ( .A(n14935), .B(n19321), .Y(n17388) );
  NOR2X1 U16554 ( .A(n13555), .B(n7518), .Y(n17350) );
  NOR2BX1 U16555 ( .AN(n17362), .B(n7519), .Y(n7518) );
  INVX1 U16556 ( .A(n13562), .Y(n7554) );
  NOR2X1 U16557 ( .A(n7502), .B(n17334), .Y(n7501) );
  INVXL U16558 ( .A(n17300), .Y(n7494) );
  INVXL U16559 ( .A(n13872), .Y(n13858) );
  NOR2X1 U16560 ( .A(n19979), .B(n14926), .Y(n20405) );
  NOR2X1 U16561 ( .A(n20390), .B(n14880), .Y(n14882) );
  NAND2XL U16562 ( .A(n20072), .B(n20356), .Y(n20309) );
  NOR2X1 U16563 ( .A(n20317), .B(n20309), .Y(n20318) );
  NOR2XL U16564 ( .A(n13669), .B(U1_A_i_d0[2]), .Y(n17288) );
  INVXL U16565 ( .A(n17242), .Y(n17256) );
  NOR2X1 U16566 ( .A(n13683), .B(U1_A_i_d0[10]), .Y(n17245) );
  OAI21XL U16567 ( .A0(n9452), .A1(n17542), .B0(n9451), .Y(n9453) );
  NAND2X1 U16568 ( .A(n7007), .B(n17530), .Y(n9458) );
  INVX1 U16569 ( .A(n13692), .Y(n9501) );
  AOI21XL U16570 ( .A0(n17700), .A1(n12795), .B0(n12887), .Y(n12888) );
  INVXL U16571 ( .A(n17702), .Y(n12887) );
  INVXL U16572 ( .A(n13632), .Y(n13619) );
  NAND2XL U16573 ( .A(n14968), .B(n19237), .Y(n17300) );
  NAND2XL U16574 ( .A(n19737), .B(U1_A_r_d0[8]), .Y(n19886) );
  AOI2BB1X2 U16575 ( .A0N(n13912), .A1N(n17103), .B0(n7515), .Y(n17084) );
  NAND2XL U16576 ( .A(n13987), .B(n7509), .Y(n7508) );
  INVXL U16577 ( .A(n16790), .Y(n7509) );
  INVXL U16578 ( .A(n12288), .Y(n19711) );
  OAI21XL U16579 ( .A0(n8655), .A1(n16736), .B0(n8654), .Y(n16702) );
  NAND2X1 U16580 ( .A(n6907), .B(n16669), .Y(n16658) );
  AOI21XL U16581 ( .A0(n6907), .A1(n6675), .B0(n7019), .Y(n16657) );
  AND2XL U16582 ( .A(n7543), .B(U1_A_i_d0[18]), .Y(n7019) );
  NAND2XL U16583 ( .A(n14942), .B(n16860), .Y(n14943) );
  INVXL U16584 ( .A(n16892), .Y(n14924) );
  NOR2X1 U16585 ( .A(n16800), .B(n14965), .Y(n16793) );
  INVXL U16586 ( .A(n13626), .Y(n13612) );
  INVXL U16587 ( .A(n13976), .Y(n13973) );
  INVXL U16588 ( .A(n13990), .Y(n13986) );
  INVXL U16589 ( .A(n13653), .Y(n13642) );
  NAND2X1 U16590 ( .A(n16793), .B(n14967), .Y(n16788) );
  OR2XL U16591 ( .A(n19724), .B(n7063), .Y(n19918) );
  OR2X2 U16592 ( .A(n19738), .B(n7065), .Y(n19893) );
  AOI21XL U16593 ( .A0(n12310), .A1(n20245), .B0(n12312), .Y(n20233) );
  NAND2XL U16594 ( .A(n19839), .B(n19843), .Y(n20211) );
  AOI21XL U16595 ( .A0(n19829), .A1(n12321), .B0(n12320), .Y(n12322) );
  NOR2XL U16596 ( .A(n13669), .B(U1_A_r_d0[2]), .Y(n19221) );
  INVX1 U16597 ( .A(n13675), .Y(n9665) );
  OAI21XL U16598 ( .A0(n9672), .A1(n19186), .B0(n9671), .Y(n19152) );
  AND2XL U16599 ( .A(n7627), .B(U1_A_r_d0[14]), .Y(n9691) );
  NOR2XL U16600 ( .A(n19330), .B(n14783), .Y(n19316) );
  NAND2X1 U16601 ( .A(n19304), .B(n19306), .Y(n14792) );
  NOR2X1 U16602 ( .A(n19302), .B(n14792), .Y(n7846) );
  OAI2BB1XL U16603 ( .A0N(n19306), .A1N(n8146), .B0(n19305), .Y(n7845) );
  NAND2X1 U16604 ( .A(n14757), .B(n7850), .Y(n19301) );
  NAND3BXL U16605 ( .AN(n19334), .B(n19336), .C(n19338), .Y(n7850) );
  INVXL U16606 ( .A(n19337), .Y(n14756) );
  INVXL U16607 ( .A(n14841), .Y(n14843) );
  NOR2XL U16608 ( .A(n14851), .B(n19557), .Y(n19251) );
  AOI21X1 U16609 ( .A0(n6985), .A1(n19258), .B0(n6899), .Y(n14836) );
  AND2XL U16610 ( .A(n19259), .B(n5857), .Y(n6899) );
  NAND2X1 U16611 ( .A(n6985), .B(n19263), .Y(n14837) );
  XOR2X1 U16612 ( .A(n8472), .B(n8471), .Y(n12295) );
  INVXL U16613 ( .A(n8468), .Y(n8470) );
  OR2X2 U16614 ( .A(n19738), .B(n7064), .Y(n16723) );
  INVXL U16615 ( .A(n8548), .Y(n8550) );
  NAND2X1 U16616 ( .A(n16708), .B(n8553), .Y(n8559) );
  AOI21XL U16617 ( .A0(n16708), .A1(n16997), .B0(n8557), .Y(n8558) );
  AOI21XL U16618 ( .A0(n8580), .A1(n16987), .B0(n8605), .Y(n16976) );
  NAND2X1 U16619 ( .A(n6906), .B(n16665), .Y(n8614) );
  XOR2X1 U16620 ( .A(n12773), .B(n12772), .Y(n14921) );
  INVXL U16621 ( .A(n12777), .Y(n12771) );
  INVXL U16622 ( .A(n12780), .Y(n12706) );
  OAI21XL U16623 ( .A0(n13846), .A1(n17131), .B0(n13845), .Y(n17107) );
  NAND2XL U16624 ( .A(n7431), .B(n7681), .Y(n9358) );
  NOR2X1 U16625 ( .A(n13683), .B(U1_A_r_d0[10]), .Y(n19172) );
  NAND2X1 U16626 ( .A(n19158), .B(n13680), .Y(n13690) );
  NAND2XL U16627 ( .A(n7024), .B(n19444), .Y(n19431) );
  AOI21XL U16628 ( .A0(n19134), .A1(n13695), .B0(n7688), .Y(n13696) );
  AOI21X1 U16629 ( .A0(n19118), .A1(n13701), .B0(n13700), .Y(n19411) );
  INVXL U16630 ( .A(n14696), .Y(n14698) );
  NOR2X1 U16631 ( .A(n19243), .B(n20041), .Y(n19562) );
  NOR2XL U16632 ( .A(n11957), .B(n28642), .Y(n28663) );
  NOR2XL U16633 ( .A(n11958), .B(n28639), .Y(n28650) );
  NOR2XL U16634 ( .A(n11957), .B(n28637), .Y(n28645) );
  NOR2XL U16635 ( .A(n11957), .B(n28636), .Y(n28648) );
  NOR2XL U16636 ( .A(ram_sel_reg[1]), .B(n11633), .Y(n11986) );
  OAI2BB1XL U16637 ( .A0N(n7305), .A1N(ram_sel_reg[0]), .B0(n11985), .Y(n11982) );
  NAND2XL U16638 ( .A(CQ0[8]), .B(n28921), .Y(n27847) );
  INVXL U16639 ( .A(n27847), .Y(n27848) );
  INVXL U16640 ( .A(n28040), .Y(n28042) );
  NAND2XL U16641 ( .A(CQ0[49]), .B(n28921), .Y(n28040) );
  NAND2XL U16642 ( .A(CQ0[47]), .B(n28921), .Y(n28030) );
  NAND2XL U16643 ( .A(n28921), .B(n28030), .Y(n28031) );
  INVXL U16644 ( .A(n28030), .Y(n28032) );
  NAND2XL U16645 ( .A(CQ0[42]), .B(n28921), .Y(n28005) );
  NAND2XL U16646 ( .A(n28921), .B(n28005), .Y(n28006) );
  INVXL U16647 ( .A(n28005), .Y(n28007) );
  NAND2XL U16648 ( .A(CQ0[38]), .B(n28921), .Y(n27985) );
  NAND2XL U16649 ( .A(n28921), .B(n27985), .Y(n27986) );
  INVXL U16650 ( .A(n27985), .Y(n27987) );
  NAND2XL U16651 ( .A(CQ0[37]), .B(n28921), .Y(n27980) );
  NAND2XL U16652 ( .A(n28921), .B(n27980), .Y(n27981) );
  INVXL U16653 ( .A(n27980), .Y(n27982) );
  NAND2XL U16654 ( .A(CQ0[33]), .B(n28921), .Y(n27963) );
  INVXL U16655 ( .A(n27963), .Y(n27964) );
  NAND2XL U16656 ( .A(CQ0[28]), .B(n28921), .Y(n27942) );
  NAND2XL U16657 ( .A(CQ0[26]), .B(n28921), .Y(n27934) );
  INVXL U16658 ( .A(n27934), .Y(n27935) );
  NAND2XL U16659 ( .A(CQ0[23]), .B(n28921), .Y(n27919) );
  INVXL U16660 ( .A(n27919), .Y(n27921) );
  NAND2XL U16661 ( .A(CQ0[20]), .B(n28921), .Y(n27904) );
  INVXL U16662 ( .A(n27904), .Y(n27906) );
  NAND2XL U16663 ( .A(CQ0[15]), .B(n28921), .Y(n27879) );
  NAND2XL U16664 ( .A(n28921), .B(n27879), .Y(n27880) );
  INVXL U16665 ( .A(n27879), .Y(n27881) );
  NAND2XL U16666 ( .A(CQ0[13]), .B(n28921), .Y(n27869) );
  NAND2XL U16667 ( .A(n28921), .B(n27869), .Y(n27870) );
  INVXL U16668 ( .A(n27869), .Y(n27871) );
  NOR2XL U16669 ( .A(n11896), .B(n28659), .Y(n28669) );
  INVXL U16670 ( .A(n11973), .Y(n11959) );
  INVXL U16671 ( .A(n11640), .Y(n11641) );
  NOR2XL U16672 ( .A(n7863), .B(n20026), .Y(n7937) );
  NOR2X1 U16673 ( .A(n24703), .B(n24690), .Y(n24691) );
  NOR2X1 U16674 ( .A(n24688), .B(n24687), .Y(n24690) );
  NAND2XL U16675 ( .A(n14974), .B(n29008), .Y(n7646) );
  AND2X1 U16676 ( .A(n9548), .B(n9547), .Y(n7653) );
  NOR2XL U16677 ( .A(n14974), .B(n29008), .Y(n7652) );
  INVXL U16678 ( .A(n17462), .Y(n17463) );
  NOR2X1 U16679 ( .A(n13709), .B(U1_A_i_d0[21]), .Y(n17189) );
  NAND2XL U16680 ( .A(n17195), .B(n17191), .Y(n17182) );
  NAND2XL U16681 ( .A(cnt[4]), .B(n11961), .Y(n11969) );
  NOR2XL U16682 ( .A(n28673), .B(n11969), .Y(n11640) );
  INVXL U16683 ( .A(n28630), .Y(n11966) );
  NAND2XL U16684 ( .A(n28705), .B(n28679), .Y(n11965) );
  INVXL U16685 ( .A(n11961), .Y(n11967) );
  NAND2XL U16686 ( .A(n26975), .B(n26974), .Y(n27013) );
  AOI21XL U16687 ( .A0(n26932), .A1(n26891), .B0(n26931), .Y(n26972) );
  INVXL U16688 ( .A(n26930), .Y(n26931) );
  NOR2XL U16689 ( .A(n26934), .B(n26933), .Y(n26971) );
  NAND2XL U16690 ( .A(n26934), .B(n26933), .Y(n26970) );
  NAND2XL U16691 ( .A(n26893), .B(n26892), .Y(n26930) );
  AOI21XL U16692 ( .A0(n26845), .A1(n26798), .B0(n26844), .Y(n26890) );
  INVXL U16693 ( .A(n26843), .Y(n26844) );
  NOR2XL U16694 ( .A(n26847), .B(n26846), .Y(n26889) );
  NAND2XL U16695 ( .A(n26847), .B(n26846), .Y(n26888) );
  INVXL U16696 ( .A(n26734), .Y(n26679) );
  INVXL U16697 ( .A(n26731), .Y(n26680) );
  INVXL U16698 ( .A(n26733), .Y(n26683) );
  NOR2XL U16699 ( .A(n26626), .B(n26629), .Y(n26675) );
  NAND2XL U16700 ( .A(n26632), .B(n26631), .Y(n26676) );
  INVXL U16701 ( .A(n26628), .Y(n26563) );
  NAND2XL U16702 ( .A(n26566), .B(n26565), .Y(n26627) );
  INVXL U16703 ( .A(n26629), .Y(n26567) );
  NAND2XL U16704 ( .A(n26500), .B(n26499), .Y(n26628) );
  INVXL U16705 ( .A(n26626), .Y(n26564) );
  INVXL U16706 ( .A(n26488), .Y(n26433) );
  NAND2XL U16707 ( .A(n26437), .B(n26436), .Y(n26487) );
  INVXL U16708 ( .A(n26489), .Y(n26438) );
  NAND2XL U16709 ( .A(n26388), .B(n26387), .Y(n26488) );
  INVXL U16710 ( .A(n26485), .Y(n26385) );
  INVXL U16711 ( .A(n26491), .Y(n26384) );
  INVXL U16712 ( .A(n26484), .Y(n26434) );
  INVXL U16713 ( .A(n26382), .Y(n26324) );
  NAND2XL U16714 ( .A(n26328), .B(n26327), .Y(n26381) );
  INVXL U16715 ( .A(n26383), .Y(n26329) );
  INVXL U16716 ( .A(n26326), .Y(n26386) );
  NAND2XL U16717 ( .A(n26266), .B(n26265), .Y(n26382) );
  INVXL U16718 ( .A(n26380), .Y(n26325) );
  INVXL U16719 ( .A(n26259), .Y(n26206) );
  NAND2XL U16720 ( .A(n26210), .B(n26209), .Y(n26258) );
  INVXL U16721 ( .A(n26260), .Y(n26211) );
  NAND2XL U16722 ( .A(n26173), .B(n26172), .Y(n26259) );
  INVXL U16723 ( .A(n26257), .Y(n26171) );
  INVXL U16724 ( .A(n26262), .Y(n26170) );
  INVXL U16725 ( .A(n26256), .Y(n26207) );
  INVXL U16726 ( .A(n26444), .Y(n26391) );
  INVXL U16727 ( .A(n26445), .Y(n26396) );
  INVXL U16728 ( .A(n26442), .Y(n26392) );
  INVXL U16729 ( .A(n26314), .Y(n26278) );
  NAND2XL U16730 ( .A(n26282), .B(n26281), .Y(n26313) );
  INVXL U16731 ( .A(n26315), .Y(n26283) );
  NAND2XL U16732 ( .A(n26232), .B(n26231), .Y(n26314) );
  INVXL U16733 ( .A(n26312), .Y(n26230) );
  INVXL U16734 ( .A(n26317), .Y(n26229) );
  INVXL U16735 ( .A(n26311), .Y(n26279) );
  INVXL U16736 ( .A(n25995), .Y(n25975) );
  NAND2XL U16737 ( .A(n25978), .B(n25977), .Y(n25994) );
  INVXL U16738 ( .A(n25996), .Y(n25979) );
  NAND2XL U16739 ( .A(n25933), .B(n25932), .Y(n25995) );
  INVXL U16740 ( .A(n26136), .Y(n25997) );
  INVXL U16741 ( .A(n25993), .Y(n25976) );
  NAND2XL U16742 ( .A(n24308), .B(n24307), .Y(n24346) );
  AOI21XL U16743 ( .A0(n24280), .A1(n24239), .B0(n24279), .Y(n24305) );
  INVXL U16744 ( .A(n24278), .Y(n24279) );
  NOR2XL U16745 ( .A(n24282), .B(n24281), .Y(n24304) );
  NAND2XL U16746 ( .A(n24282), .B(n24281), .Y(n24303) );
  NAND2XL U16747 ( .A(n24241), .B(n24240), .Y(n24278) );
  NOR2XL U16748 ( .A(n24195), .B(n24194), .Y(n24237) );
  NAND2XL U16749 ( .A(n24195), .B(n24194), .Y(n24236) );
  NAND2XL U16750 ( .A(n24126), .B(n24125), .Y(n24191) );
  NAND2XL U16751 ( .A(n24117), .B(n24085), .Y(n24122) );
  AOI21XL U16752 ( .A0(n24120), .A1(n24085), .B0(n24119), .Y(n24121) );
  INVXL U16753 ( .A(n24118), .Y(n24119) );
  INVXL U16754 ( .A(n24083), .Y(n24004) );
  INVXL U16755 ( .A(n24080), .Y(n24005) );
  INVXL U16756 ( .A(n24082), .Y(n24008) );
  NOR2XL U16757 ( .A(n23969), .B(n23972), .Y(n24000) );
  NAND2XL U16758 ( .A(n23975), .B(n23974), .Y(n24001) );
  INVXL U16759 ( .A(n23971), .Y(n23914) );
  NAND2XL U16760 ( .A(n23917), .B(n23916), .Y(n23970) );
  INVXL U16761 ( .A(n23972), .Y(n23918) );
  NAND2XL U16762 ( .A(n23826), .B(n23825), .Y(n23971) );
  INVXL U16763 ( .A(n23969), .Y(n23915) );
  INVXL U16764 ( .A(n23814), .Y(n23761) );
  NAND2XL U16765 ( .A(n23765), .B(n23764), .Y(n23813) );
  INVXL U16766 ( .A(n23815), .Y(n23766) );
  NAND2XL U16767 ( .A(n23736), .B(n23735), .Y(n23814) );
  INVXL U16768 ( .A(n23811), .Y(n23733) );
  INVXL U16769 ( .A(n23817), .Y(n23732) );
  INVXL U16770 ( .A(n23810), .Y(n23762) );
  INVXL U16771 ( .A(n23656), .Y(n23734) );
  INVXL U16772 ( .A(n23585), .Y(n23561) );
  NAND2XL U16773 ( .A(n23565), .B(n23564), .Y(n23584) );
  INVXL U16774 ( .A(n23586), .Y(n23566) );
  NAND2XL U16775 ( .A(n23521), .B(n23520), .Y(n23585) );
  INVXL U16776 ( .A(n23583), .Y(n23519) );
  INVXL U16777 ( .A(n23588), .Y(n23518) );
  INVXL U16778 ( .A(n23582), .Y(n23562) );
  NAND2XL U16779 ( .A(n26983), .B(n26982), .Y(n27021) );
  NAND2XL U16780 ( .A(n26885), .B(n26884), .Y(n26922) );
  NOR2XL U16781 ( .A(n26839), .B(n26838), .Y(n26881) );
  NAND2XL U16782 ( .A(n26839), .B(n26838), .Y(n26880) );
  NAND2XL U16783 ( .A(n26788), .B(n26787), .Y(n26835) );
  NAND2XL U16784 ( .A(n26779), .B(n26747), .Y(n26784) );
  AOI21XL U16785 ( .A0(n26782), .A1(n26747), .B0(n26781), .Y(n26783) );
  INVXL U16786 ( .A(n26780), .Y(n26781) );
  NOR2XL U16787 ( .A(n26742), .B(n26744), .Y(n26779) );
  NAND2XL U16788 ( .A(n26749), .B(n26748), .Y(n26780) );
  INVXL U16789 ( .A(n26742), .Y(n26668) );
  INVXL U16790 ( .A(n26745), .Y(n26667) );
  NAND2XL U16791 ( .A(n26670), .B(n26669), .Y(n26743) );
  INVXL U16792 ( .A(n26744), .Y(n26671) );
  INVXL U16793 ( .A(n26619), .Y(n26666) );
  NAND2XL U16794 ( .A(n26622), .B(n26621), .Y(n26664) );
  NAND2XL U16795 ( .A(n26588), .B(n26587), .Y(n26619) );
  INVXL U16796 ( .A(n26575), .Y(n26503) );
  NAND2XL U16797 ( .A(n26507), .B(n26506), .Y(n26574) );
  INVXL U16798 ( .A(n26576), .Y(n26508) );
  NAND2XL U16799 ( .A(n26430), .B(n26429), .Y(n26575) );
  INVXL U16800 ( .A(n26572), .Y(n26427) );
  INVXL U16801 ( .A(n26578), .Y(n26426) );
  INVXL U16802 ( .A(n26571), .Y(n26504) );
  INVXL U16803 ( .A(n26424), .Y(n26371) );
  NAND2XL U16804 ( .A(n26375), .B(n26374), .Y(n26423) );
  INVXL U16805 ( .A(n26425), .Y(n26376) );
  INVXL U16806 ( .A(n26373), .Y(n26428) );
  NAND2XL U16807 ( .A(n26343), .B(n26342), .Y(n26424) );
  INVXL U16808 ( .A(n26422), .Y(n26372) );
  INVXL U16809 ( .A(n26336), .Y(n26247) );
  NAND2XL U16810 ( .A(n26251), .B(n26250), .Y(n26335) );
  INVXL U16811 ( .A(n26337), .Y(n26252) );
  NAND2XL U16812 ( .A(n26203), .B(n26202), .Y(n26336) );
  INVXL U16813 ( .A(n26339), .Y(n26200) );
  INVXL U16814 ( .A(n26334), .Y(n26201) );
  INVXL U16815 ( .A(n26333), .Y(n26248) );
  INVXL U16816 ( .A(n26022), .Y(n25949) );
  NAND2XL U16817 ( .A(n25952), .B(n25951), .Y(n26021) );
  INVXL U16818 ( .A(n26023), .Y(n25953) );
  NAND2XL U16819 ( .A(n25903), .B(n25902), .Y(n26022) );
  INVXL U16820 ( .A(n26098), .Y(n26024) );
  INVXL U16821 ( .A(n26020), .Y(n25950) );
  AOI21XL U16822 ( .A0(n25796), .A1(n25795), .B0(n25794), .Y(n25831) );
  OR2XL U16823 ( .A(U0_pipe9[1]), .B(U0_pipe8[1]), .Y(n25796) );
  AND2XL U16824 ( .A(U0_pipe9[1]), .B(U0_pipe8[1]), .Y(n25794) );
  NOR2XL U16825 ( .A(n25792), .B(n28896), .Y(n25830) );
  NAND2XL U16826 ( .A(n25792), .B(n28896), .Y(n25829) );
  NAND2XL U16827 ( .A(n24316), .B(n24315), .Y(n24354) );
  AOI21XL U16828 ( .A0(n24272), .A1(n24231), .B0(n24271), .Y(n24313) );
  INVXL U16829 ( .A(n24270), .Y(n24271) );
  NOR2XL U16830 ( .A(n24274), .B(n24273), .Y(n24312) );
  NAND2XL U16831 ( .A(n24274), .B(n24273), .Y(n24311) );
  NAND2XL U16832 ( .A(n24233), .B(n24232), .Y(n24270) );
  NOR2XL U16833 ( .A(n24187), .B(n24186), .Y(n24229) );
  NAND2XL U16834 ( .A(n24187), .B(n24186), .Y(n24228) );
  NAND2XL U16835 ( .A(n24139), .B(n24138), .Y(n24183) );
  NAND2XL U16836 ( .A(n24130), .B(n24074), .Y(n24135) );
  AOI21XL U16837 ( .A0(n24133), .A1(n24074), .B0(n24132), .Y(n24134) );
  INVXL U16838 ( .A(n24131), .Y(n24132) );
  INVXL U16839 ( .A(n24072), .Y(n24016) );
  INVXL U16840 ( .A(n24069), .Y(n24017) );
  INVXL U16841 ( .A(n24071), .Y(n24020) );
  NOR2XL U16842 ( .A(n23959), .B(n23962), .Y(n24012) );
  NAND2XL U16843 ( .A(n23965), .B(n23964), .Y(n24013) );
  INVXL U16844 ( .A(n23961), .Y(n23906) );
  NAND2XL U16845 ( .A(n23909), .B(n23908), .Y(n23960) );
  INVXL U16846 ( .A(n23962), .Y(n23910) );
  NAND2XL U16847 ( .A(n23845), .B(n23844), .Y(n23961) );
  INVXL U16848 ( .A(n23959), .Y(n23907) );
  INVXL U16849 ( .A(n23833), .Y(n23770) );
  NAND2XL U16850 ( .A(n23774), .B(n23773), .Y(n23832) );
  INVXL U16851 ( .A(n23834), .Y(n23775) );
  NAND2XL U16852 ( .A(n23725), .B(n23724), .Y(n23833) );
  INVXL U16853 ( .A(n23830), .Y(n23722) );
  INVXL U16854 ( .A(n23836), .Y(n23721) );
  INVXL U16855 ( .A(n23829), .Y(n23771) );
  INVXL U16856 ( .A(n23665), .Y(n23723) );
  INVXL U16857 ( .A(n23598), .Y(n23541) );
  NAND2XL U16858 ( .A(n23545), .B(n23544), .Y(n23597) );
  INVXL U16859 ( .A(n23599), .Y(n23546) );
  NAND2XL U16860 ( .A(n23505), .B(n23504), .Y(n23598) );
  INVXL U16861 ( .A(n23596), .Y(n23503) );
  INVXL U16862 ( .A(n23601), .Y(n23502) );
  INVXL U16863 ( .A(n23595), .Y(n23542) );
  NAND2XL U16864 ( .A(n24300), .B(n24299), .Y(n24338) );
  AOI21XL U16865 ( .A0(n24256), .A1(n24215), .B0(n24255), .Y(n24297) );
  INVXL U16866 ( .A(n24254), .Y(n24255) );
  NOR2XL U16867 ( .A(n24258), .B(n24257), .Y(n24296) );
  NAND2XL U16868 ( .A(n24258), .B(n24257), .Y(n24295) );
  NAND2XL U16869 ( .A(n24217), .B(n24216), .Y(n24254) );
  NOR2XL U16870 ( .A(n24171), .B(n24170), .Y(n24213) );
  NAND2XL U16871 ( .A(n24171), .B(n24170), .Y(n24212) );
  NAND2XL U16872 ( .A(n24114), .B(n24113), .Y(n24167) );
  NAND2XL U16873 ( .A(n24105), .B(n24052), .Y(n24110) );
  AOI21XL U16874 ( .A0(n24108), .A1(n24052), .B0(n24107), .Y(n24109) );
  INVXL U16875 ( .A(n24106), .Y(n24107) );
  NOR2XL U16876 ( .A(n24047), .B(n24049), .Y(n24105) );
  NAND2XL U16877 ( .A(n24054), .B(n24053), .Y(n24106) );
  INVXL U16878 ( .A(n24047), .Y(n23993) );
  INVXL U16879 ( .A(n24050), .Y(n23992) );
  NAND2XL U16880 ( .A(n23995), .B(n23994), .Y(n24048) );
  INVXL U16881 ( .A(n24049), .Y(n23996) );
  INVXL U16882 ( .A(n23882), .Y(n23801) );
  NAND2XL U16883 ( .A(n23805), .B(n23804), .Y(n23881) );
  INVXL U16884 ( .A(n23883), .Y(n23806) );
  NAND2XL U16885 ( .A(n23758), .B(n23757), .Y(n23882) );
  INVXL U16886 ( .A(n23879), .Y(n23755) );
  INVXL U16887 ( .A(n23885), .Y(n23754) );
  INVXL U16888 ( .A(n23878), .Y(n23802) );
  INVXL U16889 ( .A(n23752), .Y(n23697) );
  NAND2XL U16890 ( .A(n23701), .B(n23700), .Y(n23751) );
  INVXL U16891 ( .A(n23753), .Y(n23702) );
  INVXL U16892 ( .A(n23699), .Y(n23756) );
  NAND2XL U16893 ( .A(n23651), .B(n23650), .Y(n23752) );
  INVXL U16894 ( .A(n23750), .Y(n23698) );
  INVXL U16895 ( .A(n23644), .Y(n23608) );
  NAND2XL U16896 ( .A(n23612), .B(n23611), .Y(n23643) );
  INVXL U16897 ( .A(n23645), .Y(n23613) );
  NAND2XL U16898 ( .A(n23557), .B(n23556), .Y(n23644) );
  INVXL U16899 ( .A(n23642), .Y(n23555) );
  INVXL U16900 ( .A(n23647), .Y(n23554) );
  INVXL U16901 ( .A(n23641), .Y(n23609) );
  INVXL U16902 ( .A(n23345), .Y(n23301) );
  NAND2XL U16903 ( .A(n23304), .B(n23303), .Y(n23344) );
  INVXL U16904 ( .A(n23346), .Y(n23305) );
  NAND2XL U16905 ( .A(n23257), .B(n23256), .Y(n23345) );
  INVXL U16906 ( .A(n23458), .Y(n23347) );
  INVXL U16907 ( .A(n23343), .Y(n23302) );
  NAND2XL U16908 ( .A(n26959), .B(n26958), .Y(n26997) );
  AOI21XL U16909 ( .A0(n26916), .A1(n26875), .B0(n26915), .Y(n26956) );
  INVXL U16910 ( .A(n26914), .Y(n26915) );
  NOR2XL U16911 ( .A(n26918), .B(n26917), .Y(n26955) );
  NAND2XL U16912 ( .A(n26918), .B(n26917), .Y(n26954) );
  NAND2XL U16913 ( .A(n26877), .B(n26876), .Y(n26914) );
  NOR2XL U16914 ( .A(n26831), .B(n26830), .Y(n26873) );
  NAND2XL U16915 ( .A(n26831), .B(n26830), .Y(n26872) );
  NAND2XL U16916 ( .A(n26776), .B(n26775), .Y(n26827) );
  NAND2XL U16917 ( .A(n26767), .B(n26714), .Y(n26772) );
  INVXL U16918 ( .A(n26768), .Y(n26769) );
  NOR2XL U16919 ( .A(n26709), .B(n26711), .Y(n26767) );
  NAND2XL U16920 ( .A(n26716), .B(n26715), .Y(n26768) );
  INVXL U16921 ( .A(n26709), .Y(n26657) );
  INVXL U16922 ( .A(n26712), .Y(n26656) );
  NAND2XL U16923 ( .A(n26659), .B(n26658), .Y(n26710) );
  INVXL U16924 ( .A(n26711), .Y(n26660) );
  INVXL U16925 ( .A(n26612), .Y(n26655) );
  NAND2XL U16926 ( .A(n26615), .B(n26614), .Y(n26653) );
  NAND2XL U16927 ( .A(n26540), .B(n26539), .Y(n26612) );
  INVXL U16928 ( .A(n26527), .Y(n26466) );
  NAND2XL U16929 ( .A(n26470), .B(n26469), .Y(n26526) );
  INVXL U16930 ( .A(n26528), .Y(n26471) );
  NAND2XL U16931 ( .A(n26419), .B(n26418), .Y(n26527) );
  INVXL U16932 ( .A(n26524), .Y(n26416) );
  INVXL U16933 ( .A(n26530), .Y(n26415) );
  INVXL U16934 ( .A(n26523), .Y(n26467) );
  INVXL U16935 ( .A(n26413), .Y(n26362) );
  NAND2XL U16936 ( .A(n26366), .B(n26365), .Y(n26412) );
  INVXL U16937 ( .A(n26414), .Y(n26367) );
  INVXL U16938 ( .A(n26301), .Y(n26269) );
  NAND2XL U16939 ( .A(n26273), .B(n26272), .Y(n26300) );
  INVXL U16940 ( .A(n26302), .Y(n26274) );
  NAND2XL U16941 ( .A(n26222), .B(n26221), .Y(n26301) );
  INVXL U16942 ( .A(n26299), .Y(n26220) );
  INVXL U16943 ( .A(n26304), .Y(n26219) );
  INVXL U16944 ( .A(n26298), .Y(n26270) );
  INVXL U16945 ( .A(n26012), .Y(n25967) );
  NAND2XL U16946 ( .A(n25970), .B(n25969), .Y(n26011) );
  INVXL U16947 ( .A(n26013), .Y(n25971) );
  NAND2XL U16948 ( .A(n25922), .B(n25921), .Y(n26012) );
  INVXL U16949 ( .A(n26120), .Y(n26014) );
  INVXL U16950 ( .A(n26010), .Y(n25968) );
  NAND2XL U16951 ( .A(n24324), .B(n24323), .Y(n24362) );
  AOI21XL U16952 ( .A0(n24264), .A1(n24223), .B0(n24263), .Y(n24321) );
  INVXL U16953 ( .A(n24262), .Y(n24263) );
  NOR2XL U16954 ( .A(n24266), .B(n24265), .Y(n24320) );
  NAND2XL U16955 ( .A(n24266), .B(n24265), .Y(n24319) );
  NAND2XL U16956 ( .A(n24225), .B(n24224), .Y(n24262) );
  NOR2XL U16957 ( .A(n24179), .B(n24178), .Y(n24221) );
  NAND2XL U16958 ( .A(n24179), .B(n24178), .Y(n24220) );
  NAND2XL U16959 ( .A(n24151), .B(n24150), .Y(n24175) );
  NAND2XL U16960 ( .A(n24142), .B(n24063), .Y(n24147) );
  AOI21XL U16961 ( .A0(n24145), .A1(n24063), .B0(n24144), .Y(n24146) );
  INVXL U16962 ( .A(n24143), .Y(n24144) );
  NOR2XL U16963 ( .A(n24058), .B(n24060), .Y(n24142) );
  NAND2XL U16964 ( .A(n24065), .B(n24064), .Y(n24143) );
  INVXL U16965 ( .A(n24061), .Y(n24028) );
  INVXL U16966 ( .A(n24058), .Y(n24029) );
  NAND2XL U16967 ( .A(n24031), .B(n24030), .Y(n24059) );
  INVXL U16968 ( .A(n24060), .Y(n24032) );
  NOR2XL U16969 ( .A(n23949), .B(n23952), .Y(n24024) );
  NAND2XL U16970 ( .A(n23955), .B(n23954), .Y(n24025) );
  INVXL U16971 ( .A(n23951), .Y(n23898) );
  NAND2XL U16972 ( .A(n23901), .B(n23900), .Y(n23950) );
  INVXL U16973 ( .A(n23952), .Y(n23902) );
  INVXL U16974 ( .A(n23852), .Y(n23779) );
  NAND2XL U16975 ( .A(n23783), .B(n23782), .Y(n23851) );
  INVXL U16976 ( .A(n23853), .Y(n23784) );
  NAND2XL U16977 ( .A(n23714), .B(n23713), .Y(n23852) );
  INVXL U16978 ( .A(n23849), .Y(n23711) );
  INVXL U16979 ( .A(n23855), .Y(n23710) );
  INVXL U16980 ( .A(n23848), .Y(n23780) );
  INVXL U16981 ( .A(n23708), .Y(n23672) );
  NAND2XL U16982 ( .A(n23676), .B(n23675), .Y(n23707) );
  INVXL U16983 ( .A(n23709), .Y(n23677) );
  INVXL U16984 ( .A(n23674), .Y(n23712) );
  NAND2XL U16985 ( .A(n23627), .B(n23626), .Y(n23708) );
  INVXL U16986 ( .A(n23706), .Y(n23673) );
  NAND2XL U16987 ( .A(n26967), .B(n26966), .Y(n27005) );
  AOI21XL U16988 ( .A0(n26940), .A1(n26899), .B0(n26939), .Y(n26964) );
  INVXL U16989 ( .A(n26938), .Y(n26939) );
  NOR2XL U16990 ( .A(n26942), .B(n26941), .Y(n26963) );
  NAND2XL U16991 ( .A(n26942), .B(n26941), .Y(n26962) );
  NAND2XL U16992 ( .A(n26901), .B(n26900), .Y(n26938) );
  NOR2XL U16993 ( .A(n26855), .B(n26854), .Y(n26897) );
  NAND2XL U16994 ( .A(n26855), .B(n26854), .Y(n26896) );
  NAND2XL U16995 ( .A(n26812), .B(n26811), .Y(n26851) );
  NAND2XL U16996 ( .A(n26803), .B(n26725), .Y(n26808) );
  AOI21XL U16997 ( .A0(n26806), .A1(n26725), .B0(n26805), .Y(n26807) );
  INVXL U16998 ( .A(n26804), .Y(n26805) );
  NOR2XL U16999 ( .A(n26720), .B(n26722), .Y(n26803) );
  NAND2XL U17000 ( .A(n26727), .B(n26726), .Y(n26804) );
  INVXL U17001 ( .A(n26636), .Y(n26689) );
  NAND2XL U17002 ( .A(n26639), .B(n26638), .Y(n26687) );
  NAND2XL U17003 ( .A(n26560), .B(n26559), .Y(n26636) );
  INVXL U17004 ( .A(n26547), .Y(n26475) );
  NAND2XL U17005 ( .A(n26479), .B(n26478), .Y(n26546) );
  INVXL U17006 ( .A(n26548), .Y(n26480) );
  NAND2XL U17007 ( .A(n26450), .B(n26449), .Y(n26547) );
  INVXL U17008 ( .A(n26544), .Y(n26447) );
  INVXL U17009 ( .A(n26550), .Y(n26446) );
  INVXL U17010 ( .A(n26543), .Y(n26476) );
  NAND2XL U17011 ( .A(n21115), .B(n21114), .Y(n21220) );
  INVXL U17012 ( .A(n21216), .Y(n21167) );
  INVXL U17013 ( .A(n21220), .Y(n21166) );
  NAND2XL U17014 ( .A(n21170), .B(n21169), .Y(n21219) );
  INVXL U17015 ( .A(n21221), .Y(n21171) );
  INVXL U17016 ( .A(n21217), .Y(n21112) );
  INVXL U17017 ( .A(n21223), .Y(n21111) );
  NAND2XL U17018 ( .A(n21233), .B(n21232), .Y(n21297) );
  INVXL U17019 ( .A(n21297), .Y(n21328) );
  NAND2XL U17020 ( .A(n21300), .B(n21299), .Y(n21326) );
  INVXL U17021 ( .A(n21383), .Y(n21329) );
  INVXL U17022 ( .A(n21380), .Y(n21330) );
  INVXL U17023 ( .A(n21382), .Y(n21333) );
  NAND2XL U17024 ( .A(n21450), .B(n21449), .Y(n21510) );
  NAND2XL U17025 ( .A(n21441), .B(n21385), .Y(n21446) );
  AOI21XL U17026 ( .A0(n21444), .A1(n21385), .B0(n21443), .Y(n21445) );
  INVXL U17027 ( .A(n21442), .Y(n21443) );
  AOI21XL U17028 ( .A0(n21512), .A1(n21448), .B0(n21511), .Y(n21562) );
  INVXL U17029 ( .A(n21510), .Y(n21511) );
  NOR2XL U17030 ( .A(n21514), .B(n21513), .Y(n21561) );
  NAND2XL U17031 ( .A(n21514), .B(n21513), .Y(n21560) );
  NAND2XL U17032 ( .A(n21565), .B(n21564), .Y(n21604) );
  AOI21XL U17033 ( .A0(n21606), .A1(n21563), .B0(n21605), .Y(n21632) );
  INVXL U17034 ( .A(n21604), .Y(n21605) );
  NOR2XL U17035 ( .A(n21608), .B(n21607), .Y(n21631) );
  NAND2XL U17036 ( .A(n21608), .B(n21607), .Y(n21630) );
  NAND2XL U17037 ( .A(n21635), .B(n21634), .Y(n21668) );
  NAND2XL U17038 ( .A(n17805), .B(n17804), .Y(n17925) );
  INVXL U17039 ( .A(n17923), .Y(n17851) );
  INVXL U17040 ( .A(n17925), .Y(n17850) );
  NAND2XL U17041 ( .A(n17853), .B(n17852), .Y(n17924) );
  INVXL U17042 ( .A(n17926), .Y(n17854) );
  INVXL U17043 ( .A(n17995), .Y(n17927) );
  NAND2XL U17044 ( .A(n18107), .B(n18106), .Y(n18234) );
  INVXL U17045 ( .A(n18231), .Y(n18149) );
  INVXL U17046 ( .A(n18234), .Y(n18148) );
  NAND2XL U17047 ( .A(n18152), .B(n18151), .Y(n18233) );
  INVXL U17048 ( .A(n18235), .Y(n18153) );
  INVXL U17049 ( .A(n18232), .Y(n18105) );
  INVXL U17050 ( .A(n18237), .Y(n18104) );
  NAND2XL U17051 ( .A(n18327), .B(n18326), .Y(n18428) );
  INVXL U17052 ( .A(n18424), .Y(n18396) );
  INVXL U17053 ( .A(n18428), .Y(n18395) );
  NAND2XL U17054 ( .A(n18399), .B(n18398), .Y(n18427) );
  INVXL U17055 ( .A(n18429), .Y(n18400) );
  INVXL U17056 ( .A(n18425), .Y(n18324) );
  INVXL U17057 ( .A(n18431), .Y(n18323) );
  NAND2XL U17058 ( .A(n18440), .B(n18439), .Y(n18583) );
  INVXL U17059 ( .A(n18581), .Y(n18521) );
  INVXL U17060 ( .A(n18583), .Y(n18520) );
  NAND2XL U17061 ( .A(n18523), .B(n18522), .Y(n18582) );
  INVXL U17062 ( .A(n18584), .Y(n18524) );
  NOR2XL U17063 ( .A(n18581), .B(n18584), .Y(n18613) );
  NAND2XL U17064 ( .A(n18587), .B(n18586), .Y(n18614) );
  INVXL U17065 ( .A(n18692), .Y(n18617) );
  INVXL U17066 ( .A(n18689), .Y(n18618) );
  INVXL U17067 ( .A(n18691), .Y(n18621) );
  NAND2XL U17068 ( .A(n18762), .B(n18761), .Y(n18782) );
  NAND2XL U17069 ( .A(n18753), .B(n18694), .Y(n18758) );
  AOI21XL U17070 ( .A0(n18756), .A1(n18694), .B0(n18755), .Y(n18757) );
  INVXL U17071 ( .A(n18754), .Y(n18755) );
  AOI21XL U17072 ( .A0(n18784), .A1(n18760), .B0(n18783), .Y(n18850) );
  INVXL U17073 ( .A(n18782), .Y(n18783) );
  NOR2XL U17074 ( .A(n18786), .B(n18785), .Y(n18849) );
  NAND2XL U17075 ( .A(n18786), .B(n18785), .Y(n18848) );
  NAND2XL U17076 ( .A(n18853), .B(n18852), .Y(n18895) );
  NAND2XL U17077 ( .A(n18940), .B(n18939), .Y(n18971) );
  AND2XL U17078 ( .A(U1_pipe13[1]), .B(U1_pipe12[1]), .Y(n20183) );
  NOR2XL U17079 ( .A(n20181), .B(n28902), .Y(n20490) );
  NAND2XL U17080 ( .A(n20181), .B(n28902), .Y(n20489) );
  NAND2XL U17081 ( .A(n20587), .B(n20586), .Y(n20676) );
  INVXL U17082 ( .A(n20674), .Y(n20630) );
  INVXL U17083 ( .A(n20676), .Y(n20629) );
  NAND2XL U17084 ( .A(n20632), .B(n20631), .Y(n20675) );
  INVXL U17085 ( .A(n20677), .Y(n20633) );
  INVXL U17086 ( .A(n20790), .Y(n20678) );
  NAND2XL U17087 ( .A(n20886), .B(n20885), .Y(n20968) );
  INVXL U17088 ( .A(n20965), .Y(n20933) );
  INVXL U17089 ( .A(n20968), .Y(n20932) );
  NAND2XL U17090 ( .A(n20936), .B(n20935), .Y(n20967) );
  INVXL U17091 ( .A(n20969), .Y(n20937) );
  INVXL U17092 ( .A(n20966), .Y(n20884) );
  INVXL U17093 ( .A(n20971), .Y(n20883) );
  INVXL U17094 ( .A(n21078), .Y(n21025) );
  INVXL U17095 ( .A(n21079), .Y(n21030) );
  NAND2XL U17096 ( .A(n21084), .B(n21083), .Y(n21200) );
  INVXL U17097 ( .A(n21196), .Y(n21130) );
  INVXL U17098 ( .A(n21200), .Y(n21129) );
  NAND2XL U17099 ( .A(n21133), .B(n21132), .Y(n21199) );
  INVXL U17100 ( .A(n21201), .Y(n21134) );
  INVXL U17101 ( .A(n21197), .Y(n21081) );
  INVXL U17102 ( .A(n21203), .Y(n21080) );
  NAND2XL U17103 ( .A(n21213), .B(n21212), .Y(n21273) );
  INVXL U17104 ( .A(n21273), .Y(n21317) );
  NAND2XL U17105 ( .A(n21276), .B(n21275), .Y(n21315) );
  INVXL U17106 ( .A(n21369), .Y(n21319) );
  INVXL U17107 ( .A(n21372), .Y(n21318) );
  INVXL U17108 ( .A(n21371), .Y(n21322) );
  NAND2XL U17109 ( .A(n21438), .B(n21437), .Y(n21486) );
  NAND2XL U17110 ( .A(n21429), .B(n21374), .Y(n21434) );
  AOI21XL U17111 ( .A0(n21432), .A1(n21374), .B0(n21431), .Y(n21433) );
  INVXL U17112 ( .A(n21430), .Y(n21431) );
  NOR2XL U17113 ( .A(n21490), .B(n21489), .Y(n21537) );
  NAND2XL U17114 ( .A(n21490), .B(n21489), .Y(n21536) );
  INVXL U17115 ( .A(n21580), .Y(n21581) );
  NOR2XL U17116 ( .A(n21584), .B(n21583), .Y(n21623) );
  NAND2XL U17117 ( .A(n21584), .B(n21583), .Y(n21622) );
  NAND2XL U17118 ( .A(n21627), .B(n21626), .Y(n21660) );
  NAND2XL U17119 ( .A(n17874), .B(n17873), .Y(n17961) );
  INVXL U17120 ( .A(n17959), .Y(n17916) );
  INVXL U17121 ( .A(n17961), .Y(n17915) );
  NAND2XL U17122 ( .A(n17918), .B(n17917), .Y(n17960) );
  INVXL U17123 ( .A(n17962), .Y(n17919) );
  INVXL U17124 ( .A(n18080), .Y(n17963) );
  NAND2XL U17125 ( .A(n18173), .B(n18172), .Y(n18262) );
  INVXL U17126 ( .A(n18259), .Y(n18223) );
  INVXL U17127 ( .A(n18262), .Y(n18222) );
  NAND2XL U17128 ( .A(n18226), .B(n18225), .Y(n18261) );
  INVXL U17129 ( .A(n18263), .Y(n18227) );
  INVXL U17130 ( .A(n18260), .Y(n18171) );
  INVXL U17131 ( .A(n18265), .Y(n18170) );
  INVXL U17132 ( .A(n18366), .Y(n18311) );
  INVXL U17133 ( .A(n18368), .Y(n18310) );
  INVXL U17134 ( .A(n18369), .Y(n18315) );
  NAND2XL U17135 ( .A(n18374), .B(n18373), .Y(n18504) );
  INVXL U17136 ( .A(n18500), .Y(n18416) );
  INVXL U17137 ( .A(n18504), .Y(n18415) );
  NAND2XL U17138 ( .A(n18419), .B(n18418), .Y(n18503) );
  INVXL U17139 ( .A(n18505), .Y(n18420) );
  INVXL U17140 ( .A(n18501), .Y(n18371) );
  INVXL U17141 ( .A(n18507), .Y(n18370) );
  INVXL U17142 ( .A(n18554), .Y(n18604) );
  NAND2XL U17143 ( .A(n18557), .B(n18556), .Y(n18602) );
  INVXL U17144 ( .A(n18656), .Y(n18606) );
  INVXL U17145 ( .A(n18659), .Y(n18605) );
  INVXL U17146 ( .A(n18658), .Y(n18609) );
  NAND2XL U17147 ( .A(n18725), .B(n18724), .Y(n18774) );
  NAND2XL U17148 ( .A(n18716), .B(n18661), .Y(n18721) );
  AOI21XL U17149 ( .A0(n18719), .A1(n18661), .B0(n18718), .Y(n18720) );
  INVXL U17150 ( .A(n18717), .Y(n18718) );
  AOI21XL U17151 ( .A0(n18776), .A1(n18723), .B0(n18775), .Y(n18826) );
  INVXL U17152 ( .A(n18774), .Y(n18775) );
  NOR2XL U17153 ( .A(n18778), .B(n18777), .Y(n18825) );
  NAND2XL U17154 ( .A(n18778), .B(n18777), .Y(n18824) );
  NAND2XL U17155 ( .A(n18829), .B(n18828), .Y(n18870) );
  AOI21XL U17156 ( .A0(n18872), .A1(n18827), .B0(n18871), .Y(n18913) );
  INVXL U17157 ( .A(n18870), .Y(n18871) );
  NOR2XL U17158 ( .A(n18874), .B(n18873), .Y(n18912) );
  NAND2XL U17159 ( .A(n18874), .B(n18873), .Y(n18911) );
  NAND2XL U17160 ( .A(n18916), .B(n18915), .Y(n18947) );
  NAND2XL U17161 ( .A(n18117), .B(n18116), .Y(n18212) );
  INVXL U17162 ( .A(n18209), .Y(n18158) );
  INVXL U17163 ( .A(n18212), .Y(n18157) );
  NAND2XL U17164 ( .A(n18161), .B(n18160), .Y(n18211) );
  INVXL U17165 ( .A(n18213), .Y(n18162) );
  INVXL U17166 ( .A(n18210), .Y(n18115) );
  INVXL U17167 ( .A(n18215), .Y(n18114) );
  NAND2XL U17168 ( .A(n18219), .B(n18218), .Y(n18332) );
  INVXL U17169 ( .A(n18330), .Y(n18282) );
  INVXL U17170 ( .A(n18332), .Y(n18281) );
  NAND2XL U17171 ( .A(n18285), .B(n18284), .Y(n18331) );
  INVXL U17172 ( .A(n18333), .Y(n18286) );
  NAND2XL U17173 ( .A(n18459), .B(n18458), .Y(n18573) );
  INVXL U17174 ( .A(n18571), .Y(n18529) );
  INVXL U17175 ( .A(n18573), .Y(n18528) );
  NAND2XL U17176 ( .A(n18531), .B(n18530), .Y(n18572) );
  INVXL U17177 ( .A(n18574), .Y(n18532) );
  NOR2XL U17178 ( .A(n18571), .B(n18574), .Y(n18625) );
  NAND2XL U17179 ( .A(n18577), .B(n18576), .Y(n18626) );
  INVXL U17180 ( .A(n18681), .Y(n18629) );
  INVXL U17181 ( .A(n18678), .Y(n18630) );
  INVXL U17182 ( .A(n18680), .Y(n18633) );
  NAND2XL U17183 ( .A(n18750), .B(n18749), .Y(n18790) );
  NAND2XL U17184 ( .A(n18741), .B(n18683), .Y(n18746) );
  AOI21XL U17185 ( .A0(n18744), .A1(n18683), .B0(n18743), .Y(n18745) );
  INVXL U17186 ( .A(n18742), .Y(n18743) );
  AOI21XL U17187 ( .A0(n18792), .A1(n18748), .B0(n18791), .Y(n18842) );
  INVXL U17188 ( .A(n18790), .Y(n18791) );
  NOR2XL U17189 ( .A(n18794), .B(n18793), .Y(n18841) );
  NAND2XL U17190 ( .A(n18794), .B(n18793), .Y(n18840) );
  NAND2XL U17191 ( .A(n18845), .B(n18844), .Y(n18886) );
  AOI21XL U17192 ( .A0(n18888), .A1(n18843), .B0(n18887), .Y(n18929) );
  INVXL U17193 ( .A(n18886), .Y(n18887) );
  NOR2XL U17194 ( .A(n18890), .B(n18889), .Y(n18928) );
  NAND2XL U17195 ( .A(n18890), .B(n18889), .Y(n18927) );
  NAND2XL U17196 ( .A(n18932), .B(n18931), .Y(n18963) );
  AOI21XL U17197 ( .A0(n20463), .A1(n20462), .B0(n20461), .Y(n20499) );
  OR2XL U17198 ( .A(U1_pipe9[1]), .B(U1_pipe8[1]), .Y(n20463) );
  AND2XL U17199 ( .A(U1_pipe9[1]), .B(U1_pipe8[1]), .Y(n20461) );
  OR2XL U17200 ( .A(n28908), .B(U1_pipe8[0]), .Y(n20462) );
  NOR2XL U17201 ( .A(n20459), .B(n28900), .Y(n20498) );
  NAND2XL U17202 ( .A(n20459), .B(n28900), .Y(n20497) );
  NAND2XL U17203 ( .A(n20568), .B(n20567), .Y(n20686) );
  INVXL U17204 ( .A(n20684), .Y(n20638) );
  INVXL U17205 ( .A(n20686), .Y(n20637) );
  NAND2XL U17206 ( .A(n20640), .B(n20639), .Y(n20685) );
  INVXL U17207 ( .A(n20687), .Y(n20641) );
  INVXL U17208 ( .A(n20768), .Y(n20688) );
  NAND2XL U17209 ( .A(n20896), .B(n20895), .Y(n20981) );
  INVXL U17210 ( .A(n20978), .Y(n20942) );
  INVXL U17211 ( .A(n20981), .Y(n20941) );
  NAND2XL U17212 ( .A(n20945), .B(n20944), .Y(n20980) );
  INVXL U17213 ( .A(n20982), .Y(n20946) );
  INVXL U17214 ( .A(n20984), .Y(n20893) );
  INVXL U17215 ( .A(n20979), .Y(n20894) );
  INVXL U17216 ( .A(n21087), .Y(n21035) );
  INVXL U17217 ( .A(n21089), .Y(n21034) );
  INVXL U17218 ( .A(n21090), .Y(n21039) );
  NAND2XL U17219 ( .A(n21095), .B(n21094), .Y(n21248) );
  INVXL U17220 ( .A(n21244), .Y(n21139) );
  INVXL U17221 ( .A(n21248), .Y(n21138) );
  NAND2XL U17222 ( .A(n21142), .B(n21141), .Y(n21247) );
  INVXL U17223 ( .A(n21249), .Y(n21143) );
  INVXL U17224 ( .A(n21245), .Y(n21092) );
  INVXL U17225 ( .A(n21251), .Y(n21091) );
  NAND2XL U17226 ( .A(n21261), .B(n21260), .Y(n21280) );
  INVXL U17227 ( .A(n21280), .Y(n21351) );
  NAND2XL U17228 ( .A(n21283), .B(n21282), .Y(n21349) );
  INVXL U17229 ( .A(n21402), .Y(n21353) );
  INVXL U17230 ( .A(n21405), .Y(n21352) );
  INVXL U17231 ( .A(n21404), .Y(n21356) );
  NAND2XL U17232 ( .A(n21474), .B(n21473), .Y(n21494) );
  NAND2XL U17233 ( .A(n21465), .B(n21407), .Y(n21470) );
  AOI21XL U17234 ( .A0(n21468), .A1(n21407), .B0(n21467), .Y(n21469) );
  INVXL U17235 ( .A(n21466), .Y(n21467) );
  AOI21XL U17236 ( .A0(n21496), .A1(n21472), .B0(n21495), .Y(n21546) );
  INVXL U17237 ( .A(n21494), .Y(n21495) );
  NOR2XL U17238 ( .A(n21498), .B(n21497), .Y(n21545) );
  NAND2XL U17239 ( .A(n21498), .B(n21497), .Y(n21544) );
  NAND2XL U17240 ( .A(n21549), .B(n21548), .Y(n21588) );
  NAND2XL U17241 ( .A(n21651), .B(n21650), .Y(n21684) );
  NAND2XL U17242 ( .A(n17834), .B(n17833), .Y(n17897) );
  INVXL U17243 ( .A(n17895), .Y(n17878) );
  INVXL U17244 ( .A(n17897), .Y(n17877) );
  NAND2XL U17245 ( .A(n17880), .B(n17879), .Y(n17896) );
  INVXL U17246 ( .A(n17898), .Y(n17881) );
  INVXL U17247 ( .A(n18034), .Y(n17899) );
  INVXL U17248 ( .A(n18199), .Y(n18176) );
  NAND2XL U17249 ( .A(n18180), .B(n18179), .Y(n18198) );
  INVXL U17250 ( .A(n18200), .Y(n18181) );
  INVXL U17251 ( .A(n18341), .Y(n18291) );
  INVXL U17252 ( .A(n18343), .Y(n18290) );
  INVXL U17253 ( .A(n18344), .Y(n18295) );
  NAND2XL U17254 ( .A(n18349), .B(n18348), .Y(n18466) );
  INVXL U17255 ( .A(n18462), .Y(n18378) );
  INVXL U17256 ( .A(n18466), .Y(n18377) );
  NAND2XL U17257 ( .A(n18381), .B(n18380), .Y(n18465) );
  INVXL U17258 ( .A(n18467), .Y(n18382) );
  INVXL U17259 ( .A(n18463), .Y(n18346) );
  INVXL U17260 ( .A(n18469), .Y(n18345) );
  NAND2XL U17261 ( .A(n18478), .B(n18477), .Y(n18563) );
  INVXL U17262 ( .A(n18561), .Y(n18537) );
  INVXL U17263 ( .A(n18563), .Y(n18536) );
  NAND2XL U17264 ( .A(n18539), .B(n18538), .Y(n18562) );
  INVXL U17265 ( .A(n18564), .Y(n18540) );
  NOR2XL U17266 ( .A(n18561), .B(n18564), .Y(n18637) );
  NAND2XL U17267 ( .A(n18567), .B(n18566), .Y(n18638) );
  INVXL U17268 ( .A(n18670), .Y(n18641) );
  INVXL U17269 ( .A(n18667), .Y(n18642) );
  NAND2XL U17270 ( .A(n18644), .B(n18643), .Y(n18668) );
  INVXL U17271 ( .A(n18669), .Y(n18645) );
  NOR2XL U17272 ( .A(n18667), .B(n18669), .Y(n18728) );
  NAND2XL U17273 ( .A(n18674), .B(n18673), .Y(n18729) );
  NAND2XL U17274 ( .A(n18737), .B(n18736), .Y(n18798) );
  NAND2XL U17275 ( .A(n18837), .B(n18836), .Y(n18878) );
  AOI21XL U17276 ( .A0(n18880), .A1(n18835), .B0(n18879), .Y(n18921) );
  INVXL U17277 ( .A(n18878), .Y(n18879) );
  NOR2XL U17278 ( .A(n18882), .B(n18881), .Y(n18920) );
  NAND2XL U17279 ( .A(n18882), .B(n18881), .Y(n18919) );
  NAND2XL U17280 ( .A(n18924), .B(n18923), .Y(n18955) );
  AOI21XL U17281 ( .A0(n19382), .A1(n19381), .B0(n19380), .Y(n20476) );
  OR2XL U17282 ( .A(U1_pipe3[1]), .B(U1_pipe2[1]), .Y(n19382) );
  AND2XL U17283 ( .A(U1_pipe3[1]), .B(U1_pipe2[1]), .Y(n19380) );
  OR2XL U17284 ( .A(n28909), .B(U1_pipe2[0]), .Y(n19381) );
  NOR2XL U17285 ( .A(n19378), .B(n28901), .Y(n20475) );
  NAND2XL U17286 ( .A(n19378), .B(n28901), .Y(n20474) );
  NAND2XL U17287 ( .A(n20598), .B(n20597), .Y(n20659) );
  INVXL U17288 ( .A(n20657), .Y(n20612) );
  INVXL U17289 ( .A(n20659), .Y(n20611) );
  NAND2XL U17290 ( .A(n20614), .B(n20613), .Y(n20658) );
  INVXL U17291 ( .A(n20660), .Y(n20615) );
  INVXL U17292 ( .A(n20806), .Y(n20661) );
  NAND2XL U17293 ( .A(n20867), .B(n20866), .Y(n21003) );
  INVXL U17294 ( .A(n21000), .Y(n20911) );
  INVXL U17295 ( .A(n21003), .Y(n20910) );
  NAND2XL U17296 ( .A(n20914), .B(n20913), .Y(n21002) );
  INVXL U17297 ( .A(n21004), .Y(n20915) );
  INVXL U17298 ( .A(n21001), .Y(n20865) );
  INVXL U17299 ( .A(n21006), .Y(n20864) );
  NAND2XL U17300 ( .A(n21010), .B(n21009), .Y(n21109) );
  INVXL U17301 ( .A(n21056), .Y(n21113) );
  INVXL U17302 ( .A(n21107), .Y(n21055) );
  INVXL U17303 ( .A(n21109), .Y(n21054) );
  NAND2XL U17304 ( .A(n21058), .B(n21057), .Y(n21108) );
  INVXL U17305 ( .A(n21110), .Y(n21059) );
  INVXL U17306 ( .A(n20621), .Y(n20571) );
  NAND2XL U17307 ( .A(n20574), .B(n20573), .Y(n20620) );
  INVXL U17308 ( .A(n20622), .Y(n20575) );
  NAND2XL U17309 ( .A(n20833), .B(n20832), .Y(n20922) );
  INVXL U17310 ( .A(n20919), .Y(n20871) );
  INVXL U17311 ( .A(n20922), .Y(n20870) );
  NAND2XL U17312 ( .A(n20874), .B(n20873), .Y(n20921) );
  INVXL U17313 ( .A(n20923), .Y(n20875) );
  INVXL U17314 ( .A(n20920), .Y(n20831) );
  INVXL U17315 ( .A(n20925), .Y(n20830) );
  INVXL U17316 ( .A(n21045), .Y(n20991) );
  INVXL U17317 ( .A(n21046), .Y(n20996) );
  NAND2XL U17318 ( .A(n21051), .B(n21050), .Y(n21151) );
  INVXL U17319 ( .A(n21147), .Y(n21099) );
  INVXL U17320 ( .A(n21151), .Y(n21098) );
  NAND2XL U17321 ( .A(n21102), .B(n21101), .Y(n21150) );
  INVXL U17322 ( .A(n21152), .Y(n21103) );
  INVXL U17323 ( .A(n21154), .Y(n21047) );
  INVXL U17324 ( .A(n21148), .Y(n21048) );
  NAND2XL U17325 ( .A(n21163), .B(n21162), .Y(n21289) );
  INVXL U17326 ( .A(n21287), .Y(n21237) );
  INVXL U17327 ( .A(n21289), .Y(n21236) );
  NAND2XL U17328 ( .A(n21239), .B(n21238), .Y(n21288) );
  INVXL U17329 ( .A(n21290), .Y(n21240) );
  NOR2XL U17330 ( .A(n21287), .B(n21290), .Y(n21337) );
  NAND2XL U17331 ( .A(n21293), .B(n21292), .Y(n21338) );
  INVXL U17332 ( .A(n21394), .Y(n21341) );
  INVXL U17333 ( .A(n21391), .Y(n21342) );
  INVXL U17334 ( .A(n21393), .Y(n21345) );
  NAND2XL U17335 ( .A(n21462), .B(n21461), .Y(n21502) );
  NAND2XL U17336 ( .A(n21453), .B(n21396), .Y(n21458) );
  AOI21XL U17337 ( .A0(n21456), .A1(n21396), .B0(n21455), .Y(n21457) );
  INVXL U17338 ( .A(n21454), .Y(n21455) );
  AOI21XL U17339 ( .A0(n21504), .A1(n21460), .B0(n21503), .Y(n21554) );
  INVXL U17340 ( .A(n21502), .Y(n21503) );
  NOR2XL U17341 ( .A(n21506), .B(n21505), .Y(n21553) );
  NAND2XL U17342 ( .A(n21506), .B(n21505), .Y(n21552) );
  NAND2XL U17343 ( .A(n21557), .B(n21556), .Y(n21596) );
  AOI21XL U17344 ( .A0(n21598), .A1(n21555), .B0(n21597), .Y(n21640) );
  INVXL U17345 ( .A(n21596), .Y(n21597) );
  NOR2XL U17346 ( .A(n21600), .B(n21599), .Y(n21639) );
  NAND2XL U17347 ( .A(n21600), .B(n21599), .Y(n21638) );
  NAND2XL U17348 ( .A(n21643), .B(n21642), .Y(n21676) );
  NAND2XL U17349 ( .A(n20530), .B(n20529), .Y(n20621) );
  INVXL U17350 ( .A(n20720), .Y(n20623) );
  INVXL U17351 ( .A(n20619), .Y(n20572) );
  INVXL U17352 ( .A(n26032), .Y(n25983) );
  INVXL U17353 ( .A(n26033), .Y(n25989) );
  INVXL U17354 ( .A(n26947), .Y(n26912) );
  NAND2XL U17355 ( .A(n26911), .B(n26910), .Y(n26946) );
  NAND2XL U17356 ( .A(n26951), .B(n26950), .Y(n26986) );
  INVXL U17357 ( .A(n23174), .Y(n21732) );
  INVXL U17358 ( .A(n23131), .Y(n23166) );
  INVXL U17359 ( .A(n23360), .Y(n23320) );
  INVXL U17360 ( .A(n23362), .Y(n23319) );
  NAND2XL U17361 ( .A(n24292), .B(n24291), .Y(n24327) );
  NOR2XL U17362 ( .A(U2_A_r_d[0]), .B(n19065), .Y(n20467) );
  NAND2XL U17363 ( .A(U2_A_r_d[0]), .B(n19065), .Y(n20466) );
  INVXL U17364 ( .A(n20645), .Y(n20602) );
  INVXL U17365 ( .A(n20647), .Y(n20601) );
  INVXL U17366 ( .A(n20953), .Y(n20899) );
  INVXL U17367 ( .A(n20954), .Y(n20906) );
  NAND2XL U17368 ( .A(n21577), .B(n21576), .Y(n21612) );
  NOR2XL U17369 ( .A(U2_A_i_d[0]), .B(n16624), .Y(n17751) );
  NAND2XL U17370 ( .A(U2_A_i_d[0]), .B(n16624), .Y(n17750) );
  INVXL U17371 ( .A(n17933), .Y(n17886) );
  INVXL U17372 ( .A(n17935), .Y(n17885) );
  INVXL U17373 ( .A(n17936), .Y(n17891) );
  INVXL U17374 ( .A(n18485), .Y(n18404) );
  NAND2XL U17375 ( .A(n18856), .B(n6935), .Y(n18861) );
  NAND2XL U17376 ( .A(n18905), .B(n18865), .Y(n7376) );
  INVXL U17377 ( .A(n25799), .Y(n25837) );
  INVXL U17378 ( .A(n25845), .Y(n24411) );
  INVXL U17379 ( .A(n26030), .Y(n25984) );
  INVXL U17380 ( .A(n25087), .Y(n25080) );
  INVXL U17381 ( .A(n25079), .Y(n25088) );
  INVXL U17382 ( .A(n24865), .Y(n13530) );
  NAND2XL U17383 ( .A(n22456), .B(n29010), .Y(n24860) );
  INVXL U17384 ( .A(n24959), .Y(n24952) );
  INVXL U17385 ( .A(n24951), .Y(n24960) );
  INVXL U17386 ( .A(n22401), .Y(n22394) );
  INVXL U17387 ( .A(n22393), .Y(n22402) );
  INVXL U17388 ( .A(n22108), .Y(n22254) );
  INVXL U17389 ( .A(n22121), .Y(n22272) );
  AND2X2 U17390 ( .A(n24632), .B(n24631), .Y(n24778) );
  NAND2XL U17391 ( .A(n25062), .B(n25060), .Y(n25066) );
  NAND2XL U17392 ( .A(n24611), .B(n24610), .Y(n24813) );
  NAND2XL U17393 ( .A(n24839), .B(n25094), .Y(n25103) );
  INVXL U17394 ( .A(n25095), .Y(n24839) );
  OAI21XL U17395 ( .A0(n24465), .A1(n24453), .B0(n24452), .Y(n24463) );
  NAND2XL U17396 ( .A(n13507), .B(n24513), .Y(n24926) );
  NAND2XL U17397 ( .A(n24533), .B(n24929), .Y(n24940) );
  INVXL U17398 ( .A(n24553), .Y(n24546) );
  INVXL U17399 ( .A(n25553), .Y(n25556) );
  INVXL U17400 ( .A(n25473), .Y(n25608) );
  INVXL U17401 ( .A(n22040), .Y(n22043) );
  NAND2XL U17402 ( .A(n22054), .B(n22372), .Y(n22383) );
  INVXL U17403 ( .A(n22073), .Y(n22066) );
  NAND2XL U17404 ( .A(n22087), .B(n22407), .Y(n22415) );
  NAND2XL U17405 ( .A(n22165), .B(n22191), .Y(n22196) );
  NAND2XL U17406 ( .A(n22231), .B(n22143), .Y(n22235) );
  AND2XL U17407 ( .A(n14386), .B(U2_A_i_d[11]), .Y(n21884) );
  NAND2XL U17408 ( .A(n22242), .B(n22113), .Y(n22246) );
  INVXL U17409 ( .A(n21897), .Y(n21898) );
  NAND2XL U17410 ( .A(n21900), .B(n22109), .Y(n22255) );
  NAND2XL U17411 ( .A(n22254), .B(n22252), .Y(n22258) );
  NAND2XL U17412 ( .A(n22118), .B(n22250), .Y(n22261) );
  INVXL U17413 ( .A(n21916), .Y(n21919) );
  INVXL U17414 ( .A(n21917), .Y(n21918) );
  NAND2XL U17415 ( .A(n21920), .B(n22130), .Y(n22273) );
  NAND2XL U17416 ( .A(n22272), .B(n22270), .Y(n22276) );
  NAND2BXL U17417 ( .AN(n22323), .B(n22322), .Y(n22326) );
  NAND2XL U17418 ( .A(n21996), .B(n22329), .Y(n22335) );
  NAND2XL U17419 ( .A(n22365), .B(n22034), .Y(n22369) );
  INVXL U17420 ( .A(n25222), .Y(n25225) );
  INVXL U17421 ( .A(n25223), .Y(n25224) );
  NAND2XL U17422 ( .A(n25608), .B(n25606), .Y(n25613) );
  INVXL U17423 ( .A(n25247), .Y(n25250) );
  INVXL U17424 ( .A(n25248), .Y(n25249) );
  NAND2XL U17425 ( .A(n25270), .B(n25635), .Y(n25640) );
  INVXL U17426 ( .A(n25636), .Y(n25270) );
  NAND2X1 U17427 ( .A(n22931), .B(n5819), .Y(n23010) );
  INVXL U17428 ( .A(n23074), .Y(n23067) );
  INVXL U17429 ( .A(n23099), .Y(n23092) );
  INVXL U17430 ( .A(n23091), .Y(n23100) );
  INVXL U17431 ( .A(n22855), .Y(n22847) );
  INVXL U17432 ( .A(n22846), .Y(n22856) );
  INVXL U17433 ( .A(n25770), .Y(n25763) );
  INVXL U17434 ( .A(n25764), .Y(n25766) );
  INVXL U17435 ( .A(n25762), .Y(n25771) );
  NAND2XL U17436 ( .A(n5814), .B(n21946), .Y(n22591) );
  NAND2XL U17437 ( .A(n7735), .B(n22596), .Y(n22979) );
  INVXL U17438 ( .A(n22702), .Y(n22695) );
  INVXL U17439 ( .A(n22694), .Y(n22703) );
  NOR2XL U17440 ( .A(n22456), .B(n29009), .Y(n22459) );
  INVXL U17441 ( .A(n22518), .Y(n22513) );
  NAND2XL U17442 ( .A(n22519), .B(n22518), .Y(n22803) );
  NAND2XL U17443 ( .A(n14029), .B(n22529), .Y(n22816) );
  NAND2XL U17444 ( .A(n22541), .B(n22540), .Y(n22830) );
  NAND2XL U17445 ( .A(n22546), .B(n22545), .Y(n22834) );
  INVXL U17446 ( .A(n22564), .Y(n22557) );
  INVXL U17447 ( .A(n22558), .Y(n22560) );
  INVXL U17448 ( .A(n22556), .Y(n22565) );
  NOR2XL U17449 ( .A(n14577), .B(n24677), .Y(n12401) );
  NAND2XL U17450 ( .A(n25343), .B(n25691), .Y(n25697) );
  NAND2XL U17451 ( .A(n25433), .B(n25776), .Y(n25781) );
  INVXL U17452 ( .A(n25777), .Y(n25433) );
  NAND2XL U17453 ( .A(n25487), .B(n25578), .Y(n25583) );
  NAND2XL U17454 ( .A(n25587), .B(n25490), .Y(n25591) );
  INVXL U17455 ( .A(n20143), .Y(n20152) );
  INVXL U17456 ( .A(n20151), .Y(n20144) );
  INVXL U17457 ( .A(n20145), .Y(n20147) );
  INVXL U17458 ( .A(n20121), .Y(n20123) );
  INVXL U17459 ( .A(n17266), .Y(n17274) );
  CLKINVX2 U17460 ( .A(n17180), .Y(n17196) );
  INVXL U17461 ( .A(n17418), .Y(n17411) );
  INVXL U17462 ( .A(n17410), .Y(n17419) );
  NAND2XL U17463 ( .A(n14935), .B(n19321), .Y(n17389) );
  INVXL U17464 ( .A(n17388), .Y(n17390) );
  INVXL U17465 ( .A(n20442), .Y(n20165) );
  INVXL U17466 ( .A(n20434), .Y(n20427) );
  INVXL U17467 ( .A(n20426), .Y(n20435) );
  INVXL U17468 ( .A(n20405), .Y(n20407) );
  NAND2XL U17469 ( .A(n17285), .B(n17284), .Y(n17583) );
  INVXL U17470 ( .A(n17283), .Y(n17285) );
  NAND2XL U17471 ( .A(n17274), .B(n17273), .Y(n17572) );
  NAND2XL U17472 ( .A(n17256), .B(n17255), .Y(n17553) );
  NAND2XL U17473 ( .A(n17252), .B(n17251), .Y(n17549) );
  OR2XL U17474 ( .A(n9680), .B(U1_A_i_d0[11]), .Y(n17530) );
  NAND2XL U17475 ( .A(n17221), .B(n17220), .Y(n17512) );
  INVXL U17476 ( .A(n17706), .Y(n17715) );
  INVXL U17477 ( .A(n17714), .Y(n17707) );
  INVXL U17478 ( .A(n17708), .Y(n17710) );
  INVXL U17479 ( .A(n17699), .Y(n17717) );
  INVXL U17480 ( .A(n17682), .Y(n17691) );
  OAI21X1 U17481 ( .A0(n17603), .A1(n14512), .B0(n14511), .Y(n7932) );
  NOR2X1 U17482 ( .A(n19237), .B(n14510), .Y(n14512) );
  INVXL U17483 ( .A(n19913), .Y(n19916) );
  INVXL U17484 ( .A(n19914), .Y(n19915) );
  INVXL U17485 ( .A(n19888), .Y(n19891) );
  INVXL U17486 ( .A(n19889), .Y(n19890) );
  AOI21X2 U17487 ( .A0(n17081), .A1(n14010), .B0(n14009), .Y(n17072) );
  INVXL U17488 ( .A(n14008), .Y(n14010) );
  INVXL U17489 ( .A(n16744), .Y(n16747) );
  INVXL U17490 ( .A(n16745), .Y(n16746) );
  NOR2XL U17491 ( .A(n8652), .B(n16744), .Y(n16738) );
  INVXL U17492 ( .A(n16736), .Y(n16755) );
  INVXL U17493 ( .A(n16719), .Y(n16720) );
  OAI21XL U17494 ( .A0(n16668), .A1(n16658), .B0(n16657), .Y(n16666) );
  INVXL U17495 ( .A(n16896), .Y(n16905) );
  INVXL U17496 ( .A(n16904), .Y(n16897) );
  INVXL U17497 ( .A(n16898), .Y(n16900) );
  INVXL U17498 ( .A(n16871), .Y(n16874) );
  INVXL U17499 ( .A(n16872), .Y(n16873) );
  NAND2XL U17500 ( .A(n14513), .B(n20028), .Y(n16783) );
  NAND2XL U17501 ( .A(n20023), .B(n14972), .Y(n16782) );
  NAND2XL U17502 ( .A(n19936), .B(n20293), .Y(n20298) );
  INVXL U17503 ( .A(n20294), .Y(n19936) );
  NAND2XL U17504 ( .A(n20285), .B(n20283), .Y(n20289) );
  NAND2XL U17505 ( .A(n19919), .B(n19918), .Y(n20286) );
  INVXL U17506 ( .A(n19917), .Y(n19919) );
  INVXL U17507 ( .A(n19923), .Y(n20285) );
  INVXL U17508 ( .A(n20277), .Y(n20290) );
  NAND2XL U17509 ( .A(n19902), .B(n20263), .Y(n20274) );
  NAND2XL U17510 ( .A(n20267), .B(n20265), .Y(n20271) );
  NAND2XL U17511 ( .A(n19894), .B(n19893), .Y(n20268) );
  INVXL U17512 ( .A(n19892), .Y(n19894) );
  INVXL U17513 ( .A(n19898), .Y(n20267) );
  NAND2XL U17514 ( .A(n12300), .B(n19882), .Y(n20260) );
  NAND2XL U17515 ( .A(n20246), .B(n19868), .Y(n20250) );
  NAND2XL U17516 ( .A(n19858), .B(n20236), .Y(n20242) );
  NAND2XL U17517 ( .A(n19843), .B(n20223), .Y(n20229) );
  NAND2XL U17518 ( .A(n19818), .B(n20200), .Y(n20205) );
  NOR2X1 U17519 ( .A(n7877), .B(n19564), .Y(n7876) );
  INVXL U17520 ( .A(n19193), .Y(n19196) );
  INVXL U17521 ( .A(n19194), .Y(n19195) );
  INVXL U17522 ( .A(n19342), .Y(n19351) );
  INVXL U17523 ( .A(n19350), .Y(n19343) );
  INVXL U17524 ( .A(n19344), .Y(n19346) );
  INVXL U17525 ( .A(n19318), .Y(n19319) );
  NAND2XL U17526 ( .A(n14851), .B(n19557), .Y(n19252) );
  INVXL U17527 ( .A(n19251), .Y(n7790) );
  NOR2X1 U17528 ( .A(n7038), .B(n19236), .Y(n7904) );
  INVXL U17529 ( .A(n14864), .Y(n7854) );
  NAND2XL U17530 ( .A(n16766), .B(n17035), .Y(n17040) );
  INVXL U17531 ( .A(n17036), .Y(n16766) );
  NAND2XL U17532 ( .A(n17026), .B(n17024), .Y(n17030) );
  NAND2XL U17533 ( .A(n16749), .B(n16748), .Y(n17027) );
  INVXL U17534 ( .A(n16753), .Y(n17026) );
  NAND2XL U17535 ( .A(n16732), .B(n17004), .Y(n17015) );
  NAND2XL U17536 ( .A(n17008), .B(n17006), .Y(n17012) );
  NAND2XL U17537 ( .A(n16724), .B(n16723), .Y(n17009) );
  INVXL U17538 ( .A(n16722), .Y(n16724) );
  INVXL U17539 ( .A(n16728), .Y(n17008) );
  NAND2XL U17540 ( .A(n16988), .B(n16698), .Y(n16992) );
  NAND2XL U17541 ( .A(n6906), .B(n16661), .Y(n16962) );
  NAND2BX1 U17542 ( .AN(n16635), .B(n8631), .Y(n7534) );
  NAND2XL U17543 ( .A(n16918), .B(n17152), .Y(n17157) );
  INVXL U17544 ( .A(n17153), .Y(n16918) );
  INVXL U17545 ( .A(n17138), .Y(n17147) );
  INVXL U17546 ( .A(n17146), .Y(n17139) );
  NAND2XL U17547 ( .A(n17121), .B(n17119), .Y(n17125) );
  NAND2XL U17548 ( .A(n19217), .B(n19490), .Y(n19495) );
  INVXL U17549 ( .A(n19491), .Y(n19217) );
  NAND2XL U17550 ( .A(n19199), .B(n19198), .Y(n19483) );
  NAND2XL U17551 ( .A(n19182), .B(n19460), .Y(n19471) );
  NAND2XL U17552 ( .A(n19464), .B(n19462), .Y(n19468) );
  NAND2XL U17553 ( .A(n13680), .B(n19162), .Y(n19457) );
  NAND2XL U17554 ( .A(n19138), .B(n19435), .Y(n19440) );
  NAND2XL U17555 ( .A(n19123), .B(n19422), .Y(n19428) );
  NAND2XL U17556 ( .A(n19364), .B(n19685), .Y(n19690) );
  INVXL U17557 ( .A(n19686), .Y(n19364) );
  INVXL U17558 ( .A(n19679), .Y(n19672) );
  INVXL U17559 ( .A(n19671), .Y(n19680) );
  NAND2XL U17560 ( .A(n19654), .B(n19652), .Y(n19658) );
  NAND2XL U17561 ( .A(n19322), .B(n19526), .Y(n19655) );
  INVXL U17562 ( .A(n19524), .Y(n19654) );
  INVXL U17563 ( .A(n19588), .Y(n7271) );
  AOI22XL U17564 ( .A0(B7_q[0]), .A1(n5803), .B0(B3_q[0]), .B1(n5833), .Y(
        n11715) );
  AOI22XL U17565 ( .A0(B5_q[10]), .A1(n11864), .B0(B1_q[10]), .B1(n5832), .Y(
        n11724) );
  AOI22XL U17566 ( .A0(B3_q[11]), .A1(n5833), .B0(B0_q[11]), .B1(n5828), .Y(
        n11788) );
  AOI22XL U17567 ( .A0(B5_q[12]), .A1(n11864), .B0(B0_q[12]), .B1(n5828), .Y(
        n11832) );
  AOI22XL U17568 ( .A0(B5_q[13]), .A1(n11864), .B0(B6_q[13]), .B1(n5801), .Y(
        n11740) );
  AOI22XL U17569 ( .A0(B3_q[14]), .A1(n5833), .B0(B1_q[14]), .B1(n5832), .Y(
        n11711) );
  AOI22XL U17570 ( .A0(B7_q[15]), .A1(n5803), .B0(B0_q[15]), .B1(n5828), .Y(
        n11869) );
  AOI22XL U17571 ( .A0(B6_q[16]), .A1(n5801), .B0(B0_q[16]), .B1(n5828), .Y(
        n11865) );
  AOI22XL U17572 ( .A0(B1_q[17]), .A1(n5832), .B0(B0_q[17]), .B1(n5828), .Y(
        n11800) );
  AOI22XL U17573 ( .A0(B7_q[18]), .A1(n5803), .B0(B1_q[18]), .B1(n5832), .Y(
        n11860) );
  AOI22XL U17574 ( .A0(B6_q[19]), .A1(n5801), .B0(B7_q[19]), .B1(n5803), .Y(
        n11812) );
  AOI22XL U17575 ( .A0(B4_q[1]), .A1(n5802), .B0(B1_q[1]), .B1(n5832), .Y(
        n11668) );
  AOI22XL U17576 ( .A0(B6_q[20]), .A1(n5801), .B0(B3_q[20]), .B1(n5833), .Y(
        n11840) );
  AOI22XL U17577 ( .A0(B0_q[21]), .A1(n5828), .B0(B2_q[21]), .B1(n5831), .Y(
        n11808) );
  AOI22XL U17578 ( .A0(B7_q[22]), .A1(n5803), .B0(B1_q[22]), .B1(n5832), .Y(
        n11720) );
  AOI22XL U17579 ( .A0(B2_q[23]), .A1(n5831), .B0(B0_q[23]), .B1(n5828), .Y(
        n11804) );
  AOI22XL U17580 ( .A0(B3_q[24]), .A1(n5833), .B0(B0_q[24]), .B1(n5828), .Y(
        n11836) );
  AOI22XL U17581 ( .A0(B1_q[25]), .A1(n5832), .B0(B2_q[25]), .B1(n5831), .Y(
        n11780) );
  AOI22XL U17582 ( .A0(B6_q[26]), .A1(n5801), .B0(B4_q[26]), .B1(n5802), .Y(
        n11856) );
  AOI22XL U17583 ( .A0(B4_q[27]), .A1(n5802), .B0(B1_q[27]), .B1(n5832), .Y(
        n11736) );
  AOI22XL U17584 ( .A0(B4_q[28]), .A1(n5802), .B0(B3_q[28]), .B1(n5833), .Y(
        n11685) );
  AOI22XL U17585 ( .A0(B4_q[29]), .A1(n5802), .B0(B0_q[29]), .B1(n5828), .Y(
        n11693) );
  AOI22XL U17586 ( .A0(B0_q[2]), .A1(n5828), .B0(B1_q[2]), .B1(n5832), .Y(
        n11776) );
  AOI22XL U17587 ( .A0(B2_q[30]), .A1(n5831), .B0(B0_q[30]), .B1(n5828), .Y(
        n11792) );
  AOI22XL U17588 ( .A0(B5_q[31]), .A1(n11676), .B0(B0_q[31]), .B1(n5828), .Y(
        n11756) );
  AOI22XL U17589 ( .A0(B4_q[32]), .A1(n5802), .B0(B7_q[32]), .B1(n5803), .Y(
        n11744) );
  AOI22XL U17590 ( .A0(B7_q[33]), .A1(n5803), .B0(B1_q[33]), .B1(n5832), .Y(
        n11680) );
  AOI22XL U17591 ( .A0(B6_q[34]), .A1(n5801), .B0(B5_q[34]), .B1(n11676), .Y(
        n11728) );
  AOI22XL U17592 ( .A0(B5_q[35]), .A1(n11676), .B0(B2_q[35]), .B1(n5831), .Y(
        n11844) );
  AOI22XL U17593 ( .A0(B4_q[36]), .A1(n5802), .B0(B1_q[36]), .B1(n5832), .Y(
        n11816) );
  AOI22XL U17594 ( .A0(B7_q[37]), .A1(n5803), .B0(B1_q[37]), .B1(n5832), .Y(
        n11764) );
  AOI22XL U17595 ( .A0(B7_q[38]), .A1(n5803), .B0(B3_q[38]), .B1(n5833), .Y(
        n11748) );
  AOI22XL U17596 ( .A0(B3_q[39]), .A1(n5833), .B0(B1_q[39]), .B1(n5832), .Y(
        n11672) );
  AOI22XL U17597 ( .A0(B5_q[3]), .A1(n11676), .B0(B6_q[3]), .B1(n5801), .Y(
        n11824) );
  AOI22XL U17598 ( .A0(B7_q[40]), .A1(n5803), .B0(B0_q[40]), .B1(n5828), .Y(
        n11784) );
  AOI22XL U17599 ( .A0(B4_q[41]), .A1(n5802), .B0(B2_q[41]), .B1(n5831), .Y(
        n11852) );
  AOI22XL U17600 ( .A0(B4_q[42]), .A1(n5802), .B0(B1_q[42]), .B1(n5832), .Y(
        n11660) );
  AOI22XL U17601 ( .A0(B0_q[43]), .A1(n5828), .B0(B1_q[43]), .B1(n5832), .Y(
        n11820) );
  AOI22XL U17602 ( .A0(B0_q[44]), .A1(n5828), .B0(B3_q[44]), .B1(n5833), .Y(
        n11760) );
  AOI22XL U17603 ( .A0(B4_q[45]), .A1(n5802), .B0(B7_q[45]), .B1(n5803), .Y(
        n11701) );
  AOI22XL U17604 ( .A0(B6_q[46]), .A1(n5801), .B0(B1_q[46]), .B1(n5832), .Y(
        n11705) );
  AOI22XL U17605 ( .A0(B5_q[47]), .A1(n11676), .B0(B1_q[47]), .B1(n5832), .Y(
        n11656) );
  AOI22XL U17606 ( .A0(B5_q[48]), .A1(n11676), .B0(B1_q[48]), .B1(n5832), .Y(
        n11689) );
  AOI22XL U17607 ( .A0(B5_q[49]), .A1(n11676), .B0(B7_q[49]), .B1(n5803), .Y(
        n11752) );
  AOI22XL U17608 ( .A0(B5_q[4]), .A1(n11676), .B0(B7_q[4]), .B1(n5803), .Y(
        n11732) );
  AOI22XL U17609 ( .A0(B5_q[50]), .A1(n11676), .B0(B1_q[50]), .B1(n5832), .Y(
        n11697) );
  AOI22XL U17610 ( .A0(B6_q[51]), .A1(n5801), .B0(B7_q[51]), .B1(n5803), .Y(
        n11768) );
  AOI22XL U17611 ( .A0(B2_q[5]), .A1(n5831), .B0(B0_q[5]), .B1(n5828), .Y(
        n11796) );
  AOI22XL U17612 ( .A0(B6_q[6]), .A1(n5801), .B0(B4_q[6]), .B1(n5802), .Y(
        n11848) );
  AOI22XL U17613 ( .A0(B5_q[7]), .A1(n11676), .B0(B1_q[7]), .B1(n5832), .Y(
        n11664) );
  AOI22XL U17614 ( .A0(B5_q[8]), .A1(n11676), .B0(B2_q[8]), .B1(n5831), .Y(
        n11772) );
  AOI22XL U17615 ( .A0(B1_q[9]), .A1(n5832), .B0(B2_q[9]), .B1(n5831), .Y(
        n11828) );
  NAND2XL U17616 ( .A(n11956), .B(n28669), .Y(n28670) );
  NAND2XL U17617 ( .A(n11956), .B(n28667), .Y(n28668) );
  NAND2XL U17618 ( .A(n28666), .B(n28665), .Y(n28667) );
  INVXL U17619 ( .A(n28663), .Y(n28664) );
  INVXL U17620 ( .A(n28661), .Y(n28662) );
  OAI2BB1XL U17621 ( .A0N(n28666), .A1N(n28659), .B0(n11956), .Y(n28660) );
  NAND2XL U17622 ( .A(n11956), .B(n28657), .Y(n28658) );
  AND2X1 U17623 ( .A(n5808), .B(n15025), .Y(n11997) );
  INVXL U17624 ( .A(n28650), .Y(n28654) );
  INVXL U17625 ( .A(n28648), .Y(n28652) );
  NAND2XL U17626 ( .A(n11956), .B(n28640), .Y(n28651) );
  INVXL U17627 ( .A(n28645), .Y(n28649) );
  NAND2XL U17628 ( .A(n28661), .B(n28643), .Y(n28656) );
  NAND2XL U17629 ( .A(n28663), .B(n28643), .Y(n28647) );
  NAND2BXL U17630 ( .AN(n28651), .B(n28641), .Y(n28655) );
  NAND2XL U17631 ( .A(n28650), .B(n28641), .Y(n28646) );
  NAND2XL U17632 ( .A(n28645), .B(n28638), .Y(n28653) );
  NAND2XL U17633 ( .A(n28648), .B(n28638), .Y(n28644) );
  NOR2XL U17634 ( .A(n28706), .B(n28635), .Y(n11996) );
  NOR2XL U17635 ( .A(n28631), .B(n11996), .Y(n28634) );
  NOR2XL U17636 ( .A(n28703), .B(n14977), .Y(n11972) );
  NOR2XL U17637 ( .A(n11986), .B(n11988), .Y(n11987) );
  NOR2XL U17638 ( .A(n11986), .B(n11982), .Y(n11981) );
  INVXL U17639 ( .A(n11992), .Y(n11645) );
  INVXL U17640 ( .A(n11993), .Y(n11646) );
  NOR2XL U17641 ( .A(n15027), .B(n28669), .Y(n11621) );
  OAI211XL U17642 ( .A0(n5836), .A1(n16494), .B0(n15152), .C0(n15151), .Y(
        n15153) );
  AOI21XL U17643 ( .A0(B0_q[19]), .A1(n5925), .B0(n5924), .Y(n15151) );
  AOI22XL U17644 ( .A0(B3_q[19]), .A1(n15982), .B0(B2_q[19]), .B1(n15958), .Y(
        n15152) );
  NAND4XL U17645 ( .A(n15011), .B(n15010), .C(n5913), .D(n15009), .Y(n15012)
         );
  NAND2XL U17646 ( .A(B6_q[35]), .B(n16570), .Y(n15011) );
  NAND2XL U17647 ( .A(B5_q[35]), .B(n16559), .Y(n15010) );
  OAI211XL U17648 ( .A0(n15495), .A1(n16287), .B0(n16099), .C0(n16098), .Y(
        n16100) );
  AOI21XL U17649 ( .A0(B0_q[18]), .A1(n5933), .B0(n16496), .Y(n16098) );
  AOI22XL U17650 ( .A0(B3_q[18]), .A1(n16158), .B0(B1_q[18]), .B1(n16165), .Y(
        n16099) );
  NAND4XL U17651 ( .A(n15328), .B(n15327), .C(n5800), .D(n15326), .Y(n15329)
         );
  NAND2XL U17652 ( .A(B4_q[37]), .B(n7126), .Y(n15328) );
  NAND2XL U17653 ( .A(B5_q[37]), .B(n16375), .Y(n15327) );
  NAND4XL U17654 ( .A(n15290), .B(n15289), .C(n5909), .D(n15288), .Y(n15291)
         );
  NAND2XL U17655 ( .A(B7_q[42]), .B(n7127), .Y(n15290) );
  NAND2XL U17656 ( .A(B5_q[42]), .B(n16559), .Y(n15289) );
  OAI211XL U17657 ( .A0(n5836), .A1(n15847), .B0(n15846), .C0(n15845), .Y(
        n15848) );
  AOI21XL U17658 ( .A0(B4_q[33]), .A1(n5925), .B0(n5924), .Y(n15845) );
  AOI22XL U17659 ( .A0(B7_q[33]), .A1(n5930), .B0(B6_q[33]), .B1(n15958), .Y(
        n15846) );
  NAND4XL U17660 ( .A(n15709), .B(n15708), .C(n6880), .D(n15707), .Y(n15710)
         );
  NAND2XL U17661 ( .A(B6_q[16]), .B(n16293), .Y(n15709) );
  NAND2XL U17662 ( .A(B4_q[16]), .B(n16277), .Y(n15708) );
  OAI211XL U17663 ( .A0(n5806), .A1(n15819), .B0(n15429), .C0(n15428), .Y(
        n15430) );
  AOI22XL U17664 ( .A0(B7_q[40]), .A1(n16128), .B0(B6_q[40]), .B1(n16143), .Y(
        n15429) );
  NAND4XL U17665 ( .A(n15915), .B(n15914), .C(n5800), .D(n15913), .Y(n15916)
         );
  NAND2XL U17666 ( .A(B4_q[16]), .B(n15969), .Y(n15915) );
  NAND2XL U17667 ( .A(B5_q[16]), .B(n15963), .Y(n15914) );
  OAI211XL U17668 ( .A0(n15967), .A1(n16107), .B0(n15162), .C0(n15161), .Y(
        n15163) );
  AOI21XL U17669 ( .A0(B1_q[16]), .A1(n15963), .B0(n5924), .Y(n15161) );
  AOI22XL U17670 ( .A0(B2_q[16]), .A1(n15958), .B0(B0_q[16]), .B1(n5925), .Y(
        n15162) );
  NAND4XL U17671 ( .A(n15522), .B(n15521), .C(n6880), .D(n15520), .Y(n15523)
         );
  NAND2XL U17672 ( .A(B6_q[15]), .B(n15431), .Y(n15522) );
  NAND2XL U17673 ( .A(B5_q[15]), .B(n16165), .Y(n15521) );
  OAI211XL U17674 ( .A0(n5813), .A1(n15701), .B0(n15700), .C0(n15699), .Y(
        n15702) );
  AOI21XL U17675 ( .A0(B7_q[18]), .A1(n16325), .B0(n5924), .Y(n15699) );
  AOI22XL U17676 ( .A0(B6_q[18]), .A1(n16354), .B0(B4_q[18]), .B1(n15687), .Y(
        n15700) );
  NAND4XL U17677 ( .A(n15697), .B(n15696), .C(n5800), .D(n15695), .Y(n15698)
         );
  NAND2XL U17678 ( .A(B4_q[19]), .B(n16277), .Y(n15697) );
  NAND2XL U17679 ( .A(B5_q[19]), .B(n15747), .Y(n15696) );
  INVXL U17680 ( .A(T1_rom3_q[15]), .Y(n29138) );
  INVXL U17681 ( .A(T1_rom1_q[11]), .Y(n29206) );
  INVXL U17682 ( .A(T1_rom1_q[9]), .Y(n29177) );
  NAND4XL U17683 ( .A(n15537), .B(n15536), .C(n5800), .D(n15535), .Y(n15538)
         );
  NAND2XL U17684 ( .A(B5_q[11]), .B(n16165), .Y(n15537) );
  NAND2XL U17685 ( .A(B7_q[11]), .B(n16158), .Y(n15536) );
  OAI211XL U17686 ( .A0(n5813), .A1(n15985), .B0(n15771), .C0(n15770), .Y(
        n15772) );
  AOI21XL U17687 ( .A0(B4_q[0]), .A1(n15687), .B0(n16461), .Y(n15770) );
  AOI22XL U17688 ( .A0(B7_q[0]), .A1(n16325), .B0(B6_q[0]), .B1(n5926), .Y(
        n15771) );
  INVXL U17689 ( .A(T1_rom1_q[27]), .Y(n29189) );
  OAI211XL U17690 ( .A0(n15633), .A1(n15721), .B0(n15720), .C0(n15719), .Y(
        n15722) );
  AOI21XL U17691 ( .A0(B4_q[13]), .A1(n15687), .B0(n5924), .Y(n15719) );
  AOI22XL U17692 ( .A0(B5_q[13]), .A1(n16344), .B0(B7_q[13]), .B1(n16325), .Y(
        n15720) );
  NAND4XL U17693 ( .A(n15863), .B(n15862), .C(n5800), .D(n15861), .Y(n15864)
         );
  NAND2XL U17694 ( .A(B4_q[29]), .B(n15969), .Y(n15863) );
  NAND2XL U17695 ( .A(B7_q[29]), .B(n15982), .Y(n15862) );
  NAND4XL U17696 ( .A(n15754), .B(n15753), .C(n6880), .D(n15752), .Y(n15755)
         );
  NAND2XL U17697 ( .A(B4_q[5]), .B(n15687), .Y(n15754) );
  NAND2XL U17698 ( .A(B5_q[5]), .B(n16344), .Y(n15753) );
  OAI211XL U17699 ( .A0(n5813), .A1(n15815), .B0(n15617), .C0(n15616), .Y(
        n15618) );
  AOI21XL U17700 ( .A0(B6_q[41]), .A1(n5926), .B0(n28985), .Y(n15616) );
  AOI22XL U17701 ( .A0(B4_q[41]), .A1(n15687), .B0(B7_q[41]), .B1(n16325), .Y(
        n15617) );
  INVXL U17702 ( .A(T1_rom3_q[25]), .Y(n29127) );
  OAI211XL U17703 ( .A0(n5813), .A1(n15972), .B0(n15761), .C0(n15760), .Y(
        n15762) );
  AOI21XL U17704 ( .A0(B7_q[3]), .A1(n16325), .B0(n16470), .Y(n15760) );
  AOI22XL U17705 ( .A0(B4_q[3]), .A1(n15687), .B0(B6_q[3]), .B1(n5926), .Y(
        n15761) );
  INVXL U17706 ( .A(T1_rom1_q[25]), .Y(n29191) );
  AOI22XL U17707 ( .A0(B1_q[35]), .A1(n15963), .B0(B3_q[35]), .B1(n15982), .Y(
        n15096) );
  AOI21XL U17708 ( .A0(n15958), .A1(B2_q[35]), .B0(n15095), .Y(n15097) );
  INVXL U17709 ( .A(T1_rom0_q[25]), .Y(n29223) );
  OAI211XL U17710 ( .A0(n5806), .A1(n15859), .B0(n15465), .C0(n15464), .Y(
        n15466) );
  AOI22XL U17711 ( .A0(B6_q[30]), .A1(n16143), .B0(B7_q[30]), .B1(n16128), .Y(
        n15465) );
  AOI21XL U17712 ( .A0(B4_q[30]), .A1(n5933), .B0(n28985), .Y(n15464) );
  OAI211XL U17713 ( .A0(n16348), .A1(n16226), .B0(n16225), .C0(n16224), .Y(
        n16227) );
  AOI21XL U17714 ( .A0(B0_q[35]), .A1(n16277), .B0(n5924), .Y(n16224) );
  AOI22XL U17715 ( .A0(B1_q[35]), .A1(n16344), .B0(B2_q[35]), .B1(n16354), .Y(
        n16225) );
  OAI211XL U17716 ( .A0(n5836), .A1(n16543), .B0(n15195), .C0(n15194), .Y(
        n15196) );
  AOI21XL U17717 ( .A0(B0_q[7]), .A1(n5925), .B0(n5924), .Y(n15194) );
  AOI22XL U17718 ( .A0(B2_q[7]), .A1(n15958), .B0(B3_q[7]), .B1(n15982), .Y(
        n15195) );
  INVXL U17719 ( .A(T1_rom0_q[23]), .Y(n29225) );
  INVXL U17720 ( .A(T1_rom2_q[23]), .Y(n29161) );
  OAI211XL U17721 ( .A0(n15967), .A1(n15966), .B0(n15965), .C0(n15964), .Y(
        n15968) );
  AOI21XL U17722 ( .A0(B4_q[4]), .A1(n15969), .B0(n16496), .Y(n15964) );
  AOI22XL U17723 ( .A0(B6_q[4]), .A1(n15958), .B0(B5_q[4]), .B1(n15963), .Y(
        n15965) );
  OAI211XL U17724 ( .A0(n15967), .A1(n16205), .B0(n15077), .C0(n15076), .Y(
        n15078) );
  AOI21XL U17725 ( .A0(B2_q[41]), .A1(n15958), .B0(n5924), .Y(n15076) );
  AOI22XL U17726 ( .A0(B0_q[41]), .A1(n5925), .B0(B1_q[41]), .B1(n15963), .Y(
        n15077) );
  OAI211XL U17727 ( .A0(n15948), .A1(n15127), .B0(n15126), .C0(n15125), .Y(
        n15128) );
  AOI21XL U17728 ( .A0(B0_q[26]), .A1(n5925), .B0(n5924), .Y(n15125) );
  AOI22XL U17729 ( .A0(B3_q[26]), .A1(n15982), .B0(B1_q[26]), .B1(n15963), .Y(
        n15126) );
  OAI211XL U17730 ( .A0(n5841), .A1(n16034), .B0(n16033), .C0(n16032), .Y(
        n16035) );
  AOI21XL U17731 ( .A0(B0_q[37]), .A1(n5933), .B0(n5924), .Y(n16032) );
  AOI22XL U17732 ( .A0(B1_q[37]), .A1(n16165), .B0(B2_q[37]), .B1(n16143), .Y(
        n16033) );
  NAND4XL U17733 ( .A(n15660), .B(n15659), .C(n5800), .D(n15658), .Y(n15661)
         );
  NAND2XL U17734 ( .A(B4_q[29]), .B(n16277), .Y(n15660) );
  NAND2XL U17735 ( .A(B7_q[29]), .B(n16325), .Y(n15659) );
  INVXL U17736 ( .A(T1_rom1_q[23]), .Y(n29193) );
  OAI211XL U17737 ( .A0(n5813), .A1(n15859), .B0(n15656), .C0(n15655), .Y(
        n15657) );
  AOI22XL U17738 ( .A0(B6_q[30]), .A1(n16354), .B0(B7_q[30]), .B1(n16325), .Y(
        n15656) );
  OAI211XL U17739 ( .A0(n16348), .A1(n15610), .B0(n15609), .C0(n15608), .Y(
        n15611) );
  AOI21XL U17740 ( .A0(B4_q[43]), .A1(n15687), .B0(n16496), .Y(n15608) );
  AOI22XL U17741 ( .A0(B5_q[43]), .A1(n16344), .B0(B6_q[43]), .B1(n16354), .Y(
        n15609) );
  OAI211XL U17742 ( .A0(n5813), .A1(n15819), .B0(n15620), .C0(n15619), .Y(
        n15621) );
  AOI21XL U17743 ( .A0(B4_q[40]), .A1(n15687), .B0(n5924), .Y(n15619) );
  AOI22XL U17744 ( .A0(B7_q[40]), .A1(n16325), .B0(B6_q[40]), .B1(n5926), .Y(
        n15620) );
  OAI211XL U17745 ( .A0(n16348), .A1(n15664), .B0(n15663), .C0(n15662), .Y(
        n15665) );
  AOI21XL U17746 ( .A0(B4_q[28]), .A1(n15687), .B0(n5924), .Y(n15662) );
  AOI22XL U17747 ( .A0(B6_q[28]), .A1(n16354), .B0(B5_q[28]), .B1(n16344), .Y(
        n15663) );
  NAND4XL U17748 ( .A(n15631), .B(n15630), .C(n5800), .D(n15629), .Y(n15632)
         );
  NAND2XL U17749 ( .A(B4_q[37]), .B(n16277), .Y(n15631) );
  NAND2XL U17750 ( .A(B5_q[37]), .B(n15747), .Y(n15630) );
  OAI211XL U17751 ( .A0(n5813), .A1(n15650), .B0(n15649), .C0(n15648), .Y(
        n15651) );
  AOI22XL U17752 ( .A0(B6_q[32]), .A1(n16354), .B0(B4_q[32]), .B1(n15687), .Y(
        n15649) );
  NAND4XL U17753 ( .A(n15668), .B(n15667), .C(n5909), .D(n15666), .Y(n15669)
         );
  NAND2XL U17754 ( .A(B6_q[27]), .B(n16293), .Y(n15668) );
  NAND2XL U17755 ( .A(B4_q[27]), .B(n16277), .Y(n15667) );
  OAI211XL U17756 ( .A0(n5813), .A1(n15855), .B0(n15653), .C0(n15652), .Y(
        n15654) );
  AOI22XL U17757 ( .A0(B4_q[31]), .A1(n15687), .B0(B6_q[31]), .B1(n16354), .Y(
        n15653) );
  NAND4XL U17758 ( .A(n15871), .B(n15870), .C(n5908), .D(n15869), .Y(n15872)
         );
  NAND2XL U17759 ( .A(B4_q[27]), .B(n5925), .Y(n15871) );
  NAND2XL U17760 ( .A(B7_q[27]), .B(n15982), .Y(n15870) );
  NAND4XL U17761 ( .A(n15123), .B(n15122), .C(n5800), .D(n15121), .Y(n15124)
         );
  NAND2XL U17762 ( .A(B3_q[27]), .B(n15982), .Y(n15123) );
  NAND2XL U17763 ( .A(B1_q[27]), .B(n15963), .Y(n15122) );
  AOI21XL U17764 ( .A0(B2_q[32]), .A1(n15958), .B0(n15105), .Y(n15106) );
  NAND2XL U17765 ( .A(R7_valid), .B(n15104), .Y(n15105) );
  NAND2XL U17766 ( .A(n6880), .B(n16050), .Y(n16051) );
  AOI22XL U17767 ( .A0(B2_q[30]), .A1(n15958), .B0(B0_q[30]), .B1(n5925), .Y(
        n15113) );
  AOI21XL U17768 ( .A0(n15982), .A1(B3_q[30]), .B0(n15112), .Y(n15114) );
  OAI211XL U17769 ( .A0(n5836), .A1(n16435), .B0(n15102), .C0(n15101), .Y(
        n15103) );
  AOI21XL U17770 ( .A0(B0_q[33]), .A1(n5925), .B0(n5924), .Y(n15101) );
  AOI22XL U17771 ( .A0(B2_q[33]), .A1(n15958), .B0(B3_q[33]), .B1(n15982), .Y(
        n15102) );
  OAI211XL U17772 ( .A0(n15967), .A1(n15851), .B0(n15850), .C0(n15849), .Y(
        n15852) );
  AOI21XL U17773 ( .A0(B5_q[32]), .A1(n15179), .B0(n5924), .Y(n15849) );
  AOI22XL U17774 ( .A0(B6_q[32]), .A1(n15958), .B0(B4_q[32]), .B1(n5925), .Y(
        n15850) );
  OAI211XL U17775 ( .A0(n5836), .A1(n15855), .B0(n15854), .C0(n15853), .Y(
        n15856) );
  AOI21XL U17776 ( .A0(B6_q[31]), .A1(n15958), .B0(n5924), .Y(n15853) );
  AOI22XL U17777 ( .A0(B7_q[31]), .A1(n15982), .B0(B4_q[31]), .B1(n5925), .Y(
        n15854) );
  OAI211XL U17778 ( .A0(n5806), .A1(n15650), .B0(n15459), .C0(n15458), .Y(
        n15460) );
  AOI22XL U17779 ( .A0(B4_q[32]), .A1(n15557), .B0(B7_q[32]), .B1(n16128), .Y(
        n15459) );
  AOI21XL U17780 ( .A0(B6_q[32]), .A1(n16161), .B0(n28985), .Y(n15458) );
  INVXL U17781 ( .A(T1_rom3_q[8]), .Y(n29114) );
  OAI211XL U17782 ( .A0(n15387), .A1(n5914), .B0(n15386), .C0(n15385), .Y(
        n15388) );
  AOI22XL U17783 ( .A0(B7_q[0]), .A1(n7127), .B0(B5_q[0]), .B1(n16559), .Y(
        n15386) );
  INVXL U17784 ( .A(n19581), .Y(n19245) );
  XOR2X1 U17785 ( .A(n7419), .B(n22974), .Y(n7418) );
  INVXL U17786 ( .A(n25660), .Y(n25295) );
  XNOR2X1 U17787 ( .A(n25306), .B(n25305), .Y(n25307) );
  INVXL U17788 ( .A(n25666), .Y(n25305) );
  XNOR2X1 U17789 ( .A(n25313), .B(n25312), .Y(n25314) );
  INVXL U17790 ( .A(n25671), .Y(n25312) );
  INVXL U17791 ( .A(n20342), .Y(n20043) );
  INVXL U17792 ( .A(n20339), .Y(n20034) );
  INVXL U17793 ( .A(n24998), .Y(n24722) );
  XNOR2X1 U17794 ( .A(n14891), .B(n14890), .Y(n14892) );
  NAND2XL U17795 ( .A(n7025), .B(n20312), .Y(n14890) );
  INVXL U17796 ( .A(n19611), .Y(n19269) );
  XNOR2X1 U17797 ( .A(n24718), .B(n24717), .Y(n24719) );
  INVXL U17798 ( .A(n24994), .Y(n24717) );
  AOI21XL U17799 ( .A0(n24750), .A1(n5794), .B0(n24743), .Y(n24746) );
  XNOR2X1 U17800 ( .A(n22606), .B(n22605), .Y(n22607) );
  NAND2XL U17801 ( .A(n22604), .B(n22603), .Y(n22605) );
  XNOR2X1 U17802 ( .A(n24708), .B(n24707), .Y(n24709) );
  NAND2XL U17803 ( .A(n17330), .B(n17329), .Y(n17331) );
  XNOR2X1 U17804 ( .A(n22610), .B(n22991), .Y(n22611) );
  INVXL U17805 ( .A(n19621), .Y(n19283) );
  NAND2X1 U17806 ( .A(n20328), .B(n7337), .Y(n7219) );
  NAND2XL U17807 ( .A(n19263), .B(n19262), .Y(n19264) );
  XNOR2X1 U17808 ( .A(n12648), .B(n12647), .Y(n12649) );
  NAND2XL U17809 ( .A(n14117), .B(n14114), .Y(n12647) );
  INVXL U17810 ( .A(n19614), .Y(n19273) );
  INVXL U17811 ( .A(n16952), .Y(n16649) );
  OAI211XL U17812 ( .A0(n5813), .A1(n15847), .B0(n15646), .C0(n15645), .Y(
        n15647) );
  AOI22XL U17813 ( .A0(B7_q[33]), .A1(n16325), .B0(B4_q[33]), .B1(n15687), .Y(
        n15646) );
  OAI211XL U17814 ( .A0(n5813), .A1(n16447), .B0(n16243), .C0(n16242), .Y(
        n16244) );
  AOI21XL U17815 ( .A0(B3_q[30]), .A1(n16325), .B0(n5924), .Y(n16242) );
  AOI22XL U17816 ( .A0(B2_q[30]), .A1(n16354), .B0(B0_q[30]), .B1(n15687), .Y(
        n16243) );
  NAND4XL U17817 ( .A(n15639), .B(n15638), .C(n6880), .D(n15637), .Y(n15640)
         );
  NAND2XL U17818 ( .A(B4_q[35]), .B(n16277), .Y(n15639) );
  NAND2XL U17819 ( .A(B6_q[35]), .B(n5926), .Y(n15638) );
  NAND4XL U17820 ( .A(n15442), .B(n15441), .C(n6880), .D(n15440), .Y(n15443)
         );
  NAND2XL U17821 ( .A(B7_q[37]), .B(n16158), .Y(n15442) );
  NAND2XL U17822 ( .A(B5_q[37]), .B(n16165), .Y(n15441) );
  OAI211XL U17823 ( .A0(n5806), .A1(n16447), .B0(n16059), .C0(n16058), .Y(
        n16060) );
  AOI21XL U17824 ( .A0(B0_q[30]), .A1(n5933), .B0(n5924), .Y(n16058) );
  AOI22XL U17825 ( .A0(B2_q[30]), .A1(n16143), .B0(B3_q[30]), .B1(n16128), .Y(
        n16059) );
  OAI2BB1XL U17826 ( .A0N(n28706), .A1N(n28635), .B0(n28634), .Y(n5671) );
  OAI211XL U17827 ( .A0(n15835), .A1(n5813), .B0(n15635), .C0(n15634), .Y(
        n15636) );
  AOI22XL U17828 ( .A0(B6_q[36]), .A1(n16354), .B0(B7_q[36]), .B1(n16325), .Y(
        n15635) );
  OAI211XL U17829 ( .A0(n5813), .A1(n15823), .B0(n15623), .C0(n15622), .Y(
        n15624) );
  AOI22XL U17830 ( .A0(B7_q[39]), .A1(n16325), .B0(B6_q[39]), .B1(n16354), .Y(
        n15623) );
  AOI21XL U17831 ( .A0(B4_q[39]), .A1(n15687), .B0(n28985), .Y(n15622) );
  NAND4XL U17832 ( .A(n15627), .B(n15626), .C(n5800), .D(n15625), .Y(n15628)
         );
  NAND2XL U17833 ( .A(B6_q[38]), .B(n5926), .Y(n15627) );
  NAND2XL U17834 ( .A(B4_q[38]), .B(n16277), .Y(n15626) );
  OAI211XL U17835 ( .A0(n16435), .A1(n5813), .B0(n16232), .C0(n16231), .Y(
        n16233) );
  AOI21XL U17836 ( .A0(B0_q[33]), .A1(n15687), .B0(n5924), .Y(n16231) );
  AOI22XL U17837 ( .A0(B2_q[33]), .A1(n16354), .B0(B3_q[33]), .B1(n16325), .Y(
        n16232) );
  INVXL U17838 ( .A(T1_rom2_q[27]), .Y(n29157) );
  INVXL U17839 ( .A(T1_rom2_q[26]), .Y(n29158) );
  NAND4XL U17840 ( .A(n15606), .B(n15605), .C(n5906), .D(n15604), .Y(n15607)
         );
  NAND2XL U17841 ( .A(B7_q[44]), .B(n16325), .Y(n15606) );
  NAND2XL U17842 ( .A(B5_q[44]), .B(n15747), .Y(n15605) );
  OAI211XL U17843 ( .A0(n5836), .A1(n15835), .B0(n15834), .C0(n15833), .Y(
        n15836) );
  AOI22XL U17844 ( .A0(B6_q[36]), .A1(n15958), .B0(B7_q[36]), .B1(n5930), .Y(
        n15834) );
  AOI21XL U17845 ( .A0(B4_q[36]), .A1(n15969), .B0(n28985), .Y(n15833) );
  OAI211XL U17846 ( .A0(n16348), .A1(n15799), .B0(n15602), .C0(n15601), .Y(
        n15603) );
  AOI21XL U17847 ( .A0(B4_q[45]), .A1(n15687), .B0(n16496), .Y(n15601) );
  AOI22XL U17848 ( .A0(B5_q[45]), .A1(n16344), .B0(B6_q[45]), .B1(n16354), .Y(
        n15602) );
  INVXL U17849 ( .A(T1_rom1_q[19]), .Y(n29198) );
  OAI211XL U17850 ( .A0(n5836), .A1(n15859), .B0(n15858), .C0(n15857), .Y(
        n15860) );
  AOI22XL U17851 ( .A0(B6_q[30]), .A1(n15958), .B0(B7_q[30]), .B1(n15982), .Y(
        n15858) );
  OAI211XL U17852 ( .A0(n16163), .A1(n15815), .B0(n15426), .C0(n15425), .Y(
        n15427) );
  AOI22XL U17853 ( .A0(B4_q[41]), .A1(n15557), .B0(B7_q[41]), .B1(n16128), .Y(
        n15426) );
  OAI2BB2XL U17854 ( .B0(n5909), .B1(AOPD[44]), .A0N(n16012), .A1N(n16011), 
        .Y(n3374) );
  AOI22XL U17855 ( .A0(B0_q[44]), .A1(n15557), .B0(B2_q[44]), .B1(n16143), .Y(
        n16011) );
  AOI21XL U17856 ( .A0(n16136), .A1(B3_q[44]), .B0(n16010), .Y(n16012) );
  OAI211XL U17857 ( .A0(n5841), .A1(n15799), .B0(n15412), .C0(n15411), .Y(
        n15413) );
  AOI21XL U17858 ( .A0(B4_q[45]), .A1(n5933), .B0(n16496), .Y(n15411) );
  AOI22XL U17859 ( .A0(B5_q[45]), .A1(n16165), .B0(B6_q[45]), .B1(n16143), .Y(
        n15412) );
  NAND4XL U17860 ( .A(n16240), .B(n16239), .C(n5910), .D(n16238), .Y(n16241)
         );
  NAND2XL U17861 ( .A(B2_q[31]), .B(n16293), .Y(n16240) );
  NAND2XL U17862 ( .A(B0_q[31]), .B(n16277), .Y(n16239) );
  NAND4XL U17863 ( .A(n16056), .B(n16055), .C(n5907), .D(n16054), .Y(n16057)
         );
  NAND2XL U17864 ( .A(B1_q[31]), .B(n16165), .Y(n16056) );
  NAND2XL U17865 ( .A(B0_q[31]), .B(n15557), .Y(n16055) );
  OAI211XL U17866 ( .A0(n15967), .A1(n15799), .B0(n15798), .C0(n15797), .Y(
        n15800) );
  AOI21XL U17867 ( .A0(B4_q[45]), .A1(n5925), .B0(n16496), .Y(n15797) );
  AOI22XL U17868 ( .A0(B5_q[45]), .A1(n15963), .B0(B6_q[45]), .B1(n15958), .Y(
        n15798) );
  OAI211XL U17869 ( .A0(n5841), .A1(n16048), .B0(n16047), .C0(n16046), .Y(
        n16049) );
  AOI21XL U17870 ( .A0(B1_q[33]), .A1(n16165), .B0(n5924), .Y(n16046) );
  AOI22XL U17871 ( .A0(B2_q[33]), .A1(n16161), .B0(B0_q[33]), .B1(n15557), .Y(
        n16047) );
  INVXL U17872 ( .A(T1_rom1_q[18]), .Y(n29199) );
  NAND4XL U17873 ( .A(n15110), .B(n15109), .C(n5800), .D(n15108), .Y(n15111)
         );
  NAND2XL U17874 ( .A(B3_q[31]), .B(n15982), .Y(n15110) );
  NAND2XL U17875 ( .A(B0_q[31]), .B(n5925), .Y(n15109) );
  OAI2BB2XL U17876 ( .B0(n5909), .B1(AOPD[7]), .A0N(n16138), .A1N(n16137), .Y(
        n3418) );
  AOI22XL U17877 ( .A0(B2_q[7]), .A1(n16143), .B0(B0_q[7]), .B1(n15557), .Y(
        n16137) );
  AOI21XL U17878 ( .A0(n16136), .A1(B3_q[7]), .B0(n16135), .Y(n16138) );
  OAI211XL U17879 ( .A0(n5813), .A1(n16410), .B0(n16211), .C0(n16210), .Y(
        n16212) );
  AOI21XL U17880 ( .A0(B2_q[39]), .A1(n5926), .B0(n5924), .Y(n16210) );
  AOI22XL U17881 ( .A0(B3_q[39]), .A1(n16325), .B0(B0_q[39]), .B1(n15687), .Y(
        n16211) );
  OAI211XL U17882 ( .A0(n5806), .A1(n15855), .B0(n15462), .C0(n15461), .Y(
        n15463) );
  AOI21XL U17883 ( .A0(B6_q[31]), .A1(n16161), .B0(n16487), .Y(n15461) );
  AOI22XL U17884 ( .A0(B7_q[31]), .A1(n16128), .B0(B4_q[31]), .B1(n15557), .Y(
        n15462) );
  INVXL U17885 ( .A(T1_rom0_q[19]), .Y(n29230) );
  OAI211XL U17886 ( .A0(n15446), .A1(n5841), .B0(n15445), .C0(n15444), .Y(
        n15447) );
  AOI21XL U17887 ( .A0(B5_q[36]), .A1(n16165), .B0(n5924), .Y(n15444) );
  AOI22XL U17888 ( .A0(B6_q[36]), .A1(n16143), .B0(B4_q[36]), .B1(n15557), .Y(
        n15445) );
  OAI211XL U17889 ( .A0(n16215), .A1(n16348), .B0(n16214), .C0(n16213), .Y(
        n16216) );
  AOI21XL U17890 ( .A0(B0_q[38]), .A1(n15687), .B0(n5924), .Y(n16213) );
  AOI22XL U17891 ( .A0(B2_q[38]), .A1(n16354), .B0(B1_q[38]), .B1(n16344), .Y(
        n16214) );
  OAI211XL U17892 ( .A0(n5806), .A1(n16406), .B0(n16024), .C0(n16023), .Y(
        n16025) );
  AOI21XL U17893 ( .A0(B0_q[40]), .A1(n15557), .B0(n5924), .Y(n16023) );
  AOI22XL U17894 ( .A0(B3_q[40]), .A1(n16158), .B0(B2_q[40]), .B1(n16143), .Y(
        n16024) );
  OAI211XL U17895 ( .A0(n5836), .A1(n15819), .B0(n15818), .C0(n15817), .Y(
        n15820) );
  AOI22XL U17896 ( .A0(B7_q[40]), .A1(n5930), .B0(B4_q[40]), .B1(n5925), .Y(
        n15818) );
  AOI21XL U17897 ( .A0(B6_q[40]), .A1(n15958), .B0(n28985), .Y(n15817) );
  AOI31XL U17898 ( .A0(cnt[10]), .A1(n11951), .A2(n28922), .B0(n11950), .Y(
        n5682) );
  OAI211XL U17899 ( .A0(n5799), .A1(n15758), .B0(n15369), .C0(n15368), .Y(
        n15370) );
  AOI21XL U17900 ( .A0(B4_q[4]), .A1(n7126), .B0(n28985), .Y(n15368) );
  AOI22XL U17901 ( .A0(B7_q[4]), .A1(n7127), .B0(B6_q[4]), .B1(n16570), .Y(
        n15369) );
  NAND4XL U17902 ( .A(n15363), .B(n15362), .C(n5800), .D(n15361), .Y(n15364)
         );
  NAND2XL U17903 ( .A(B4_q[5]), .B(n7126), .Y(n15363) );
  NAND2XL U17904 ( .A(B5_q[5]), .B(n16559), .Y(n15362) );
  NAND4XL U17905 ( .A(n15356), .B(n15355), .C(n5915), .D(n15354), .Y(n15357)
         );
  NAND2XL U17906 ( .A(B4_q[6]), .B(n7126), .Y(n15356) );
  NAND2XL U17907 ( .A(B5_q[6]), .B(n16559), .Y(n15355) );
  OAI211XL U17908 ( .A0(n15352), .A1(n5914), .B0(n15351), .C0(n15350), .Y(
        n15353) );
  AOI21XL U17909 ( .A0(B5_q[7]), .A1(n16559), .B0(n15349), .Y(n15350) );
  AOI22XL U17910 ( .A0(B7_q[7]), .A1(n7127), .B0(B6_q[7]), .B1(n16570), .Y(
        n15351) );
  INVXL U17911 ( .A(T1_rom3_q[13]), .Y(n29140) );
  OAI211XL U17912 ( .A0(n5799), .A1(n15980), .B0(n15383), .C0(n15382), .Y(
        n15384) );
  AOI21XL U17913 ( .A0(B4_q[1]), .A1(n7126), .B0(n5924), .Y(n15382) );
  AOI22XL U17914 ( .A0(B7_q[1]), .A1(n7127), .B0(B6_q[1]), .B1(n16570), .Y(
        n15383) );
  NAND4XL U17915 ( .A(n15380), .B(n15379), .C(n5910), .D(n15378), .Y(n15381)
         );
  NAND2XL U17916 ( .A(B6_q[2]), .B(n16570), .Y(n15380) );
  NAND2XL U17917 ( .A(B5_q[2]), .B(n16375), .Y(n15379) );
  OAI211XL U17918 ( .A0(n5799), .A1(n15972), .B0(n15376), .C0(n15375), .Y(
        n15377) );
  AOI21XL U17919 ( .A0(B7_q[3]), .A1(n16569), .B0(n16496), .Y(n15375) );
  AOI22XL U17920 ( .A0(B4_q[3]), .A1(n7126), .B0(B6_q[3]), .B1(n16570), .Y(
        n15376) );
  NAND2XL U17921 ( .A(n29112), .B(DATA0[0]), .Y(n5748) );
  NAND2XL U17922 ( .A(n29112), .B(DATA0[10]), .Y(n5738) );
  NAND2XL U17923 ( .A(n29112), .B(DATA0[12]), .Y(n5736) );
  NAND2XL U17924 ( .A(n29112), .B(DATA0[14]), .Y(n5734) );
  NAND2XL U17925 ( .A(n29112), .B(DATA0[15]), .Y(n5733) );
  NAND2XL U17926 ( .A(n29112), .B(DATA0[16]), .Y(n5732) );
  NAND2XL U17927 ( .A(n29112), .B(DATA0[17]), .Y(n5731) );
  NAND2XL U17928 ( .A(n29112), .B(DATA0[18]), .Y(n5730) );
  NAND2XL U17929 ( .A(n29112), .B(DATA0[20]), .Y(n5728) );
  NAND2XL U17930 ( .A(n29112), .B(DATA0[22]), .Y(n5726) );
  NAND2XL U17931 ( .A(n29112), .B(DATA0[24]), .Y(n5724) );
  NAND2XL U17932 ( .A(n29112), .B(DATA0[25]), .Y(n5723) );
  NAND2XL U17933 ( .A(n29112), .B(DATA0[26]), .Y(n5722) );
  NAND2XL U17934 ( .A(n29112), .B(DATA0[28]), .Y(n5720) );
  NAND2XL U17935 ( .A(n29112), .B(DATA0[2]), .Y(n5746) );
  NAND2XL U17936 ( .A(n29112), .B(DATA0[30]), .Y(n5718) );
  NAND2XL U17937 ( .A(n29112), .B(DATA0[32]), .Y(n5716) );
  NAND2XL U17938 ( .A(n29112), .B(DATA0[33]), .Y(n5715) );
  NAND2XL U17939 ( .A(n29112), .B(DATA0[34]), .Y(n5714) );
  NAND2XL U17940 ( .A(n29112), .B(DATA0[35]), .Y(n5713) );
  NAND2XL U17941 ( .A(n29112), .B(DATA0[36]), .Y(n5712) );
  NAND2XL U17942 ( .A(n29112), .B(DATA0[38]), .Y(n5710) );
  NAND2XL U17943 ( .A(n29112), .B(DATA0[40]), .Y(n5708) );
  NAND2XL U17944 ( .A(n29112), .B(DATA0[42]), .Y(n5706) );
  NAND2XL U17945 ( .A(n29112), .B(DATA0[43]), .Y(n5705) );
  NAND2XL U17946 ( .A(n29112), .B(DATA0[44]), .Y(n5704) );
  NAND2XL U17947 ( .A(n29112), .B(DATA0[46]), .Y(n5702) );
  NAND2XL U17948 ( .A(n29112), .B(DATA0[48]), .Y(n5700) );
  NAND2XL U17949 ( .A(n29112), .B(DATA0[4]), .Y(n5744) );
  NAND2XL U17950 ( .A(n29112), .B(DATA0[50]), .Y(n5698) );
  NAND2XL U17951 ( .A(n29112), .B(DATA0[51]), .Y(n5697) );
  NAND2XL U17952 ( .A(n29112), .B(DATA0[6]), .Y(n5742) );
  NAND2XL U17953 ( .A(n29112), .B(DATA0[7]), .Y(n5741) );
  NAND2XL U17954 ( .A(n29112), .B(DATA0[8]), .Y(n5740) );
  MXI2XL U17955 ( .A(n6914), .B(U1_pipe10[21]), .S0(n8053), .Y(n4859) );
  MXI2XL U17956 ( .A(n7637), .B(U1_pipe14[25]), .S0(n7096), .Y(n4776) );
  INVXL U17957 ( .A(n19400), .Y(n19095) );
  XOR2X1 U17958 ( .A(n17454), .B(n7012), .Y(n7661) );
  XNOR2X1 U17959 ( .A(n19079), .B(n19078), .Y(n19080) );
  NAND3XL U17960 ( .A(n17454), .B(n7654), .C(n9547), .Y(n7624) );
  OAI211XL U17961 ( .A0(n5799), .A1(n15819), .B0(n15304), .C0(n15303), .Y(
        n15305) );
  AOI21XL U17962 ( .A0(B6_q[40]), .A1(n16570), .B0(n5924), .Y(n15303) );
  AOI22XL U17963 ( .A0(B4_q[40]), .A1(n7126), .B0(B7_q[40]), .B1(n7127), .Y(
        n15304) );
  OAI211XL U17964 ( .A0(n15252), .A1(n5914), .B0(n15251), .C0(n15250), .Y(
        n15253) );
  AOI21XL U17965 ( .A0(B5_q[47]), .A1(n16375), .B0(n5924), .Y(n15250) );
  AOI22XL U17966 ( .A0(B7_q[47]), .A1(n7127), .B0(B6_q[47]), .B1(n16570), .Y(
        n15251) );
  OAI211XL U17967 ( .A0(n5914), .A1(n15268), .B0(n15267), .C0(n15266), .Y(
        n15269) );
  AOI21XL U17968 ( .A0(B6_q[45]), .A1(n16570), .B0(n15349), .Y(n15266) );
  AOI22XL U17969 ( .A0(B7_q[45]), .A1(n7127), .B0(B5_q[45]), .B1(n16559), .Y(
        n15267) );
  AOI22XL U17970 ( .A0(n12000), .A1(C_sel_reg[0]), .B0(C_sel_reg[2]), .B1(
        n5829), .Y(n5412) );
  NAND4XL U17971 ( .A(n15260), .B(n15259), .C(n5917), .D(n15258), .Y(n15261)
         );
  NAND2XL U17972 ( .A(B7_q[46]), .B(n16569), .Y(n15260) );
  NAND2XL U17973 ( .A(B5_q[46]), .B(n16559), .Y(n15259) );
  OAI211XL U17974 ( .A0(n5799), .A1(n15859), .B0(n15366), .C0(n15365), .Y(
        n15367) );
  AOI21XL U17975 ( .A0(B7_q[30]), .A1(n16569), .B0(n16496), .Y(n15365) );
  AOI22XL U17976 ( .A0(B4_q[30]), .A1(n7126), .B0(B6_q[30]), .B1(n16570), .Y(
        n15366) );
  INVXL U17977 ( .A(T1_rom3_q[11]), .Y(n29142) );
  OAI211XL U17978 ( .A0(n5799), .A1(n15815), .B0(n15297), .C0(n15296), .Y(
        n15298) );
  AOI21XL U17979 ( .A0(B6_q[41]), .A1(n16570), .B0(n5924), .Y(n15296) );
  AOI22XL U17980 ( .A0(B4_q[41]), .A1(n7126), .B0(B7_q[41]), .B1(n7127), .Y(
        n15297) );
  OAI211XL U17981 ( .A0(n5799), .A1(n15835), .B0(n15335), .C0(n15334), .Y(
        n15336) );
  AOI21XL U17982 ( .A0(B4_q[36]), .A1(n7126), .B0(n16496), .Y(n15334) );
  AOI22XL U17983 ( .A0(B7_q[36]), .A1(n7127), .B0(B6_q[36]), .B1(n16570), .Y(
        n15335) );
  INVXL U17984 ( .A(T1_rom3_q[7]), .Y(n29115) );
  INVXL U17985 ( .A(T1_rom2_q[15]), .Y(n29170) );
  OAI211XL U17986 ( .A0(n15967), .A1(n16168), .B0(n15221), .C0(n15220), .Y(
        n15222) );
  AOI22XL U17987 ( .A0(B2_q[0]), .A1(n15958), .B0(B1_q[0]), .B1(n15963), .Y(
        n15221) );
  AOI21XL U17988 ( .A0(B0_q[0]), .A1(n15969), .B0(n28985), .Y(n15220) );
  OAI211XL U17989 ( .A0(n16357), .A1(n5813), .B0(n16356), .C0(n16355), .Y(
        n16358) );
  AOI22XL U17990 ( .A0(B2_q[0]), .A1(n16354), .B0(B3_q[0]), .B1(n16325), .Y(
        n16356) );
  INVXL U17991 ( .A(B1_q[0]), .Y(n16357) );
  OAI211XL U17992 ( .A0(n5841), .A1(n16168), .B0(n16167), .C0(n16166), .Y(
        n16169) );
  AOI21XL U17993 ( .A0(B0_q[0]), .A1(n15557), .B0(n5924), .Y(n16166) );
  AOI22XL U17994 ( .A0(B2_q[0]), .A1(n16143), .B0(B1_q[0]), .B1(n16165), .Y(
        n16167) );
  OAI211XL U17995 ( .A0(n5914), .A1(n16573), .B0(n16572), .C0(n16571), .Y(
        n16574) );
  AOI22XL U17996 ( .A0(B1_q[0]), .A1(n16375), .B0(B2_q[0]), .B1(n16570), .Y(
        n16571) );
  OAI211XL U17997 ( .A0(n15967), .A1(n15185), .B0(n15184), .C0(n15183), .Y(
        n15186) );
  AOI22XL U17998 ( .A0(B1_q[10]), .A1(n15963), .B0(B0_q[10]), .B1(n5925), .Y(
        n15184) );
  OAI211XL U17999 ( .A0(n5813), .A1(n16531), .B0(n16315), .C0(n16314), .Y(
        n16316) );
  AOI21XL U18000 ( .A0(B3_q[10]), .A1(n16325), .B0(n5807), .Y(n16314) );
  AOI22XL U18001 ( .A0(B2_q[10]), .A1(n16354), .B0(B0_q[10]), .B1(n15687), .Y(
        n16315) );
  OAI211XL U18002 ( .A0(n5806), .A1(n16531), .B0(n16126), .C0(n16125), .Y(
        n16127) );
  AOI22XL U18003 ( .A0(B3_q[10]), .A1(n16158), .B0(B0_q[10]), .B1(n15557), .Y(
        n16126) );
  AOI21XL U18004 ( .A0(B2_q[10]), .A1(n16161), .B0(n28985), .Y(n16125) );
  OAI211XL U18005 ( .A0(n5799), .A1(n16531), .B0(n16530), .C0(n16529), .Y(
        n16532) );
  AOI21XL U18006 ( .A0(B0_q[10]), .A1(n7126), .B0(n16564), .Y(n16530) );
  AOI22XL U18007 ( .A0(B3_q[10]), .A1(n7127), .B0(B2_q[10]), .B1(n16570), .Y(
        n16529) );
  OAI211XL U18008 ( .A0(n5836), .A1(n16527), .B0(n15181), .C0(n15180), .Y(
        n15182) );
  AOI21XL U18009 ( .A0(B0_q[11]), .A1(n5925), .B0(n5924), .Y(n15180) );
  AOI22XL U18010 ( .A0(B2_q[11]), .A1(n15958), .B0(B3_q[11]), .B1(n15982), .Y(
        n15181) );
  OAI211XL U18011 ( .A0(n5813), .A1(n16527), .B0(n16312), .C0(n16311), .Y(
        n16313) );
  AOI21XL U18012 ( .A0(B2_q[11]), .A1(n5926), .B0(n5807), .Y(n16311) );
  AOI22XL U18013 ( .A0(B3_q[11]), .A1(n16325), .B0(B0_q[11]), .B1(n15687), .Y(
        n16312) );
  OAI211XL U18014 ( .A0(n5806), .A1(n16527), .B0(n16123), .C0(n16122), .Y(
        n16124) );
  AOI22XL U18015 ( .A0(B2_q[11]), .A1(n16143), .B0(B3_q[11]), .B1(n16128), .Y(
        n16123) );
  AOI21XL U18016 ( .A0(B0_q[11]), .A1(n15557), .B0(n28985), .Y(n16122) );
  OAI211XL U18017 ( .A0(n5799), .A1(n16527), .B0(n16526), .C0(n16525), .Y(
        n16528) );
  AOI21XL U18018 ( .A0(B0_q[11]), .A1(n7126), .B0(n28985), .Y(n16526) );
  AOI22XL U18019 ( .A0(B3_q[11]), .A1(n7127), .B0(B2_q[11]), .B1(n16570), .Y(
        n16525) );
  OAI211XL U18020 ( .A0(n15948), .A1(n15177), .B0(n15176), .C0(n15175), .Y(
        n15178) );
  AOI21XL U18021 ( .A0(B0_q[12]), .A1(n5925), .B0(n5924), .Y(n15175) );
  AOI22XL U18022 ( .A0(B1_q[12]), .A1(n15963), .B0(B3_q[12]), .B1(n15982), .Y(
        n15176) );
  OAI211XL U18023 ( .A0(n5813), .A1(n16523), .B0(n16309), .C0(n16308), .Y(
        n16310) );
  AOI21XL U18024 ( .A0(B0_q[12]), .A1(n15687), .B0(n5807), .Y(n16308) );
  AOI22XL U18025 ( .A0(B3_q[12]), .A1(n16325), .B0(B2_q[12]), .B1(n5926), .Y(
        n16309) );
  OAI211XL U18026 ( .A0(n5806), .A1(n16523), .B0(n16120), .C0(n16119), .Y(
        n16121) );
  AOI22XL U18027 ( .A0(B0_q[12]), .A1(n15557), .B0(B3_q[12]), .B1(n16128), .Y(
        n16120) );
  AOI21XL U18028 ( .A0(B2_q[12]), .A1(n16161), .B0(n28985), .Y(n16119) );
  OAI211XL U18029 ( .A0(n5799), .A1(n16523), .B0(n16522), .C0(n16521), .Y(
        n16524) );
  AOI21XL U18030 ( .A0(B2_q[12]), .A1(n16570), .B0(n28985), .Y(n16522) );
  AOI22XL U18031 ( .A0(B0_q[12]), .A1(n7126), .B0(B3_q[12]), .B1(n7127), .Y(
        n16521) );
  OAI211XL U18032 ( .A0(n15967), .A1(n15173), .B0(n15172), .C0(n15171), .Y(
        n15174) );
  AOI21XL U18033 ( .A0(B1_q[13]), .A1(n15963), .B0(n5924), .Y(n15171) );
  AOI22XL U18034 ( .A0(B0_q[13]), .A1(n5925), .B0(B2_q[13]), .B1(n15958), .Y(
        n15172) );
  OAI211XL U18035 ( .A0(n5813), .A1(n16519), .B0(n16306), .C0(n16305), .Y(
        n16307) );
  AOI21XL U18036 ( .A0(B3_q[13]), .A1(n16325), .B0(n5807), .Y(n16305) );
  AOI22XL U18037 ( .A0(B0_q[13]), .A1(n15687), .B0(B2_q[13]), .B1(n16354), .Y(
        n16306) );
  OAI211XL U18038 ( .A0(n5806), .A1(n16519), .B0(n16117), .C0(n16116), .Y(
        n16118) );
  AOI21XL U18039 ( .A0(B0_q[13]), .A1(n15557), .B0(n5924), .Y(n16116) );
  AOI22XL U18040 ( .A0(B2_q[13]), .A1(n16143), .B0(B3_q[13]), .B1(n16128), .Y(
        n16117) );
  OAI211XL U18041 ( .A0(n5799), .A1(n16519), .B0(n16518), .C0(n16517), .Y(
        n16520) );
  AOI21XL U18042 ( .A0(B3_q[13]), .A1(n7127), .B0(n5807), .Y(n16518) );
  AOI22XL U18043 ( .A0(B0_q[13]), .A1(n7126), .B0(B2_q[13]), .B1(n16570), .Y(
        n16517) );
  OAI211XL U18044 ( .A0(n5836), .A1(n16303), .B0(n15169), .C0(n15168), .Y(
        n15170) );
  AOI21XL U18045 ( .A0(B0_q[14]), .A1(n5925), .B0(n5924), .Y(n15168) );
  AOI22XL U18046 ( .A0(B3_q[14]), .A1(n15982), .B0(B2_q[14]), .B1(n15214), .Y(
        n15169) );
  OAI211XL U18047 ( .A0(n5813), .A1(n16303), .B0(n16302), .C0(n16301), .Y(
        n16304) );
  AOI21XL U18048 ( .A0(B0_q[14]), .A1(n15687), .B0(n5807), .Y(n16301) );
  AOI22XL U18049 ( .A0(B3_q[14]), .A1(n16325), .B0(B2_q[14]), .B1(n5926), .Y(
        n16302) );
  OAI211XL U18050 ( .A0(n5806), .A1(n16303), .B0(n16114), .C0(n16113), .Y(
        n16115) );
  AOI21XL U18051 ( .A0(B0_q[14]), .A1(n15557), .B0(n5924), .Y(n16113) );
  AOI22XL U18052 ( .A0(B3_q[14]), .A1(n16158), .B0(B2_q[14]), .B1(n16161), .Y(
        n16114) );
  OAI211XL U18053 ( .A0(n5914), .A1(n16515), .B0(n16514), .C0(n16513), .Y(
        n16516) );
  AOI21XL U18054 ( .A0(B1_q[14]), .A1(n16559), .B0(n28985), .Y(n16514) );
  AOI22XL U18055 ( .A0(B3_q[14]), .A1(n7127), .B0(B2_q[14]), .B1(n16570), .Y(
        n16513) );
  NAND3XL U18056 ( .A(n15166), .B(n15165), .C(n15164), .Y(n15167) );
  NAND2XL U18057 ( .A(B1_q[15]), .B(n15963), .Y(n15164) );
  AOI21XL U18058 ( .A0(B0_q[15]), .A1(n5925), .B0(n5924), .Y(n15165) );
  OAI211XL U18059 ( .A0(n15633), .A1(n16299), .B0(n16298), .C0(n16297), .Y(
        n16300) );
  AOI21XL U18060 ( .A0(B0_q[15]), .A1(n16277), .B0(n5807), .Y(n16297) );
  AOI22XL U18061 ( .A0(B3_q[15]), .A1(n16325), .B0(B1_q[15]), .B1(n16344), .Y(
        n16298) );
  OAI211XL U18062 ( .A0(n5806), .A1(n16111), .B0(n16110), .C0(n16109), .Y(
        n16112) );
  AOI21XL U18063 ( .A0(B0_q[15]), .A1(n5933), .B0(n16564), .Y(n16109) );
  AOI22XL U18064 ( .A0(B2_q[15]), .A1(n16143), .B0(B3_q[15]), .B1(n16128), .Y(
        n16110) );
  OAI211XL U18065 ( .A0(n5799), .A1(n16111), .B0(n16511), .C0(n16510), .Y(
        n16512) );
  AOI21XL U18066 ( .A0(B0_q[15]), .A1(n7126), .B0(n5924), .Y(n16511) );
  AOI22XL U18067 ( .A0(B3_q[15]), .A1(n7127), .B0(B2_q[15]), .B1(n16570), .Y(
        n16510) );
  OAI211XL U18068 ( .A0(n5813), .A1(n16508), .B0(n16295), .C0(n16294), .Y(
        n16296) );
  AOI21XL U18069 ( .A0(B3_q[16]), .A1(n16325), .B0(n5807), .Y(n16294) );
  AOI22XL U18070 ( .A0(B2_q[16]), .A1(n16293), .B0(B0_q[16]), .B1(n15687), .Y(
        n16295) );
  OAI211XL U18071 ( .A0(n5841), .A1(n16107), .B0(n16106), .C0(n16105), .Y(
        n16108) );
  AOI21XL U18072 ( .A0(B1_q[16]), .A1(n16165), .B0(n5807), .Y(n16105) );
  AOI22XL U18073 ( .A0(B2_q[16]), .A1(n16143), .B0(B0_q[16]), .B1(n15557), .Y(
        n16106) );
  OAI211XL U18074 ( .A0(n5799), .A1(n16508), .B0(n16507), .C0(n16506), .Y(
        n16509) );
  AOI21XL U18075 ( .A0(B0_q[16]), .A1(n7126), .B0(n5924), .Y(n16507) );
  AOI22XL U18076 ( .A0(B3_q[16]), .A1(n7127), .B0(B2_q[16]), .B1(n16570), .Y(
        n16506) );
  AOI21XL U18077 ( .A0(B0_q[17]), .A1(n5925), .B0(n15158), .Y(n15159) );
  NAND2XL U18078 ( .A(n6880), .B(n15157), .Y(n15158) );
  AOI21XL U18079 ( .A0(B2_q[17]), .A1(n5926), .B0(n16290), .Y(n16291) );
  NAND2XL U18080 ( .A(R7_valid), .B(n16289), .Y(n16290) );
  NAND4XL U18081 ( .A(n16103), .B(n16102), .C(n5906), .D(n16101), .Y(n16104)
         );
  NAND2XL U18082 ( .A(B3_q[17]), .B(n16158), .Y(n16103) );
  NAND2XL U18083 ( .A(B1_q[17]), .B(n16165), .Y(n16102) );
  OAI211XL U18084 ( .A0(n5799), .A1(n16504), .B0(n16503), .C0(n16502), .Y(
        n16505) );
  AOI21XL U18085 ( .A0(B0_q[17]), .A1(n7126), .B0(n16501), .Y(n16503) );
  AOI22XL U18086 ( .A0(B3_q[17]), .A1(n7127), .B0(B2_q[17]), .B1(n16570), .Y(
        n16502) );
  OAI211XL U18087 ( .A0(n15948), .A1(n16287), .B0(n15155), .C0(n15154), .Y(
        n15156) );
  AOI21XL U18088 ( .A0(B0_q[18]), .A1(n5925), .B0(n5924), .Y(n15154) );
  AOI22XL U18089 ( .A0(B3_q[18]), .A1(n5930), .B0(B1_q[18]), .B1(n15963), .Y(
        n15155) );
  OAI211XL U18090 ( .A0(n15633), .A1(n16287), .B0(n16286), .C0(n16285), .Y(
        n16288) );
  AOI21XL U18091 ( .A0(B0_q[18]), .A1(n15687), .B0(n5807), .Y(n16285) );
  AOI22XL U18092 ( .A0(B3_q[18]), .A1(n16325), .B0(B1_q[18]), .B1(n16344), .Y(
        n16286) );
  OAI211XL U18093 ( .A0(n5914), .A1(n16499), .B0(n16498), .C0(n16497), .Y(
        n16500) );
  AOI21XL U18094 ( .A0(B1_q[18]), .A1(n16559), .B0(n16496), .Y(n16498) );
  AOI22XL U18095 ( .A0(B3_q[18]), .A1(n7127), .B0(B2_q[18]), .B1(n16570), .Y(
        n16497) );
  OAI211XL U18096 ( .A0(n5813), .A1(n16494), .B0(n16283), .C0(n16282), .Y(
        n16284) );
  AOI21XL U18097 ( .A0(B3_q[19]), .A1(n16325), .B0(n5807), .Y(n16282) );
  AOI22XL U18098 ( .A0(B0_q[19]), .A1(n15687), .B0(B2_q[19]), .B1(n16354), .Y(
        n16283) );
  OAI2BB2XL U18099 ( .B0(n5915), .B1(AOPD[19]), .A0N(n16097), .A1N(n16096), 
        .Y(n3262) );
  AOI22XL U18100 ( .A0(B0_q[19]), .A1(n15557), .B0(B2_q[19]), .B1(n16143), .Y(
        n16096) );
  AOI21XL U18101 ( .A0(n16158), .A1(B3_q[19]), .B0(n16095), .Y(n16097) );
  OAI211XL U18102 ( .A0(n5799), .A1(n16494), .B0(n16493), .C0(n16492), .Y(
        n16495) );
  AOI21XL U18103 ( .A0(B2_q[19]), .A1(n16570), .B0(n5924), .Y(n16493) );
  AOI22XL U18104 ( .A0(B0_q[19]), .A1(n7126), .B0(B3_q[19]), .B1(n7127), .Y(
        n16492) );
  AOI21XL U18105 ( .A0(B0_q[1]), .A1(n5925), .B0(n15216), .Y(n15217) );
  NAND2XL U18106 ( .A(n6880), .B(n15215), .Y(n15216) );
  AOI21XL U18107 ( .A0(B3_q[1]), .A1(n16325), .B0(n16351), .Y(n16352) );
  NAND2XL U18108 ( .A(R7_valid), .B(n16350), .Y(n16351) );
  AOI21XL U18109 ( .A0(B2_q[1]), .A1(n16161), .B0(n16160), .Y(n16162) );
  NAND2XL U18110 ( .A(n6880), .B(n16159), .Y(n16160) );
  OAI211XL U18111 ( .A0(n5799), .A1(n16567), .B0(n16566), .C0(n16565), .Y(
        n16568) );
  AOI22XL U18112 ( .A0(B0_q[1]), .A1(n7126), .B0(B3_q[1]), .B1(n7127), .Y(
        n16565) );
  NAND4XL U18113 ( .A(n15149), .B(n15148), .C(n5913), .D(n15147), .Y(n15150)
         );
  NAND2XL U18114 ( .A(B1_q[20]), .B(n15963), .Y(n15149) );
  NAND2XL U18115 ( .A(B0_q[20]), .B(n5925), .Y(n15148) );
  NAND4XL U18116 ( .A(n16280), .B(n16279), .C(n5906), .D(n16278), .Y(n16281)
         );
  NAND2XL U18117 ( .A(B2_q[20]), .B(n16293), .Y(n16280) );
  NAND2XL U18118 ( .A(B0_q[20]), .B(n16277), .Y(n16279) );
  NAND4XL U18119 ( .A(n16093), .B(n16092), .C(n5906), .D(n16091), .Y(n16094)
         );
  NAND2XL U18120 ( .A(B3_q[20]), .B(n16158), .Y(n16093) );
  NAND2XL U18121 ( .A(B0_q[20]), .B(n15557), .Y(n16092) );
  OAI211XL U18122 ( .A0(n5914), .A1(n16490), .B0(n16489), .C0(n16488), .Y(
        n16491) );
  AOI22XL U18123 ( .A0(B3_q[20]), .A1(n7127), .B0(B2_q[20]), .B1(n16570), .Y(
        n16488) );
  OAI211XL U18124 ( .A0(n15967), .A1(n15145), .B0(n15144), .C0(n15143), .Y(
        n15146) );
  AOI21XL U18125 ( .A0(B1_q[21]), .A1(n15963), .B0(n5924), .Y(n15143) );
  AOI22XL U18126 ( .A0(B0_q[21]), .A1(n5925), .B0(B2_q[21]), .B1(n15958), .Y(
        n15144) );
  OAI211XL U18127 ( .A0(n5813), .A1(n16485), .B0(n16275), .C0(n16274), .Y(
        n16276) );
  AOI21XL U18128 ( .A0(B3_q[21]), .A1(n16325), .B0(n5807), .Y(n16274) );
  AOI22XL U18129 ( .A0(B0_q[21]), .A1(n15687), .B0(B2_q[21]), .B1(n16354), .Y(
        n16275) );
  OAI211XL U18130 ( .A0(n5806), .A1(n16485), .B0(n16089), .C0(n16088), .Y(
        n16090) );
  AOI21XL U18131 ( .A0(B2_q[21]), .A1(n16161), .B0(n28985), .Y(n16088) );
  AOI22XL U18132 ( .A0(B3_q[21]), .A1(n16158), .B0(B0_q[21]), .B1(n15557), .Y(
        n16089) );
  OAI211XL U18133 ( .A0(n5799), .A1(n16485), .B0(n16484), .C0(n16483), .Y(
        n16486) );
  AOI21XL U18134 ( .A0(B2_q[21]), .A1(n16570), .B0(n5924), .Y(n16484) );
  AOI22XL U18135 ( .A0(B0_q[21]), .A1(n7126), .B0(B3_q[21]), .B1(n7127), .Y(
        n16483) );
  OAI211XL U18136 ( .A0(n15967), .A1(n16086), .B0(n15141), .C0(n15140), .Y(
        n15142) );
  AOI21XL U18137 ( .A0(B1_q[22]), .A1(n15963), .B0(n5924), .Y(n15140) );
  AOI22XL U18138 ( .A0(B0_q[22]), .A1(n5925), .B0(B2_q[22]), .B1(n15958), .Y(
        n15141) );
  OAI211XL U18139 ( .A0(n5813), .A1(n16481), .B0(n16272), .C0(n16271), .Y(
        n16273) );
  AOI21XL U18140 ( .A0(B3_q[22]), .A1(n16325), .B0(n5924), .Y(n16271) );
  AOI22XL U18141 ( .A0(B0_q[22]), .A1(n15687), .B0(B2_q[22]), .B1(n16354), .Y(
        n16272) );
  OAI211XL U18142 ( .A0(n5841), .A1(n16086), .B0(n16085), .C0(n16084), .Y(
        n16087) );
  AOI21XL U18143 ( .A0(B1_q[22]), .A1(n16165), .B0(n28985), .Y(n16084) );
  AOI22XL U18144 ( .A0(B0_q[22]), .A1(n15557), .B0(B2_q[22]), .B1(n16161), .Y(
        n16085) );
  OAI211XL U18145 ( .A0(n14997), .A1(n16481), .B0(n16480), .C0(n16479), .Y(
        n16482) );
  AOI21XL U18146 ( .A0(B2_q[22]), .A1(n16570), .B0(n5924), .Y(n16480) );
  AOI22XL U18147 ( .A0(B0_q[22]), .A1(n7126), .B0(B3_q[22]), .B1(n7127), .Y(
        n16479) );
  OAI211XL U18148 ( .A0(n15967), .A1(n15138), .B0(n15137), .C0(n15136), .Y(
        n15139) );
  AOI21XL U18149 ( .A0(B1_q[23]), .A1(n15963), .B0(n5924), .Y(n15136) );
  AOI22XL U18150 ( .A0(B2_q[23]), .A1(n15958), .B0(B0_q[23]), .B1(n5925), .Y(
        n15137) );
  OAI211XL U18151 ( .A0(n16477), .A1(n5813), .B0(n16269), .C0(n16268), .Y(
        n16270) );
  AOI22XL U18152 ( .A0(B3_q[23]), .A1(n16325), .B0(B2_q[23]), .B1(n16354), .Y(
        n16269) );
  AOI21XL U18153 ( .A0(B0_q[23]), .A1(n15687), .B0(n28985), .Y(n16268) );
  OAI211XL U18154 ( .A0(n5806), .A1(n16477), .B0(n16082), .C0(n16081), .Y(
        n16083) );
  AOI22XL U18155 ( .A0(B3_q[23]), .A1(n16158), .B0(B2_q[23]), .B1(n16143), .Y(
        n16082) );
  AOI21XL U18156 ( .A0(B0_q[23]), .A1(n15557), .B0(n28985), .Y(n16081) );
  OAI211XL U18157 ( .A0(n5799), .A1(n16477), .B0(n16476), .C0(n16475), .Y(
        n16478) );
  AOI21XL U18158 ( .A0(B0_q[23]), .A1(n7126), .B0(n5924), .Y(n16476) );
  AOI22XL U18159 ( .A0(B3_q[23]), .A1(n7127), .B0(B2_q[23]), .B1(n16570), .Y(
        n16475) );
  OAI2BB2XL U18160 ( .B0(n5909), .B1(AOPB[24]), .A0N(n15135), .A1N(n15134), 
        .Y(n3284) );
  AOI22XL U18161 ( .A0(B0_q[24]), .A1(n5925), .B0(B2_q[24]), .B1(n15958), .Y(
        n15134) );
  AOI21XL U18162 ( .A0(n5930), .A1(B3_q[24]), .B0(n15133), .Y(n15135) );
  OAI211XL U18163 ( .A0(n5813), .A1(n16473), .B0(n16266), .C0(n16265), .Y(
        n16267) );
  AOI22XL U18164 ( .A0(B0_q[24]), .A1(n15687), .B0(B2_q[24]), .B1(n16354), .Y(
        n16266) );
  AOI21XL U18165 ( .A0(B3_q[24]), .A1(n16325), .B0(n28985), .Y(n16265) );
  OAI211XL U18166 ( .A0(n5806), .A1(n16473), .B0(n16079), .C0(n16078), .Y(
        n16080) );
  AOI22XL U18167 ( .A0(B3_q[24]), .A1(n16128), .B0(B0_q[24]), .B1(n15557), .Y(
        n16079) );
  AOI21XL U18168 ( .A0(B2_q[24]), .A1(n16161), .B0(n28985), .Y(n16078) );
  OAI211XL U18169 ( .A0(n5799), .A1(n16473), .B0(n16472), .C0(n16471), .Y(
        n16474) );
  AOI21XL U18170 ( .A0(B2_q[24]), .A1(n16570), .B0(n16470), .Y(n16472) );
  AOI22XL U18171 ( .A0(B0_q[24]), .A1(n7126), .B0(B3_q[24]), .B1(n7127), .Y(
        n16471) );
  OAI2BB2XL U18172 ( .B0(n5909), .B1(AOPB[25]), .A0N(n15132), .A1N(n15131), 
        .Y(n3288) );
  AOI22XL U18173 ( .A0(B3_q[25]), .A1(n5930), .B0(B2_q[25]), .B1(n15958), .Y(
        n15131) );
  AOI21XL U18174 ( .A0(n15963), .A1(B1_q[25]), .B0(n15130), .Y(n15132) );
  OAI211XL U18175 ( .A0(n16348), .A1(n16263), .B0(n16262), .C0(n16261), .Y(
        n16264) );
  AOI21XL U18176 ( .A0(B0_q[25]), .A1(n15687), .B0(n5924), .Y(n16261) );
  AOI22XL U18177 ( .A0(B1_q[25]), .A1(n16344), .B0(B2_q[25]), .B1(n16354), .Y(
        n16262) );
  OAI2BB2XL U18178 ( .B0(n5909), .B1(AOPD[25]), .A0N(n16077), .A1N(n16076), 
        .Y(n3290) );
  AOI22XL U18179 ( .A0(B3_q[25]), .A1(n16158), .B0(B2_q[25]), .B1(n16143), .Y(
        n16076) );
  AOI21XL U18180 ( .A0(n5931), .A1(B1_q[25]), .B0(n16075), .Y(n16077) );
  OAI211XL U18181 ( .A0(n5914), .A1(n16468), .B0(n16467), .C0(n16466), .Y(
        n16469) );
  AOI21XL U18182 ( .A0(B2_q[25]), .A1(n16570), .B0(n28985), .Y(n16467) );
  AOI22XL U18183 ( .A0(B3_q[25]), .A1(n7127), .B0(B1_q[25]), .B1(n16559), .Y(
        n16466) );
  OAI211XL U18184 ( .A0(n16348), .A1(n16259), .B0(n16258), .C0(n16257), .Y(
        n16260) );
  AOI21XL U18185 ( .A0(B0_q[26]), .A1(n15687), .B0(n5924), .Y(n16257) );
  AOI22XL U18186 ( .A0(B2_q[26]), .A1(n16354), .B0(B1_q[26]), .B1(n16344), .Y(
        n16258) );
  OAI211XL U18187 ( .A0(n5841), .A1(n16259), .B0(n16073), .C0(n16072), .Y(
        n16074) );
  AOI21XL U18188 ( .A0(B0_q[26]), .A1(n15557), .B0(n16487), .Y(n16072) );
  AOI22XL U18189 ( .A0(B2_q[26]), .A1(n16143), .B0(B1_q[26]), .B1(n16165), .Y(
        n16073) );
  AOI21XL U18190 ( .A0(B1_q[26]), .A1(n16559), .B0(n16461), .Y(n16463) );
  AOI22XL U18191 ( .A0(B3_q[26]), .A1(n7127), .B0(B2_q[26]), .B1(n16570), .Y(
        n16462) );
  NAND4XL U18192 ( .A(n16255), .B(n16254), .C(n5910), .D(n16253), .Y(n16256)
         );
  NAND2XL U18193 ( .A(B2_q[27]), .B(n16293), .Y(n16255) );
  NAND2XL U18194 ( .A(B0_q[27]), .B(n16277), .Y(n16254) );
  AOI21XL U18195 ( .A0(B0_q[27]), .A1(n5933), .B0(n16069), .Y(n16070) );
  NAND2XL U18196 ( .A(R7_valid), .B(n16068), .Y(n16069) );
  OAI211XL U18197 ( .A0(n14997), .A1(n16459), .B0(n16458), .C0(n16457), .Y(
        n16460) );
  AOI21XL U18198 ( .A0(B0_q[27]), .A1(n7126), .B0(n5924), .Y(n16458) );
  AOI22XL U18199 ( .A0(B3_q[27]), .A1(n7127), .B0(B2_q[27]), .B1(n16570), .Y(
        n16457) );
  OAI211XL U18200 ( .A0(n15967), .A1(n16251), .B0(n15119), .C0(n15118), .Y(
        n15120) );
  AOI21XL U18201 ( .A0(B2_q[28]), .A1(n15958), .B0(n5924), .Y(n15118) );
  AOI22XL U18202 ( .A0(B0_q[28]), .A1(n5925), .B0(B1_q[28]), .B1(n15963), .Y(
        n15119) );
  OAI211XL U18203 ( .A0(n16348), .A1(n16251), .B0(n16250), .C0(n16249), .Y(
        n16252) );
  AOI21XL U18204 ( .A0(B0_q[28]), .A1(n15687), .B0(n5924), .Y(n16249) );
  AOI22XL U18205 ( .A0(B2_q[28]), .A1(n16354), .B0(B1_q[28]), .B1(n16344), .Y(
        n16250) );
  OAI211XL U18206 ( .A0(n5841), .A1(n16251), .B0(n16066), .C0(n16065), .Y(
        n16067) );
  AOI21XL U18207 ( .A0(B0_q[28]), .A1(n5933), .B0(n5924), .Y(n16065) );
  AOI22XL U18208 ( .A0(B2_q[28]), .A1(n16161), .B0(B1_q[28]), .B1(n16165), .Y(
        n16066) );
  OAI211XL U18209 ( .A0(n5914), .A1(n16455), .B0(n16454), .C0(n16453), .Y(
        n16456) );
  AOI21XL U18210 ( .A0(B3_q[28]), .A1(n7127), .B0(n5924), .Y(n16454) );
  AOI22XL U18211 ( .A0(B1_q[28]), .A1(n16375), .B0(B2_q[28]), .B1(n16570), .Y(
        n16453) );
  AOI22XL U18212 ( .A0(B3_q[29]), .A1(n15982), .B0(B2_q[29]), .B1(n15958), .Y(
        n15116) );
  AOI21XL U18213 ( .A0(n15963), .A1(B1_q[29]), .B0(n15115), .Y(n15117) );
  AOI22XL U18214 ( .A0(B3_q[29]), .A1(n16325), .B0(B2_q[29]), .B1(n5926), .Y(
        n16247) );
  AOI21XL U18215 ( .A0(n15747), .A1(B1_q[29]), .B0(n16246), .Y(n16248) );
  OAI211XL U18216 ( .A0(n16063), .A1(n15495), .B0(n16062), .C0(n16061), .Y(
        n16064) );
  AOI21XL U18217 ( .A0(B0_q[29]), .A1(n5933), .B0(n5924), .Y(n16061) );
  AOI22XL U18218 ( .A0(B3_q[29]), .A1(n16158), .B0(B1_q[29]), .B1(n16165), .Y(
        n16062) );
  OAI211XL U18219 ( .A0(n5914), .A1(n16451), .B0(n16450), .C0(n16449), .Y(
        n16452) );
  AOI21XL U18220 ( .A0(B2_q[29]), .A1(n16570), .B0(n16470), .Y(n16450) );
  AOI22XL U18221 ( .A0(B3_q[29]), .A1(n7127), .B0(B1_q[29]), .B1(n16559), .Y(
        n16449) );
  OAI211XL U18222 ( .A0(n15948), .A1(n15212), .B0(n15211), .C0(n15210), .Y(
        n15213) );
  AOI21XL U18223 ( .A0(B0_q[2]), .A1(n5925), .B0(n15349), .Y(n15210) );
  AOI22XL U18224 ( .A0(B3_q[2]), .A1(n5930), .B0(B1_q[2]), .B1(n15963), .Y(
        n15211) );
  OAI211XL U18225 ( .A0(n16348), .A1(n16347), .B0(n16346), .C0(n16345), .Y(
        n16349) );
  AOI21XL U18226 ( .A0(B0_q[2]), .A1(n15687), .B0(n5924), .Y(n16345) );
  AOI22XL U18227 ( .A0(B2_q[2]), .A1(n16354), .B0(B1_q[2]), .B1(n16344), .Y(
        n16346) );
  AOI22XL U18228 ( .A0(B2_q[2]), .A1(n16143), .B0(B1_q[2]), .B1(n16165), .Y(
        n16156) );
  AOI21XL U18229 ( .A0(n16158), .A1(B3_q[2]), .B0(n16155), .Y(n16157) );
  OAI211XL U18230 ( .A0(n5914), .A1(n16562), .B0(n16561), .C0(n16560), .Y(
        n16563) );
  AOI21XL U18231 ( .A0(B1_q[2]), .A1(n16559), .B0(n5924), .Y(n16561) );
  AOI22XL U18232 ( .A0(B3_q[2]), .A1(n7127), .B0(B2_q[2]), .B1(n16570), .Y(
        n16560) );
  OAI211XL U18233 ( .A0(n5799), .A1(n16447), .B0(n16446), .C0(n16445), .Y(
        n16448) );
  AOI21XL U18234 ( .A0(B0_q[30]), .A1(n7126), .B0(n5924), .Y(n16446) );
  AOI22XL U18235 ( .A0(B3_q[30]), .A1(n7127), .B0(B2_q[30]), .B1(n16570), .Y(
        n16445) );
  OAI211XL U18236 ( .A0(n5914), .A1(n16443), .B0(n16442), .C0(n16441), .Y(
        n16444) );
  AOI21XL U18237 ( .A0(B2_q[31]), .A1(n16570), .B0(n16501), .Y(n16442) );
  AOI22XL U18238 ( .A0(B3_q[31]), .A1(n7127), .B0(B1_q[31]), .B1(n16559), .Y(
        n16441) );
  AOI21XL U18239 ( .A0(B3_q[32]), .A1(n16325), .B0(n16235), .Y(n16236) );
  NAND2XL U18240 ( .A(n6880), .B(n16234), .Y(n16235) );
  OAI211XL U18241 ( .A0(n5799), .A1(n16439), .B0(n16438), .C0(n16437), .Y(
        n16440) );
  AOI21XL U18242 ( .A0(B0_q[32]), .A1(n7126), .B0(n5924), .Y(n16438) );
  AOI22XL U18243 ( .A0(B3_q[32]), .A1(n7127), .B0(B2_q[32]), .B1(n16570), .Y(
        n16437) );
  OAI211XL U18244 ( .A0(n5799), .A1(n16435), .B0(n16434), .C0(n16433), .Y(
        n16436) );
  AOI21XL U18245 ( .A0(B3_q[33]), .A1(n7127), .B0(n5924), .Y(n16434) );
  AOI22XL U18246 ( .A0(B0_q[33]), .A1(n7126), .B0(B2_q[33]), .B1(n16570), .Y(
        n16433) );
  OAI211XL U18247 ( .A0(n15218), .A1(n16431), .B0(n15099), .C0(n15098), .Y(
        n15100) );
  AOI21XL U18248 ( .A0(B0_q[34]), .A1(n5925), .B0(n5924), .Y(n15098) );
  AOI22XL U18249 ( .A0(B3_q[34]), .A1(n15982), .B0(B2_q[34]), .B1(n15958), .Y(
        n15099) );
  OAI211XL U18250 ( .A0(n5813), .A1(n16431), .B0(n16229), .C0(n16228), .Y(
        n16230) );
  AOI21XL U18251 ( .A0(B2_q[34]), .A1(n5926), .B0(n5924), .Y(n16228) );
  AOI22XL U18252 ( .A0(B3_q[34]), .A1(n16325), .B0(B0_q[34]), .B1(n15687), .Y(
        n16229) );
  OAI211XL U18253 ( .A0(n5806), .A1(n16431), .B0(n16044), .C0(n16043), .Y(
        n16045) );
  AOI21XL U18254 ( .A0(B0_q[34]), .A1(n15557), .B0(n5924), .Y(n16043) );
  AOI22XL U18255 ( .A0(B3_q[34]), .A1(n16158), .B0(B2_q[34]), .B1(n16161), .Y(
        n16044) );
  OAI211XL U18256 ( .A0(n5799), .A1(n16431), .B0(n16430), .C0(n16429), .Y(
        n16432) );
  AOI21XL U18257 ( .A0(B0_q[34]), .A1(n7126), .B0(n5924), .Y(n16430) );
  AOI22XL U18258 ( .A0(B3_q[34]), .A1(n7127), .B0(B2_q[34]), .B1(n16570), .Y(
        n16429) );
  AOI22XL U18259 ( .A0(B1_q[35]), .A1(n16165), .B0(B3_q[35]), .B1(n16128), .Y(
        n16041) );
  AOI21XL U18260 ( .A0(n16161), .A1(B2_q[35]), .B0(n16040), .Y(n16042) );
  OAI211XL U18261 ( .A0(n5914), .A1(n16427), .B0(n16426), .C0(n16425), .Y(
        n16428) );
  AOI21XL U18262 ( .A0(B2_q[35]), .A1(n16570), .B0(n5924), .Y(n16426) );
  AOI22XL U18263 ( .A0(B3_q[35]), .A1(n7127), .B0(B1_q[35]), .B1(n16559), .Y(
        n16425) );
  NAND4XL U18264 ( .A(n15093), .B(n15092), .C(n5910), .D(n15091), .Y(n15094)
         );
  NAND2XL U18265 ( .A(B1_q[36]), .B(n15963), .Y(n15093) );
  NAND2XL U18266 ( .A(B0_q[36]), .B(n15969), .Y(n15092) );
  NAND4XL U18267 ( .A(n16222), .B(n16221), .C(n5912), .D(n16220), .Y(n16223)
         );
  NAND2XL U18268 ( .A(B3_q[36]), .B(n16325), .Y(n16222) );
  NAND2XL U18269 ( .A(B0_q[36]), .B(n16277), .Y(n16221) );
  NAND4XL U18270 ( .A(n16038), .B(n16037), .C(n5909), .D(n16036), .Y(n16039)
         );
  NAND2XL U18271 ( .A(B2_q[36]), .B(n16143), .Y(n16038) );
  NAND2XL U18272 ( .A(B0_q[36]), .B(n15557), .Y(n16037) );
  OAI211XL U18273 ( .A0(n5914), .A1(n16423), .B0(n16422), .C0(n16421), .Y(
        n16424) );
  AOI21XL U18274 ( .A0(B1_q[36]), .A1(n16559), .B0(n5924), .Y(n16422) );
  AOI22XL U18275 ( .A0(B3_q[36]), .A1(n7127), .B0(B2_q[36]), .B1(n16570), .Y(
        n16421) );
  AOI22XL U18276 ( .A0(B3_q[37]), .A1(n15982), .B0(B2_q[37]), .B1(n15958), .Y(
        n15089) );
  AOI21XL U18277 ( .A0(n15963), .A1(B1_q[37]), .B0(n15088), .Y(n15090) );
  AOI22XL U18278 ( .A0(B3_q[37]), .A1(n16325), .B0(B2_q[37]), .B1(n16354), .Y(
        n16218) );
  AOI21XL U18279 ( .A0(n15747), .A1(B1_q[37]), .B0(n16217), .Y(n16219) );
  OAI211XL U18280 ( .A0(n5914), .A1(n16419), .B0(n16418), .C0(n16417), .Y(
        n16420) );
  AOI21XL U18281 ( .A0(B2_q[37]), .A1(n16570), .B0(n5924), .Y(n16418) );
  AOI22XL U18282 ( .A0(B3_q[37]), .A1(n7127), .B0(B1_q[37]), .B1(n16559), .Y(
        n16417) );
  AOI22XL U18283 ( .A0(B2_q[38]), .A1(n15958), .B0(B3_q[38]), .B1(n5930), .Y(
        n15086) );
  AOI21XL U18284 ( .A0(n15963), .A1(B1_q[38]), .B0(n15085), .Y(n15087) );
  AOI22XL U18285 ( .A0(B2_q[38]), .A1(n16143), .B0(B3_q[38]), .B1(n16128), .Y(
        n16030) );
  AOI21XL U18286 ( .A0(n5931), .A1(B1_q[38]), .B0(n16029), .Y(n16031) );
  AOI21XL U18287 ( .A0(B1_q[38]), .A1(n16559), .B0(n28985), .Y(n16413) );
  AOI22XL U18288 ( .A0(B3_q[38]), .A1(n7127), .B0(B2_q[38]), .B1(n16570), .Y(
        n16412) );
  AOI22XL U18289 ( .A0(B2_q[39]), .A1(n15958), .B0(B0_q[39]), .B1(n5925), .Y(
        n15083) );
  AOI21XL U18290 ( .A0(n15982), .A1(B3_q[39]), .B0(n15082), .Y(n15084) );
  AOI22XL U18291 ( .A0(B2_q[39]), .A1(n16143), .B0(B0_q[39]), .B1(n15557), .Y(
        n16027) );
  AOI21XL U18292 ( .A0(n16136), .A1(B3_q[39]), .B0(n16026), .Y(n16028) );
  OAI211XL U18293 ( .A0(n5799), .A1(n16410), .B0(n16409), .C0(n16408), .Y(
        n16411) );
  AOI21XL U18294 ( .A0(B0_q[39]), .A1(n7126), .B0(n28985), .Y(n16409) );
  AOI22XL U18295 ( .A0(B3_q[39]), .A1(n7127), .B0(B2_q[39]), .B1(n16570), .Y(
        n16408) );
  OAI211XL U18296 ( .A0(n15948), .A1(n15208), .B0(n15207), .C0(n15206), .Y(
        n15209) );
  AOI21XL U18297 ( .A0(B0_q[3]), .A1(n5925), .B0(n28985), .Y(n15206) );
  AOI22XL U18298 ( .A0(B1_q[3]), .A1(n15963), .B0(B3_q[3]), .B1(n5930), .Y(
        n15207) );
  OAI211XL U18299 ( .A0(n5813), .A1(n16342), .B0(n16341), .C0(n16340), .Y(
        n16343) );
  AOI22XL U18300 ( .A0(B3_q[3]), .A1(n16325), .B0(B2_q[3]), .B1(n16354), .Y(
        n16341) );
  AOI21XL U18301 ( .A0(B0_q[3]), .A1(n15687), .B0(n28985), .Y(n16340) );
  OAI211XL U18302 ( .A0(n5806), .A1(n16342), .B0(n16152), .C0(n16151), .Y(
        n16153) );
  AOI21XL U18303 ( .A0(B0_q[3]), .A1(n5933), .B0(n5924), .Y(n16151) );
  AOI22XL U18304 ( .A0(B3_q[3]), .A1(n16158), .B0(B2_q[3]), .B1(n16143), .Y(
        n16152) );
  OAI211XL U18305 ( .A0(n5799), .A1(n16342), .B0(n16557), .C0(n16556), .Y(
        n16558) );
  AOI21XL U18306 ( .A0(B2_q[3]), .A1(n16570), .B0(n28985), .Y(n16557) );
  AOI22XL U18307 ( .A0(B0_q[3]), .A1(n7126), .B0(B3_q[3]), .B1(n7127), .Y(
        n16556) );
  OAI211XL U18308 ( .A0(n15218), .A1(n16406), .B0(n15080), .C0(n15079), .Y(
        n15081) );
  AOI21XL U18309 ( .A0(B2_q[40]), .A1(n15958), .B0(n5924), .Y(n15079) );
  AOI22XL U18310 ( .A0(B3_q[40]), .A1(n15982), .B0(B0_q[40]), .B1(n5925), .Y(
        n15080) );
  OAI211XL U18311 ( .A0(n5813), .A1(n16406), .B0(n16208), .C0(n16207), .Y(
        n16209) );
  AOI21XL U18312 ( .A0(B0_q[40]), .A1(n15687), .B0(n5924), .Y(n16207) );
  AOI22XL U18313 ( .A0(B3_q[40]), .A1(n16325), .B0(B2_q[40]), .B1(n16354), .Y(
        n16208) );
  OAI211XL U18314 ( .A0(n5799), .A1(n16406), .B0(n16405), .C0(n16404), .Y(
        n16407) );
  AOI21XL U18315 ( .A0(B0_q[40]), .A1(n7126), .B0(n28985), .Y(n16405) );
  AOI22XL U18316 ( .A0(B3_q[40]), .A1(n7127), .B0(B2_q[40]), .B1(n16570), .Y(
        n16404) );
  OAI211XL U18317 ( .A0(n16348), .A1(n16205), .B0(n16204), .C0(n16203), .Y(
        n16206) );
  AOI22XL U18318 ( .A0(B2_q[41]), .A1(n5926), .B0(B1_q[41]), .B1(n16344), .Y(
        n16204) );
  OAI211XL U18319 ( .A0(n5841), .A1(n16205), .B0(n16021), .C0(n16020), .Y(
        n16022) );
  AOI21XL U18320 ( .A0(B0_q[41]), .A1(n5933), .B0(n16496), .Y(n16020) );
  AOI22XL U18321 ( .A0(B2_q[41]), .A1(n16143), .B0(B1_q[41]), .B1(n16165), .Y(
        n16021) );
  AOI21XL U18322 ( .A0(B1_q[41]), .A1(n16559), .B0(n5924), .Y(n16401) );
  AOI22XL U18323 ( .A0(B3_q[41]), .A1(n7127), .B0(B2_q[41]), .B1(n16570), .Y(
        n16400) );
  OAI211XL U18324 ( .A0(n5836), .A1(n16398), .B0(n15074), .C0(n15073), .Y(
        n15075) );
  AOI21XL U18325 ( .A0(B0_q[42]), .A1(n5925), .B0(n5924), .Y(n15073) );
  AOI22XL U18326 ( .A0(B2_q[42]), .A1(n15958), .B0(B3_q[42]), .B1(n5930), .Y(
        n15074) );
  OAI211XL U18327 ( .A0(n5813), .A1(n16398), .B0(n16201), .C0(n16200), .Y(
        n16202) );
  AOI21XL U18328 ( .A0(B0_q[42]), .A1(n15687), .B0(n28985), .Y(n16200) );
  AOI22XL U18329 ( .A0(B2_q[42]), .A1(n5926), .B0(B3_q[42]), .B1(n16325), .Y(
        n16201) );
  OAI211XL U18330 ( .A0(n5806), .A1(n16398), .B0(n16018), .C0(n16017), .Y(
        n16019) );
  AOI21XL U18331 ( .A0(B2_q[42]), .A1(n16161), .B0(n5924), .Y(n16017) );
  AOI22XL U18332 ( .A0(B0_q[42]), .A1(n15557), .B0(B3_q[42]), .B1(n16128), .Y(
        n16018) );
  OAI211XL U18333 ( .A0(n5799), .A1(n16398), .B0(n16397), .C0(n16396), .Y(
        n16399) );
  AOI22XL U18334 ( .A0(B0_q[42]), .A1(n7126), .B0(B2_q[42]), .B1(n16570), .Y(
        n16396) );
  NAND4XL U18335 ( .A(n15071), .B(n15070), .C(n5912), .D(n15069), .Y(n15072)
         );
  NAND2XL U18336 ( .A(B3_q[43]), .B(n15982), .Y(n15071) );
  NAND2XL U18337 ( .A(B0_q[43]), .B(n15969), .Y(n15070) );
  NAND4XL U18338 ( .A(n16198), .B(n16197), .C(n5907), .D(n16196), .Y(n16199)
         );
  NAND2XL U18339 ( .A(B1_q[43]), .B(n16344), .Y(n16198) );
  NAND2XL U18340 ( .A(B0_q[43]), .B(n15687), .Y(n16197) );
  NAND4XL U18341 ( .A(n16015), .B(n16014), .C(n5908), .D(n16013), .Y(n16016)
         );
  NAND2XL U18342 ( .A(B2_q[43]), .B(n16143), .Y(n16015) );
  NAND2XL U18343 ( .A(B0_q[43]), .B(n15557), .Y(n16014) );
  AOI21XL U18344 ( .A0(B1_q[43]), .A1(n16559), .B0(n28985), .Y(n16393) );
  AOI22XL U18345 ( .A0(B3_q[43]), .A1(n7127), .B0(B2_q[43]), .B1(n16570), .Y(
        n16392) );
  OAI211XL U18346 ( .A0(n5836), .A1(n16390), .B0(n15067), .C0(n15066), .Y(
        n15068) );
  AOI21XL U18347 ( .A0(B0_q[44]), .A1(n5925), .B0(n5924), .Y(n15066) );
  AOI22XL U18348 ( .A0(B2_q[44]), .A1(n15958), .B0(B3_q[44]), .B1(n15982), .Y(
        n15067) );
  OAI211XL U18349 ( .A0(n5813), .A1(n16390), .B0(n16194), .C0(n16193), .Y(
        n16195) );
  AOI21XL U18350 ( .A0(B3_q[44]), .A1(n16325), .B0(n5924), .Y(n16193) );
  AOI22XL U18351 ( .A0(B0_q[44]), .A1(n15687), .B0(B2_q[44]), .B1(n16354), .Y(
        n16194) );
  OAI211XL U18352 ( .A0(n5799), .A1(n16390), .B0(n16389), .C0(n16388), .Y(
        n16391) );
  AOI21XL U18353 ( .A0(B3_q[44]), .A1(n7127), .B0(n5807), .Y(n16389) );
  AOI22XL U18354 ( .A0(B0_q[44]), .A1(n7126), .B0(B2_q[44]), .B1(n16570), .Y(
        n16388) );
  OAI211XL U18355 ( .A0(n15967), .A1(n16191), .B0(n15064), .C0(n15063), .Y(
        n15065) );
  AOI21XL U18356 ( .A0(B1_q[45]), .A1(n15963), .B0(n16496), .Y(n15063) );
  AOI22XL U18357 ( .A0(B2_q[45]), .A1(n15958), .B0(B0_q[45]), .B1(n5925), .Y(
        n15064) );
  OAI211XL U18358 ( .A0(n16348), .A1(n16191), .B0(n16190), .C0(n16189), .Y(
        n16192) );
  AOI21XL U18359 ( .A0(B0_q[45]), .A1(n15687), .B0(n5924), .Y(n16189) );
  AOI22XL U18360 ( .A0(B2_q[45]), .A1(n16354), .B0(B1_q[45]), .B1(n16344), .Y(
        n16190) );
  OAI2BB2XL U18361 ( .B0(n5915), .B1(AOPD[45]), .A0N(n16009), .A1N(n16008), 
        .Y(n3378) );
  AOI22XL U18362 ( .A0(B2_q[45]), .A1(n16143), .B0(B3_q[45]), .B1(n16128), .Y(
        n16008) );
  AOI21XL U18363 ( .A0(n5931), .A1(B1_q[45]), .B0(n16007), .Y(n16009) );
  AOI21XL U18364 ( .A0(B1_q[45]), .A1(n16559), .B0(n5807), .Y(n16385) );
  AOI22XL U18365 ( .A0(B3_q[45]), .A1(n7127), .B0(B2_q[45]), .B1(n16570), .Y(
        n16384) );
  AOI21XL U18366 ( .A0(B0_q[46]), .A1(n5925), .B0(n15060), .Y(n15061) );
  NAND2XL U18367 ( .A(R7_valid), .B(n15059), .Y(n15060) );
  AOI21XL U18368 ( .A0(B2_q[46]), .A1(n5926), .B0(n16186), .Y(n16187) );
  NAND2XL U18369 ( .A(n6880), .B(n16185), .Y(n16186) );
  NAND4XL U18370 ( .A(n16005), .B(n16004), .C(R7_valid), .D(n16003), .Y(n16006) );
  NAND2XL U18371 ( .A(B3_q[46]), .B(n16158), .Y(n16005) );
  NAND2XL U18372 ( .A(B1_q[46]), .B(n16165), .Y(n16004) );
  OAI211XL U18373 ( .A0(n14997), .A1(n16382), .B0(n16381), .C0(n16380), .Y(
        n16383) );
  AOI21XL U18374 ( .A0(B3_q[46]), .A1(n7127), .B0(n5807), .Y(n16381) );
  AOI22XL U18375 ( .A0(B0_q[46]), .A1(n7126), .B0(B2_q[46]), .B1(n16570), .Y(
        n16380) );
  AOI22XL U18376 ( .A0(B2_q[47]), .A1(n15958), .B0(B0_q[47]), .B1(n5925), .Y(
        n15057) );
  OAI211XL U18377 ( .A0(n5813), .A1(n16378), .B0(n16183), .C0(n16182), .Y(
        n16184) );
  AOI21XL U18378 ( .A0(B3_q[47]), .A1(n16325), .B0(n5924), .Y(n16182) );
  AOI22XL U18379 ( .A0(B2_q[47]), .A1(n16354), .B0(B0_q[47]), .B1(n15687), .Y(
        n16183) );
  OAI211XL U18380 ( .A0(n5806), .A1(n16378), .B0(n16001), .C0(n16000), .Y(
        n16002) );
  AOI21XL U18381 ( .A0(B0_q[47]), .A1(n15557), .B0(n16496), .Y(n16000) );
  AOI22XL U18382 ( .A0(B2_q[47]), .A1(n16143), .B0(B3_q[47]), .B1(n16128), .Y(
        n16001) );
  OAI211XL U18383 ( .A0(n5799), .A1(n16378), .B0(n16377), .C0(n16376), .Y(
        n16379) );
  AOI21XL U18384 ( .A0(B3_q[47]), .A1(n7127), .B0(n5807), .Y(n16377) );
  AOI22XL U18385 ( .A0(B0_q[47]), .A1(n7126), .B0(B2_q[47]), .B1(n16570), .Y(
        n16376) );
  OAI211XL U18386 ( .A0(n15054), .A1(n15967), .B0(n15053), .C0(n15052), .Y(
        n15055) );
  AOI21XL U18387 ( .A0(B1_q[48]), .A1(n15963), .B0(n5924), .Y(n15052) );
  AOI22XL U18388 ( .A0(B2_q[48]), .A1(n15958), .B0(B0_q[48]), .B1(n5925), .Y(
        n15053) );
  OAI211XL U18389 ( .A0(n16373), .A1(n5813), .B0(n16180), .C0(n16179), .Y(
        n16181) );
  AOI21XL U18390 ( .A0(B0_q[48]), .A1(n15687), .B0(n5924), .Y(n16179) );
  AOI22XL U18391 ( .A0(B2_q[48]), .A1(n16354), .B0(B3_q[48]), .B1(n16325), .Y(
        n16180) );
  OAI211XL U18392 ( .A0(n5806), .A1(n16373), .B0(n15998), .C0(n15997), .Y(
        n15999) );
  AOI21XL U18393 ( .A0(B0_q[48]), .A1(n5933), .B0(n16496), .Y(n15997) );
  AOI22XL U18394 ( .A0(B2_q[48]), .A1(n16143), .B0(B3_q[48]), .B1(n16128), .Y(
        n15998) );
  OAI211XL U18395 ( .A0(n5799), .A1(n16373), .B0(n16372), .C0(n16371), .Y(
        n16374) );
  AOI21XL U18396 ( .A0(B0_q[48]), .A1(n7126), .B0(n5807), .Y(n16372) );
  AOI22XL U18397 ( .A0(B3_q[48]), .A1(n7127), .B0(B2_q[48]), .B1(n16570), .Y(
        n16371) );
  OAI211XL U18398 ( .A0(n5836), .A1(n16369), .B0(n15050), .C0(n15049), .Y(
        n15051) );
  AOI21XL U18399 ( .A0(B0_q[49]), .A1(n5925), .B0(n5924), .Y(n15049) );
  AOI22XL U18400 ( .A0(B2_q[49]), .A1(n15958), .B0(B3_q[49]), .B1(n15982), .Y(
        n15050) );
  OAI211XL U18401 ( .A0(n16369), .A1(n5813), .B0(n16177), .C0(n16176), .Y(
        n16178) );
  AOI21XL U18402 ( .A0(B0_q[49]), .A1(n15687), .B0(n28985), .Y(n16176) );
  AOI22XL U18403 ( .A0(B2_q[49]), .A1(n16354), .B0(B3_q[49]), .B1(n16325), .Y(
        n16177) );
  OAI211XL U18404 ( .A0(n5841), .A1(n15995), .B0(n15994), .C0(n15993), .Y(
        n15996) );
  AOI21XL U18405 ( .A0(B1_q[49]), .A1(n16165), .B0(n5924), .Y(n15993) );
  AOI22XL U18406 ( .A0(B0_q[49]), .A1(n15557), .B0(B2_q[49]), .B1(n16143), .Y(
        n15994) );
  OAI211XL U18407 ( .A0(n5799), .A1(n16369), .B0(n16368), .C0(n16367), .Y(
        n16370) );
  AOI21XL U18408 ( .A0(B3_q[49]), .A1(n7127), .B0(n5924), .Y(n16368) );
  AOI22XL U18409 ( .A0(B0_q[49]), .A1(n7126), .B0(B2_q[49]), .B1(n16570), .Y(
        n16367) );
  OAI211XL U18410 ( .A0(n15967), .A1(n16338), .B0(n15204), .C0(n15203), .Y(
        n15205) );
  AOI21XL U18411 ( .A0(B0_q[4]), .A1(n5925), .B0(n5924), .Y(n15203) );
  AOI22XL U18412 ( .A0(B2_q[4]), .A1(n15958), .B0(B1_q[4]), .B1(n15963), .Y(
        n15204) );
  OAI211XL U18413 ( .A0(n16348), .A1(n16338), .B0(n16337), .C0(n16336), .Y(
        n16339) );
  AOI22XL U18414 ( .A0(B2_q[4]), .A1(n16354), .B0(B1_q[4]), .B1(n16344), .Y(
        n16337) );
  AOI21XL U18415 ( .A0(B0_q[4]), .A1(n15687), .B0(n28985), .Y(n16336) );
  OAI211XL U18416 ( .A0(n15495), .A1(n16149), .B0(n16148), .C0(n16147), .Y(
        n16150) );
  AOI21XL U18417 ( .A0(B0_q[4]), .A1(n5933), .B0(n5924), .Y(n16147) );
  AOI22XL U18418 ( .A0(B3_q[4]), .A1(n16158), .B0(B1_q[4]), .B1(n16165), .Y(
        n16148) );
  OAI211XL U18419 ( .A0(n5914), .A1(n16554), .B0(n16553), .C0(n16552), .Y(
        n16555) );
  AOI21XL U18420 ( .A0(B1_q[4]), .A1(n16559), .B0(n5924), .Y(n16553) );
  AOI22XL U18421 ( .A0(B3_q[4]), .A1(n7127), .B0(B2_q[4]), .B1(n16570), .Y(
        n16552) );
  OAI211XL U18422 ( .A0(n15967), .A1(n15047), .B0(n15046), .C0(n15045), .Y(
        n15048) );
  AOI21XL U18423 ( .A0(B1_q[50]), .A1(n15963), .B0(n5924), .Y(n15045) );
  AOI22XL U18424 ( .A0(B2_q[50]), .A1(n15958), .B0(B0_q[50]), .B1(n5925), .Y(
        n15046) );
  OAI211XL U18425 ( .A0(n5813), .A1(n16365), .B0(n16174), .C0(n16173), .Y(
        n16175) );
  AOI21XL U18426 ( .A0(B3_q[50]), .A1(n16325), .B0(n5924), .Y(n16173) );
  AOI22XL U18427 ( .A0(B2_q[50]), .A1(n16354), .B0(B0_q[50]), .B1(n15687), .Y(
        n16174) );
  OAI211XL U18428 ( .A0(n5806), .A1(n16365), .B0(n15991), .C0(n15990), .Y(
        n15992) );
  AOI21XL U18429 ( .A0(B2_q[50]), .A1(n16161), .B0(n16496), .Y(n15990) );
  AOI22XL U18430 ( .A0(B3_q[50]), .A1(n16158), .B0(B0_q[50]), .B1(n15557), .Y(
        n15991) );
  OAI211XL U18431 ( .A0(n5799), .A1(n16365), .B0(n16364), .C0(n16363), .Y(
        n16366) );
  AOI21XL U18432 ( .A0(B0_q[50]), .A1(n7126), .B0(n5924), .Y(n16364) );
  AOI22XL U18433 ( .A0(B3_q[50]), .A1(n7127), .B0(B2_q[50]), .B1(n16570), .Y(
        n16363) );
  OAI211XL U18434 ( .A0(n15043), .A1(n15948), .B0(n15042), .C0(n15041), .Y(
        n15044) );
  AOI21XL U18435 ( .A0(B0_q[51]), .A1(n5925), .B0(n5924), .Y(n15041) );
  AOI22XL U18436 ( .A0(B3_q[51]), .A1(n15982), .B0(B1_q[51]), .B1(n15963), .Y(
        n15042) );
  OAI2BB2XL U18437 ( .B0(n5915), .B1(AOPC[51]), .A0N(n16172), .A1N(n16171), 
        .Y(n3405) );
  AOI22XL U18438 ( .A0(B2_q[51]), .A1(n5926), .B0(B1_q[51]), .B1(n16344), .Y(
        n16171) );
  AOI21XL U18439 ( .A0(n16325), .A1(B3_q[51]), .B0(n16170), .Y(n16172) );
  OAI2BB2XL U18440 ( .B0(n5915), .B1(AOPD[51]), .A0N(n15989), .A1N(n15988), 
        .Y(n3406) );
  AOI22XL U18441 ( .A0(B2_q[51]), .A1(n16143), .B0(B1_q[51]), .B1(n16165), .Y(
        n15988) );
  AOI21XL U18442 ( .A0(n16136), .A1(B3_q[51]), .B0(n15987), .Y(n15989) );
  AOI21XL U18443 ( .A0(B1_q[51]), .A1(n16559), .B0(n5924), .Y(n16360) );
  AOI22XL U18444 ( .A0(B3_q[51]), .A1(n7127), .B0(B2_q[51]), .B1(n16570), .Y(
        n16359) );
  OAI211XL U18445 ( .A0(n5836), .A1(n16550), .B0(n15201), .C0(n15200), .Y(
        n15202) );
  AOI21XL U18446 ( .A0(B2_q[5]), .A1(n15958), .B0(n5924), .Y(n15200) );
  AOI22XL U18447 ( .A0(B3_q[5]), .A1(n15982), .B0(B0_q[5]), .B1(n5925), .Y(
        n15201) );
  OAI211XL U18448 ( .A0(n5813), .A1(n16550), .B0(n16334), .C0(n16333), .Y(
        n16335) );
  AOI21XL U18449 ( .A0(B0_q[5]), .A1(n15687), .B0(n5807), .Y(n16333) );
  AOI22XL U18450 ( .A0(B3_q[5]), .A1(n16325), .B0(B2_q[5]), .B1(n16354), .Y(
        n16334) );
  OAI211XL U18451 ( .A0(n5806), .A1(n16550), .B0(n16145), .C0(n16144), .Y(
        n16146) );
  AOI21XL U18452 ( .A0(B0_q[5]), .A1(n15557), .B0(n5924), .Y(n16144) );
  AOI22XL U18453 ( .A0(B3_q[5]), .A1(n16158), .B0(B2_q[5]), .B1(n16143), .Y(
        n16145) );
  OAI211XL U18454 ( .A0(n5799), .A1(n16550), .B0(n16549), .C0(n16548), .Y(
        n16551) );
  AOI21XL U18455 ( .A0(B0_q[5]), .A1(n7126), .B0(n16496), .Y(n16549) );
  AOI22XL U18456 ( .A0(B3_q[5]), .A1(n7127), .B0(B2_q[5]), .B1(n16570), .Y(
        n16548) );
  OAI211XL U18457 ( .A0(n15948), .A1(n16331), .B0(n15198), .C0(n15197), .Y(
        n15199) );
  AOI21XL U18458 ( .A0(B0_q[6]), .A1(n5925), .B0(n5924), .Y(n15197) );
  AOI22XL U18459 ( .A0(B3_q[6]), .A1(n15982), .B0(B1_q[6]), .B1(n15963), .Y(
        n15198) );
  OAI211XL U18460 ( .A0(n15633), .A1(n16331), .B0(n16330), .C0(n16329), .Y(
        n16332) );
  AOI21XL U18461 ( .A0(B0_q[6]), .A1(n15687), .B0(n5807), .Y(n16329) );
  AOI22XL U18462 ( .A0(B3_q[6]), .A1(n16325), .B0(B1_q[6]), .B1(n16344), .Y(
        n16330) );
  OAI211XL U18463 ( .A0(n5806), .A1(n16141), .B0(n16140), .C0(n16139), .Y(
        n16142) );
  AOI22XL U18464 ( .A0(B3_q[6]), .A1(n16158), .B0(B2_q[6]), .B1(n16143), .Y(
        n16140) );
  AOI21XL U18465 ( .A0(B0_q[6]), .A1(n5933), .B0(n28985), .Y(n16139) );
  OAI211XL U18466 ( .A0(n5799), .A1(n16141), .B0(n16546), .C0(n16545), .Y(
        n16547) );
  AOI21XL U18467 ( .A0(B0_q[6]), .A1(n7126), .B0(n5924), .Y(n16546) );
  AOI22XL U18468 ( .A0(B3_q[6]), .A1(n7127), .B0(B2_q[6]), .B1(n16570), .Y(
        n16545) );
  OAI211XL U18469 ( .A0(n5813), .A1(n16543), .B0(n16327), .C0(n16326), .Y(
        n16328) );
  AOI21XL U18470 ( .A0(B3_q[7]), .A1(n16325), .B0(n5807), .Y(n16326) );
  AOI22XL U18471 ( .A0(B2_q[7]), .A1(n16354), .B0(B0_q[7]), .B1(n15687), .Y(
        n16327) );
  OAI211XL U18472 ( .A0(n5799), .A1(n16543), .B0(n16542), .C0(n16541), .Y(
        n16544) );
  AOI21XL U18473 ( .A0(B0_q[7]), .A1(n7126), .B0(n5807), .Y(n16542) );
  AOI22XL U18474 ( .A0(B3_q[7]), .A1(n7127), .B0(B2_q[7]), .B1(n16570), .Y(
        n16541) );
  OAI211XL U18475 ( .A0(n5836), .A1(n16323), .B0(n15192), .C0(n15191), .Y(
        n15193) );
  AOI21XL U18476 ( .A0(B0_q[8]), .A1(n5925), .B0(n5924), .Y(n15191) );
  AOI22XL U18477 ( .A0(B3_q[8]), .A1(n15982), .B0(B2_q[8]), .B1(n15958), .Y(
        n15192) );
  OAI211XL U18478 ( .A0(n5813), .A1(n16323), .B0(n16322), .C0(n16321), .Y(
        n16324) );
  AOI21XL U18479 ( .A0(B0_q[8]), .A1(n15687), .B0(n5807), .Y(n16321) );
  AOI22XL U18480 ( .A0(B3_q[8]), .A1(n16325), .B0(B2_q[8]), .B1(n16354), .Y(
        n16322) );
  OAI211XL U18481 ( .A0(n5806), .A1(n16323), .B0(n16133), .C0(n16132), .Y(
        n16134) );
  AOI22XL U18482 ( .A0(B3_q[8]), .A1(n16158), .B0(B2_q[8]), .B1(n16143), .Y(
        n16133) );
  AOI21XL U18483 ( .A0(B0_q[8]), .A1(n15557), .B0(n28985), .Y(n16132) );
  OAI211XL U18484 ( .A0(n5914), .A1(n16539), .B0(n16538), .C0(n16537), .Y(
        n16540) );
  AOI21XL U18485 ( .A0(B2_q[8]), .A1(n16570), .B0(n5924), .Y(n16538) );
  AOI22XL U18486 ( .A0(B3_q[8]), .A1(n7127), .B0(B1_q[8]), .B1(n16559), .Y(
        n16537) );
  OAI211XL U18487 ( .A0(n15967), .A1(n15189), .B0(n15188), .C0(n15187), .Y(
        n15190) );
  AOI22XL U18488 ( .A0(B1_q[9]), .A1(n15963), .B0(B2_q[9]), .B1(n15958), .Y(
        n15188) );
  OAI211XL U18489 ( .A0(n5813), .A1(n16319), .B0(n16318), .C0(n16317), .Y(
        n16320) );
  AOI21XL U18490 ( .A0(B0_q[9]), .A1(n15687), .B0(n5807), .Y(n16317) );
  AOI22XL U18491 ( .A0(B2_q[9]), .A1(n16354), .B0(B3_q[9]), .B1(n16325), .Y(
        n16318) );
  OAI211XL U18492 ( .A0(n5806), .A1(n16319), .B0(n16130), .C0(n16129), .Y(
        n16131) );
  AOI22XL U18493 ( .A0(B2_q[9]), .A1(n16143), .B0(B3_q[9]), .B1(n16128), .Y(
        n16130) );
  AOI21XL U18494 ( .A0(B0_q[9]), .A1(n15557), .B0(n28985), .Y(n16129) );
  OAI211XL U18495 ( .A0(n5914), .A1(n16535), .B0(n16534), .C0(n16533), .Y(
        n16536) );
  AOI21XL U18496 ( .A0(B3_q[9]), .A1(n7127), .B0(n5924), .Y(n16534) );
  AOI22XL U18497 ( .A0(B1_q[9]), .A1(n16375), .B0(B2_q[9]), .B1(n16570), .Y(
        n16533) );
  MXI2XL U18498 ( .A(Q0[30]), .B(n25871), .S0(n24128), .Y(n3428) );
  XNOR2XL U18499 ( .A(n25961), .B(n25870), .Y(n25871) );
  NAND2XL U18500 ( .A(n25907), .B(n25959), .Y(n25870) );
  XOR2XL U18501 ( .A(n28689), .B(n28993), .Y(n27062) );
  XOR2XL U18502 ( .A(n27059), .B(n27019), .Y(n27020) );
  NAND2XL U18503 ( .A(n27018), .B(n27057), .Y(n27019) );
  INVXL U18504 ( .A(n27058), .Y(n27018) );
  MXI2XL U18505 ( .A(Q0[51]), .B(n26977), .S0(n24128), .Y(n3431) );
  XNOR2XL U18506 ( .A(n27015), .B(n26976), .Y(n26977) );
  NAND2XL U18507 ( .A(n26973), .B(n27013), .Y(n26976) );
  MXI2XL U18508 ( .A(Q0[50]), .B(n26937), .S0(n23239), .Y(n3432) );
  XOR2XL U18509 ( .A(n26972), .B(n26936), .Y(n26937) );
  NAND2XL U18510 ( .A(n26935), .B(n26970), .Y(n26936) );
  INVXL U18511 ( .A(n26971), .Y(n26935) );
  MXI2XL U18512 ( .A(Q0[49]), .B(n26895), .S0(n23239), .Y(n3433) );
  XNOR2XL U18513 ( .A(n26932), .B(n26894), .Y(n26895) );
  NAND2XL U18514 ( .A(n26891), .B(n26930), .Y(n26894) );
  MXI2XL U18515 ( .A(Q0[48]), .B(n26850), .S0(n23239), .Y(n3434) );
  XOR2XL U18516 ( .A(n26890), .B(n26849), .Y(n26850) );
  NAND2XL U18517 ( .A(n26848), .B(n26888), .Y(n26849) );
  INVXL U18518 ( .A(n26889), .Y(n26848) );
  MXI2XL U18519 ( .A(Q0[47]), .B(n26802), .S0(n24128), .Y(n3435) );
  MXI2XL U18520 ( .A(Q0[46]), .B(n26741), .S0(n24128), .Y(n3436) );
  XOR2XL U18521 ( .A(n26740), .B(n26739), .Y(n26741) );
  NAND2XL U18522 ( .A(n26736), .B(n26792), .Y(n26739) );
  MXI2XL U18523 ( .A(Q0[45]), .B(n26686), .S0(n24128), .Y(n3437) );
  XOR2XL U18524 ( .A(n26685), .B(n26684), .Y(n26686) );
  NAND2XL U18525 ( .A(n26683), .B(n26732), .Y(n26684) );
  AOI21XL U18526 ( .A0(n26735), .A1(n26680), .B0(n26679), .Y(n26685) );
  MXI2XL U18527 ( .A(Q0[44]), .B(n26635), .S0(n23239), .Y(n3438) );
  XOR2XL U18528 ( .A(n26634), .B(n26633), .Y(n26635) );
  NAND2XL U18529 ( .A(n26630), .B(n26676), .Y(n26633) );
  AOI21XL U18530 ( .A0(n26735), .A1(n26675), .B0(n26678), .Y(n26634) );
  MXI2XL U18531 ( .A(Q0[43]), .B(n26570), .S0(n24128), .Y(n3439) );
  XOR2XL U18532 ( .A(n26569), .B(n26568), .Y(n26570) );
  NAND2XL U18533 ( .A(n26567), .B(n26627), .Y(n26568) );
  AOI21XL U18534 ( .A0(n26735), .A1(n26564), .B0(n26563), .Y(n26569) );
  MXI2XL U18535 ( .A(Q0[42]), .B(n26502), .S0(n24128), .Y(n3440) );
  XNOR2XL U18536 ( .A(n26735), .B(n26501), .Y(n26502) );
  NAND2XL U18537 ( .A(n26564), .B(n26628), .Y(n26501) );
  MXI2XL U18538 ( .A(Q0[41]), .B(n26441), .S0(n23239), .Y(n3441) );
  XOR2XL U18539 ( .A(n26440), .B(n26439), .Y(n26441) );
  NAND2XL U18540 ( .A(n26438), .B(n26487), .Y(n26439) );
  AOI21XL U18541 ( .A0(n26435), .A1(n26434), .B0(n26433), .Y(n26440) );
  MXI2XL U18542 ( .A(Q0[40]), .B(n26390), .S0(n23239), .Y(n3442) );
  XNOR2XL U18543 ( .A(n26435), .B(n26389), .Y(n26390) );
  NAND2XL U18544 ( .A(n26434), .B(n26488), .Y(n26389) );
  MXI2XL U18545 ( .A(Q0[39]), .B(n26332), .S0(n23239), .Y(n3443) );
  XOR2XL U18546 ( .A(n26331), .B(n26330), .Y(n26332) );
  NAND2XL U18547 ( .A(n26329), .B(n26381), .Y(n26330) );
  AOI21XL U18548 ( .A0(n26326), .A1(n26325), .B0(n26324), .Y(n26331) );
  MXI2XL U18549 ( .A(Q0[38]), .B(n26268), .S0(n24128), .Y(n3444) );
  XOR2XL U18550 ( .A(n26386), .B(n26267), .Y(n26268) );
  NAND2XL U18551 ( .A(n26325), .B(n26382), .Y(n26267) );
  MXI2XL U18552 ( .A(Q0[37]), .B(n26214), .S0(n23239), .Y(n3445) );
  XOR2XL U18553 ( .A(n26213), .B(n26212), .Y(n26214) );
  NAND2XL U18554 ( .A(n26211), .B(n26258), .Y(n26212) );
  AOI21XL U18555 ( .A0(n26208), .A1(n26207), .B0(n26206), .Y(n26213) );
  MXI2XL U18556 ( .A(Q0[36]), .B(n26175), .S0(n23239), .Y(n3446) );
  XNOR2XL U18557 ( .A(n26208), .B(n26174), .Y(n26175) );
  NAND2XL U18558 ( .A(n26207), .B(n26259), .Y(n26174) );
  MXI2XL U18559 ( .A(Q0[35]), .B(n26109), .S0(n24128), .Y(n3447) );
  XNOR2XL U18560 ( .A(n26108), .B(n26107), .Y(n26109) );
  NAND2XL U18561 ( .A(n26106), .B(n26167), .Y(n26107) );
  MXI2XL U18562 ( .A(Q0[34]), .B(n26064), .S0(U1_valid[1]), .Y(n3448) );
  XOR2XL U18563 ( .A(n26264), .B(n26063), .Y(n26064) );
  NAND2XL U18564 ( .A(n26062), .B(n26168), .Y(n26063) );
  INVXL U18565 ( .A(n26166), .Y(n26062) );
  MXI2XL U18566 ( .A(Q0[33]), .B(n26009), .S0(U1_valid[1]), .Y(n3449) );
  XNOR2XL U18567 ( .A(n26008), .B(n26007), .Y(n26009) );
  NAND2XL U18568 ( .A(n26006), .B(n26051), .Y(n26007) );
  MXI2XL U18569 ( .A(Q0[32]), .B(n25966), .S0(U1_valid[1]), .Y(n3450) );
  INVXL U18570 ( .A(n26049), .Y(n25964) );
  MXI2XL U18571 ( .A(Q0[31]), .B(n25913), .S0(n23559), .Y(n3451) );
  XOR2XL U18572 ( .A(n25912), .B(n25911), .Y(n25913) );
  NAND2XL U18573 ( .A(n25910), .B(n25958), .Y(n25911) );
  MXI2XL U18574 ( .A(Q0[29]), .B(n25820), .S0(n24128), .Y(n3452) );
  XNOR2XL U18575 ( .A(n25819), .B(n25818), .Y(n25820) );
  NAND2XL U18576 ( .A(n25817), .B(n25862), .Y(n25818) );
  MXI2XL U18577 ( .A(Q2[40]), .B(n26399), .S0(n24128), .Y(n3453) );
  XOR2XL U18578 ( .A(n26398), .B(n26397), .Y(n26399) );
  NAND2XL U18579 ( .A(n26396), .B(n26443), .Y(n26397) );
  AOI21XL U18580 ( .A0(n26393), .A1(n26392), .B0(n26391), .Y(n26398) );
  MXI2XL U18581 ( .A(Q2[39]), .B(n26323), .S0(n23239), .Y(n3454) );
  XOR2XL U18582 ( .A(n26448), .B(n26322), .Y(n26323) );
  NAND2XL U18583 ( .A(n26392), .B(n26444), .Y(n26322) );
  MXI2XL U18584 ( .A(Q2[38]), .B(n26286), .S0(n24128), .Y(n3455) );
  XOR2XL U18585 ( .A(n26285), .B(n26284), .Y(n26286) );
  NAND2XL U18586 ( .A(n26283), .B(n26313), .Y(n26284) );
  AOI21XL U18587 ( .A0(n26280), .A1(n26279), .B0(n26278), .Y(n26285) );
  MXI2XL U18588 ( .A(Q2[37]), .B(n26234), .S0(n24128), .Y(n3456) );
  XNOR2XL U18589 ( .A(n26280), .B(n26233), .Y(n26234) );
  NAND2XL U18590 ( .A(n26279), .B(n26314), .Y(n26233) );
  MXI2XL U18591 ( .A(Q2[36]), .B(n26165), .S0(n24128), .Y(n3457) );
  XNOR2XL U18592 ( .A(n26164), .B(n26163), .Y(n26165) );
  NAND2XL U18593 ( .A(n26162), .B(n26226), .Y(n26163) );
  MXI2XL U18594 ( .A(Q2[35]), .B(n26141), .S0(n23239), .Y(n3458) );
  XOR2XL U18595 ( .A(n26319), .B(n26140), .Y(n26141) );
  NAND2XL U18596 ( .A(n26139), .B(n26227), .Y(n26140) );
  INVXL U18597 ( .A(n26225), .Y(n26139) );
  MXI2XL U18598 ( .A(Q2[34]), .B(n26048), .S0(n18739), .Y(n3459) );
  XNOR2XL U18599 ( .A(n26047), .B(n26046), .Y(n26048) );
  NAND2XL U18600 ( .A(n26045), .B(n26128), .Y(n26046) );
  MXI2XL U18601 ( .A(Q2[33]), .B(n26002), .S0(n18351), .Y(n3460) );
  XOR2XL U18602 ( .A(n26042), .B(n26001), .Y(n26002) );
  NAND2XL U18603 ( .A(n26000), .B(n26129), .Y(n26001) );
  INVXL U18604 ( .A(n26126), .Y(n26000) );
  MXI2XL U18605 ( .A(Q2[32]), .B(n25982), .S0(n18893), .Y(n3461) );
  XOR2XL U18606 ( .A(n25981), .B(n25980), .Y(n25982) );
  NAND2XL U18607 ( .A(n25979), .B(n25994), .Y(n25980) );
  AOI21XL U18608 ( .A0(n25997), .A1(n25976), .B0(n25975), .Y(n25981) );
  MXI2XL U18609 ( .A(Q2[31]), .B(n25935), .S0(n24128), .Y(n3462) );
  XNOR2XL U18610 ( .A(n25997), .B(n25934), .Y(n25935) );
  NAND2XL U18611 ( .A(n25976), .B(n25995), .Y(n25934) );
  MXI2XL U18612 ( .A(Q2[30]), .B(n25885), .S0(n23239), .Y(n3463) );
  XNOR2XL U18613 ( .A(n25884), .B(n25883), .Y(n25885) );
  NAND2XL U18614 ( .A(n25882), .B(n25926), .Y(n25883) );
  MXI2XL U18615 ( .A(Q2[29]), .B(n25813), .S0(n24128), .Y(n3464) );
  XOR2XL U18616 ( .A(n25879), .B(n25812), .Y(n25813) );
  NAND2XL U18617 ( .A(n25811), .B(n25927), .Y(n25812) );
  INVXL U18618 ( .A(n25925), .Y(n25811) );
  MXI2XL U18619 ( .A(Q2[28]), .B(n24859), .S0(n23239), .Y(n3465) );
  NAND2XL U18620 ( .A(n24854), .B(n25806), .Y(n24858) );
  INVXL U18621 ( .A(n25807), .Y(n24854) );
  XOR2XL U18622 ( .A(n28691), .B(n28995), .Y(n24407) );
  XOR2XL U18623 ( .A(n24404), .B(n24352), .Y(n24353) );
  NAND2XL U18624 ( .A(n24351), .B(n24402), .Y(n24352) );
  INVXL U18625 ( .A(n24403), .Y(n24351) );
  MXI2XL U18626 ( .A(Q1[23]), .B(n24310), .S0(n23239), .Y(n3468) );
  XNOR2XL U18627 ( .A(n24348), .B(n24309), .Y(n24310) );
  NAND2XL U18628 ( .A(n24306), .B(n24346), .Y(n24309) );
  MXI2XL U18629 ( .A(Q1[22]), .B(n24285), .S0(n23239), .Y(n3469) );
  XOR2XL U18630 ( .A(n24305), .B(n24284), .Y(n24285) );
  NAND2XL U18631 ( .A(n24283), .B(n24303), .Y(n24284) );
  INVXL U18632 ( .A(n24304), .Y(n24283) );
  MXI2XL U18633 ( .A(Q1[21]), .B(n24243), .S0(n23239), .Y(n3470) );
  XNOR2XL U18634 ( .A(n24280), .B(n24242), .Y(n24243) );
  NAND2XL U18635 ( .A(n24239), .B(n24278), .Y(n24242) );
  MXI2XL U18636 ( .A(Q1[20]), .B(n24198), .S0(n23239), .Y(n3471) );
  XOR2XL U18637 ( .A(n24238), .B(n24197), .Y(n24198) );
  NAND2XL U18638 ( .A(n24196), .B(n24236), .Y(n24197) );
  INVXL U18639 ( .A(n24237), .Y(n24196) );
  MXI2XL U18640 ( .A(Q1[19]), .B(n24129), .S0(n24128), .Y(n3472) );
  XNOR2XL U18641 ( .A(n24193), .B(n24127), .Y(n24129) );
  NAND2XL U18642 ( .A(n24124), .B(n24191), .Y(n24127) );
  MXI2XL U18643 ( .A(Q1[18]), .B(n24090), .S0(n24128), .Y(n3473) );
  XOR2XL U18644 ( .A(n24089), .B(n24088), .Y(n24090) );
  NAND2XL U18645 ( .A(n24085), .B(n24118), .Y(n24088) );
  MXI2XL U18646 ( .A(Q1[17]), .B(n24011), .S0(n24128), .Y(n3474) );
  XOR2XL U18647 ( .A(n24010), .B(n24009), .Y(n24011) );
  NAND2XL U18648 ( .A(n24008), .B(n24081), .Y(n24009) );
  AOI21XL U18649 ( .A0(n24084), .A1(n24005), .B0(n24004), .Y(n24010) );
  MXI2XL U18650 ( .A(Q1[16]), .B(n23978), .S0(n24128), .Y(n3475) );
  XOR2XL U18651 ( .A(n23977), .B(n23976), .Y(n23978) );
  NAND2XL U18652 ( .A(n23973), .B(n24001), .Y(n23976) );
  AOI21XL U18653 ( .A0(n24084), .A1(n24000), .B0(n24003), .Y(n23977) );
  MXI2XL U18654 ( .A(Q1[15]), .B(n23921), .S0(n23239), .Y(n3476) );
  XOR2XL U18655 ( .A(n23920), .B(n23919), .Y(n23921) );
  NAND2XL U18656 ( .A(n23918), .B(n23970), .Y(n23919) );
  AOI21XL U18657 ( .A0(n24084), .A1(n23915), .B0(n23914), .Y(n23920) );
  MXI2XL U18658 ( .A(Q1[14]), .B(n23828), .S0(n23239), .Y(n3477) );
  XNOR2XL U18659 ( .A(n24084), .B(n23827), .Y(n23828) );
  NAND2XL U18660 ( .A(n23915), .B(n23971), .Y(n23827) );
  MXI2XL U18661 ( .A(Q1[13]), .B(n23769), .S0(n23239), .Y(n3478) );
  XOR2XL U18662 ( .A(n23768), .B(n23767), .Y(n23769) );
  NAND2XL U18663 ( .A(n23766), .B(n23813), .Y(n23767) );
  AOI21XL U18664 ( .A0(n23763), .A1(n23762), .B0(n23761), .Y(n23768) );
  MXI2XL U18665 ( .A(Q1[12]), .B(n23738), .S0(n23239), .Y(n3479) );
  XNOR2XL U18666 ( .A(n23763), .B(n23737), .Y(n23738) );
  NAND2XL U18667 ( .A(n23762), .B(n23814), .Y(n23737) );
  MXI2XL U18668 ( .A(Q1[11]), .B(n23662), .S0(n23239), .Y(n3480) );
  AOI21XL U18669 ( .A0(n23656), .A1(n23655), .B0(n23654), .Y(n23661) );
  MXI2XL U18670 ( .A(Q1[10]), .B(n23594), .S0(n24128), .Y(n3481) );
  XOR2XL U18671 ( .A(n23734), .B(n23593), .Y(n23594) );
  NAND2XL U18672 ( .A(n23655), .B(n23730), .Y(n23593) );
  MXI2XL U18673 ( .A(Q1[9]), .B(n23569), .S0(n24128), .Y(n3482) );
  XOR2XL U18674 ( .A(n23568), .B(n23567), .Y(n23569) );
  NAND2XL U18675 ( .A(n23566), .B(n23584), .Y(n23567) );
  AOI21XL U18676 ( .A0(n23563), .A1(n23562), .B0(n23561), .Y(n23568) );
  MXI2XL U18677 ( .A(Q1[8]), .B(n23523), .S0(n23559), .Y(n3483) );
  XNOR2XL U18678 ( .A(n23563), .B(n23522), .Y(n23523) );
  NAND2XL U18679 ( .A(n23562), .B(n23585), .Y(n23522) );
  MXI2XL U18680 ( .A(Q1[7]), .B(n23441), .S0(n23559), .Y(n3484) );
  XNOR2XL U18681 ( .A(n23440), .B(n23439), .Y(n23441) );
  NAND2XL U18682 ( .A(n23438), .B(n23515), .Y(n23439) );
  MXI2XL U18683 ( .A(Q1[6]), .B(n23426), .S0(n23559), .Y(n3485) );
  XOR2XL U18684 ( .A(n23590), .B(n23425), .Y(n23426) );
  NAND2XL U18685 ( .A(n23424), .B(n23516), .Y(n23425) );
  INVXL U18686 ( .A(n23514), .Y(n23424) );
  MXI2XL U18687 ( .A(Q1[5]), .B(n23359), .S0(n23239), .Y(n3486) );
  XNOR2XL U18688 ( .A(n23358), .B(n23357), .Y(n23359) );
  NAND2XL U18689 ( .A(n23356), .B(n23413), .Y(n23357) );
  MXI2XL U18690 ( .A(Q1[4]), .B(n23318), .S0(n23239), .Y(n3487) );
  XOR2XL U18691 ( .A(n23353), .B(n23317), .Y(n23318) );
  NAND2XL U18692 ( .A(n23316), .B(n23414), .Y(n23317) );
  INVXL U18693 ( .A(n23411), .Y(n23316) );
  MXI2XL U18694 ( .A(Q1[3]), .B(n23240), .S0(n23239), .Y(n3488) );
  XOR2XL U18695 ( .A(n23238), .B(n23237), .Y(n23240) );
  NAND2XL U18696 ( .A(n23236), .B(n23310), .Y(n23237) );
  MXI2XL U18697 ( .A(Q1[2]), .B(n23193), .S0(n23239), .Y(n3489) );
  XNOR2XL U18698 ( .A(n23313), .B(n23192), .Y(n23193) );
  NAND2XL U18699 ( .A(n23233), .B(n23311), .Y(n23192) );
  MXI2XL U18700 ( .A(Q1[1]), .B(n23143), .S0(n23239), .Y(n3490) );
  XNOR2XL U18701 ( .A(n23142), .B(n23141), .Y(n23143) );
  NAND2XL U18702 ( .A(n23140), .B(n23184), .Y(n23141) );
  MXI2XL U18703 ( .A(Q1[0]), .B(n23130), .S0(n23239), .Y(n3491) );
  XOR2XL U18704 ( .A(n23137), .B(n23129), .Y(n23130) );
  NAND2XL U18705 ( .A(n23128), .B(n23185), .Y(n23129) );
  INVXL U18706 ( .A(n23183), .Y(n23128) );
  XOR2XL U18707 ( .A(n28914), .B(U0_pipe9[27]), .Y(n27069) );
  XOR2XL U18708 ( .A(n27066), .B(n27027), .Y(n27028) );
  NAND2XL U18709 ( .A(n27026), .B(n27064), .Y(n27027) );
  INVXL U18710 ( .A(n27065), .Y(n27026) );
  MXI2XL U18711 ( .A(Q1[51]), .B(n26985), .S0(n23239), .Y(n3494) );
  XNOR2XL U18712 ( .A(n27023), .B(n26984), .Y(n26985) );
  NAND2XL U18713 ( .A(n26981), .B(n27021), .Y(n26984) );
  MXI2XL U18714 ( .A(Q1[50]), .B(n26929), .S0(n23239), .Y(n3495) );
  NAND2XL U18715 ( .A(n26927), .B(n26978), .Y(n26928) );
  INVXL U18716 ( .A(n26979), .Y(n26927) );
  MXI2XL U18717 ( .A(Q1[49]), .B(n26887), .S0(n24128), .Y(n3496) );
  XNOR2XL U18718 ( .A(n26924), .B(n26886), .Y(n26887) );
  NAND2XL U18719 ( .A(n26883), .B(n26922), .Y(n26886) );
  MXI2XL U18720 ( .A(Q1[48]), .B(n26842), .S0(n23239), .Y(n3497) );
  XOR2XL U18721 ( .A(n26882), .B(n26841), .Y(n26842) );
  NAND2XL U18722 ( .A(n26840), .B(n26880), .Y(n26841) );
  INVXL U18723 ( .A(n26881), .Y(n26840) );
  MXI2XL U18724 ( .A(Q1[47]), .B(n26790), .S0(n24128), .Y(n3498) );
  XNOR2XL U18725 ( .A(n26837), .B(n26789), .Y(n26790) );
  NAND2XL U18726 ( .A(n26786), .B(n26835), .Y(n26789) );
  MXI2XL U18727 ( .A(Q1[46]), .B(n26752), .S0(n24128), .Y(n3499) );
  XOR2XL U18728 ( .A(n26751), .B(n26750), .Y(n26752) );
  NAND2XL U18729 ( .A(n26747), .B(n26780), .Y(n26750) );
  AOI21XL U18730 ( .A0(n26746), .A1(n26779), .B0(n26782), .Y(n26751) );
  MXI2XL U18731 ( .A(Q1[45]), .B(n26674), .S0(n23239), .Y(n3500) );
  XOR2XL U18732 ( .A(n26673), .B(n26672), .Y(n26674) );
  NAND2XL U18733 ( .A(n26671), .B(n26743), .Y(n26672) );
  AOI21XL U18734 ( .A0(n26746), .A1(n26668), .B0(n26667), .Y(n26673) );
  MXI2XL U18735 ( .A(Q1[44]), .B(n26625), .S0(n23239), .Y(n3501) );
  XOR2XL U18736 ( .A(n26624), .B(n26623), .Y(n26625) );
  NAND2XL U18737 ( .A(n26620), .B(n26664), .Y(n26623) );
  AOI21XL U18738 ( .A0(n26746), .A1(n26586), .B0(n26666), .Y(n26624) );
  MXI2XL U18739 ( .A(Q1[43]), .B(n26590), .S0(n24128), .Y(n3502) );
  XNOR2XL U18740 ( .A(n26746), .B(n26589), .Y(n26590) );
  NAND2XL U18741 ( .A(n26586), .B(n26619), .Y(n26589) );
  MXI2XL U18742 ( .A(Q1[42]), .B(n26511), .S0(n24128), .Y(n3503) );
  XOR2XL U18743 ( .A(n26510), .B(n26509), .Y(n26511) );
  NAND2XL U18744 ( .A(n26508), .B(n26574), .Y(n26509) );
  AOI21XL U18745 ( .A0(n26505), .A1(n26504), .B0(n26503), .Y(n26510) );
  MXI2XL U18746 ( .A(Q1[41]), .B(n26432), .S0(n23239), .Y(n3504) );
  XNOR2XL U18747 ( .A(n26505), .B(n26431), .Y(n26432) );
  NAND2XL U18748 ( .A(n26504), .B(n26575), .Y(n26431) );
  MXI2XL U18749 ( .A(Q1[40]), .B(n26379), .S0(n24128), .Y(n3505) );
  XOR2XL U18750 ( .A(n26378), .B(n26377), .Y(n26379) );
  NAND2XL U18751 ( .A(n26376), .B(n26423), .Y(n26377) );
  AOI21XL U18752 ( .A0(n26373), .A1(n26372), .B0(n26371), .Y(n26378) );
  MXI2XL U18753 ( .A(Q1[39]), .B(n26345), .S0(n24128), .Y(n3506) );
  XOR2XL U18754 ( .A(n26428), .B(n26344), .Y(n26345) );
  NAND2XL U18755 ( .A(n26372), .B(n26424), .Y(n26344) );
  MXI2XL U18756 ( .A(Q1[38]), .B(n26255), .S0(n23239), .Y(n3507) );
  XOR2XL U18757 ( .A(n26254), .B(n26253), .Y(n26255) );
  NAND2XL U18758 ( .A(n26252), .B(n26335), .Y(n26253) );
  AOI21XL U18759 ( .A0(n26249), .A1(n26248), .B0(n26247), .Y(n26254) );
  MXI2XL U18760 ( .A(Q1[37]), .B(n26205), .S0(n24128), .Y(n3508) );
  XNOR2XL U18761 ( .A(n26249), .B(n26204), .Y(n26205) );
  NAND2XL U18762 ( .A(n26248), .B(n26336), .Y(n26204) );
  MXI2XL U18763 ( .A(Q1[36]), .B(n26187), .S0(n24128), .Y(n3509) );
  XNOR2XL U18764 ( .A(n26186), .B(n26185), .Y(n26187) );
  NAND2XL U18765 ( .A(n26184), .B(n26197), .Y(n26185) );
  MXI2XL U18766 ( .A(Q1[35]), .B(n26103), .S0(n23239), .Y(n3510) );
  INVXL U18767 ( .A(n26196), .Y(n26101) );
  MXI2XL U18768 ( .A(Q1[34]), .B(n26078), .S0(n23239), .Y(n3511) );
  XNOR2XL U18769 ( .A(n26077), .B(n26076), .Y(n26078) );
  NAND2XL U18770 ( .A(n26075), .B(n26090), .Y(n26076) );
  MXI2XL U18771 ( .A(Q1[33]), .B(n26029), .S0(n23239), .Y(n3512) );
  XOR2XL U18772 ( .A(n26072), .B(n26028), .Y(n26029) );
  NAND2XL U18773 ( .A(n26027), .B(n26091), .Y(n26028) );
  INVXL U18774 ( .A(n26088), .Y(n26027) );
  MXI2XL U18775 ( .A(Q1[32]), .B(n25956), .S0(n24128), .Y(n3513) );
  XOR2XL U18776 ( .A(n25955), .B(n25954), .Y(n25956) );
  NAND2XL U18777 ( .A(n25953), .B(n26021), .Y(n25954) );
  AOI21XL U18778 ( .A0(n26024), .A1(n25950), .B0(n25949), .Y(n25955) );
  MXI2XL U18779 ( .A(Q1[31]), .B(n25905), .S0(n24128), .Y(n3514) );
  XNOR2XL U18780 ( .A(n26024), .B(n25904), .Y(n25905) );
  NAND2XL U18781 ( .A(n25950), .B(n26022), .Y(n25904) );
  MXI2XL U18782 ( .A(Q1[30]), .B(n25860), .S0(n23239), .Y(n3515) );
  XNOR2XL U18783 ( .A(n25859), .B(n25858), .Y(n25860) );
  NAND2XL U18784 ( .A(n25857), .B(n25896), .Y(n25858) );
  MXI2XL U18785 ( .A(Q1[29]), .B(n25836), .S0(n24128), .Y(n3516) );
  XOR2XL U18786 ( .A(n25854), .B(n25835), .Y(n25836) );
  NAND2XL U18787 ( .A(n25834), .B(n25897), .Y(n25835) );
  INVXL U18788 ( .A(n25895), .Y(n25834) );
  MXI2XL U18789 ( .A(Q1[28]), .B(n25798), .S0(n23239), .Y(n3517) );
  XOR2XL U18790 ( .A(n25797), .B(n25831), .Y(n25798) );
  NAND2XL U18791 ( .A(n25793), .B(n25829), .Y(n25797) );
  INVXL U18792 ( .A(n25830), .Y(n25793) );
  XOR2XL U18793 ( .A(n28690), .B(n28994), .Y(n24400) );
  XOR2XL U18794 ( .A(n24397), .B(n24360), .Y(n24361) );
  NAND2XL U18795 ( .A(n24359), .B(n24395), .Y(n24360) );
  INVXL U18796 ( .A(n24396), .Y(n24359) );
  MXI2XL U18797 ( .A(Q0[23]), .B(n24318), .S0(n24128), .Y(n3520) );
  XNOR2XL U18798 ( .A(n24356), .B(n24317), .Y(n24318) );
  NAND2XL U18799 ( .A(n24314), .B(n24354), .Y(n24317) );
  MXI2XL U18800 ( .A(Q0[22]), .B(n24277), .S0(n24128), .Y(n3521) );
  XOR2XL U18801 ( .A(n24313), .B(n24276), .Y(n24277) );
  NAND2XL U18802 ( .A(n24275), .B(n24311), .Y(n24276) );
  INVXL U18803 ( .A(n24312), .Y(n24275) );
  MXI2XL U18804 ( .A(Q0[21]), .B(n24235), .S0(n24128), .Y(n3522) );
  XNOR2XL U18805 ( .A(n24272), .B(n24234), .Y(n24235) );
  NAND2XL U18806 ( .A(n24231), .B(n24270), .Y(n24234) );
  MXI2XL U18807 ( .A(Q0[20]), .B(n24190), .S0(n24128), .Y(n3523) );
  XOR2XL U18808 ( .A(n24230), .B(n24189), .Y(n24190) );
  NAND2XL U18809 ( .A(n24188), .B(n24228), .Y(n24189) );
  INVXL U18810 ( .A(n24229), .Y(n24188) );
  MXI2XL U18811 ( .A(Q0[19]), .B(n24141), .S0(n24128), .Y(n3524) );
  XNOR2XL U18812 ( .A(n24185), .B(n24140), .Y(n24141) );
  NAND2XL U18813 ( .A(n24137), .B(n24183), .Y(n24140) );
  MXI2XL U18814 ( .A(Q0[18]), .B(n24079), .S0(n24128), .Y(n3525) );
  AOI21XL U18815 ( .A0(n24073), .A1(n24130), .B0(n24133), .Y(n24078) );
  MXI2XL U18816 ( .A(Q0[17]), .B(n24023), .S0(n24128), .Y(n3526) );
  XOR2XL U18817 ( .A(n24022), .B(n24021), .Y(n24023) );
  NAND2XL U18818 ( .A(n24020), .B(n24070), .Y(n24021) );
  AOI21XL U18819 ( .A0(n24073), .A1(n24017), .B0(n24016), .Y(n24022) );
  MXI2XL U18820 ( .A(Q0[16]), .B(n23968), .S0(n24128), .Y(n3527) );
  XOR2XL U18821 ( .A(n23967), .B(n23966), .Y(n23968) );
  NAND2XL U18822 ( .A(n23963), .B(n24013), .Y(n23966) );
  AOI21XL U18823 ( .A0(n24073), .A1(n24012), .B0(n24015), .Y(n23967) );
  MXI2XL U18824 ( .A(Q0[15]), .B(n23913), .S0(n24128), .Y(n3528) );
  XOR2XL U18825 ( .A(n23912), .B(n23911), .Y(n23913) );
  NAND2XL U18826 ( .A(n23910), .B(n23960), .Y(n23911) );
  AOI21XL U18827 ( .A0(n24073), .A1(n23907), .B0(n23906), .Y(n23912) );
  MXI2XL U18828 ( .A(Q0[14]), .B(n23847), .S0(n24128), .Y(n3529) );
  XNOR2XL U18829 ( .A(n24073), .B(n23846), .Y(n23847) );
  NAND2XL U18830 ( .A(n23907), .B(n23961), .Y(n23846) );
  MXI2XL U18831 ( .A(Q0[13]), .B(n23778), .S0(n24128), .Y(n3530) );
  XOR2XL U18832 ( .A(n23777), .B(n23776), .Y(n23778) );
  NAND2XL U18833 ( .A(n23775), .B(n23832), .Y(n23776) );
  AOI21XL U18834 ( .A0(n23772), .A1(n23771), .B0(n23770), .Y(n23777) );
  MXI2XL U18835 ( .A(Q0[12]), .B(n23727), .S0(n24128), .Y(n3531) );
  XNOR2XL U18836 ( .A(n23772), .B(n23726), .Y(n23727) );
  NAND2XL U18837 ( .A(n23771), .B(n23833), .Y(n23726) );
  MXI2XL U18838 ( .A(Q0[11]), .B(n23671), .S0(n24128), .Y(n3532) );
  XOR2XL U18839 ( .A(n23670), .B(n23669), .Y(n23671) );
  NAND2XL U18840 ( .A(n23668), .B(n23718), .Y(n23669) );
  MXI2XL U18841 ( .A(Q0[10]), .B(n23607), .S0(n23239), .Y(n3533) );
  XOR2XL U18842 ( .A(n23723), .B(n23606), .Y(n23607) );
  NAND2XL U18843 ( .A(n23664), .B(n23719), .Y(n23606) );
  MXI2XL U18844 ( .A(Q0[9]), .B(n23549), .S0(n23559), .Y(n3534) );
  XOR2XL U18845 ( .A(n23548), .B(n23547), .Y(n23549) );
  NAND2XL U18846 ( .A(n23546), .B(n23597), .Y(n23547) );
  AOI21XL U18847 ( .A0(n23543), .A1(n23542), .B0(n23541), .Y(n23548) );
  MXI2XL U18848 ( .A(Q0[8]), .B(n23507), .S0(n23559), .Y(n3535) );
  XNOR2XL U18849 ( .A(n23543), .B(n23506), .Y(n23507) );
  NAND2XL U18850 ( .A(n23542), .B(n23598), .Y(n23506) );
  MXI2XL U18851 ( .A(Q0[7]), .B(n23447), .S0(n23559), .Y(n3536) );
  XNOR2XL U18852 ( .A(n23446), .B(n23445), .Y(n23447) );
  NAND2XL U18853 ( .A(n23444), .B(n23499), .Y(n23445) );
  MXI2XL U18854 ( .A(Q0[6]), .B(n23403), .S0(n23239), .Y(n3537) );
  XOR2XL U18855 ( .A(n23603), .B(n23402), .Y(n23403) );
  NAND2XL U18856 ( .A(n23401), .B(n23500), .Y(n23402) );
  INVXL U18857 ( .A(n23498), .Y(n23401) );
  MXI2XL U18858 ( .A(Q0[5]), .B(n23342), .S0(n23239), .Y(n3538) );
  XNOR2XL U18859 ( .A(n23341), .B(n23340), .Y(n23342) );
  NAND2XL U18860 ( .A(n23339), .B(n23390), .Y(n23340) );
  MXI2XL U18861 ( .A(Q0[4]), .B(n23300), .S0(n23239), .Y(n3539) );
  XOR2XL U18862 ( .A(n23336), .B(n23299), .Y(n23300) );
  NAND2XL U18863 ( .A(n23298), .B(n23391), .Y(n23299) );
  INVXL U18864 ( .A(n23388), .Y(n23298) );
  MXI2XL U18865 ( .A(Q0[3]), .B(n23248), .S0(n23239), .Y(n3540) );
  AOI21XL U18866 ( .A0(n23295), .A1(n23242), .B0(n23241), .Y(n23247) );
  MXI2XL U18867 ( .A(Q0[2]), .B(n23204), .S0(n23239), .Y(n3541) );
  XNOR2XL U18868 ( .A(n23295), .B(n23203), .Y(n23204) );
  NAND2XL U18869 ( .A(n23242), .B(n23293), .Y(n23203) );
  MXI2XL U18870 ( .A(Q0[1]), .B(n23150), .S0(n23239), .Y(n3542) );
  XNOR2XL U18871 ( .A(n23149), .B(n23148), .Y(n23150) );
  NAND2XL U18872 ( .A(n23147), .B(n23195), .Y(n23148) );
  MXI2XL U18873 ( .A(Q0[0]), .B(n22431), .S0(n23239), .Y(n3543) );
  XOR2XL U18874 ( .A(n23144), .B(n22430), .Y(n22431) );
  NAND2XL U18875 ( .A(n22429), .B(n23196), .Y(n22430) );
  INVXL U18876 ( .A(n23194), .Y(n22429) );
  MXI2XL U18877 ( .A(Q0[28]), .B(n25121), .S0(n24128), .Y(n3544) );
  XOR2XL U18878 ( .A(n25814), .B(n25120), .Y(n25121) );
  NAND2XL U18879 ( .A(n25119), .B(n25863), .Y(n25120) );
  INVXL U18880 ( .A(n25861), .Y(n25119) );
  XOR2XL U18881 ( .A(n28917), .B(U0_pipe15[27]), .Y(n24386) );
  XOR2XL U18882 ( .A(n24383), .B(n24344), .Y(n24345) );
  NAND2XL U18883 ( .A(n24343), .B(n24381), .Y(n24344) );
  INVXL U18884 ( .A(n24382), .Y(n24343) );
  MXI2XL U18885 ( .A(Q3[23]), .B(n24302), .S0(n24128), .Y(n3547) );
  XNOR2XL U18886 ( .A(n24340), .B(n24301), .Y(n24302) );
  NAND2XL U18887 ( .A(n24298), .B(n24338), .Y(n24301) );
  MXI2XL U18888 ( .A(Q3[22]), .B(n24261), .S0(n24128), .Y(n3548) );
  XOR2XL U18889 ( .A(n24297), .B(n24260), .Y(n24261) );
  NAND2XL U18890 ( .A(n24259), .B(n24295), .Y(n24260) );
  INVXL U18891 ( .A(n24296), .Y(n24259) );
  MXI2XL U18892 ( .A(Q3[21]), .B(n24219), .S0(n24128), .Y(n3549) );
  XNOR2XL U18893 ( .A(n24256), .B(n24218), .Y(n24219) );
  NAND2XL U18894 ( .A(n24215), .B(n24254), .Y(n24218) );
  MXI2XL U18895 ( .A(Q3[20]), .B(n24174), .S0(n24128), .Y(n3550) );
  XOR2XL U18896 ( .A(n24214), .B(n24173), .Y(n24174) );
  NAND2XL U18897 ( .A(n24172), .B(n24212), .Y(n24173) );
  INVXL U18898 ( .A(n24213), .Y(n24172) );
  MXI2XL U18899 ( .A(Q3[19]), .B(n24116), .S0(n24128), .Y(n3551) );
  XNOR2XL U18900 ( .A(n24169), .B(n24115), .Y(n24116) );
  NAND2XL U18901 ( .A(n24112), .B(n24167), .Y(n24115) );
  MXI2XL U18902 ( .A(Q3[18]), .B(n24057), .S0(n24128), .Y(n3552) );
  XOR2XL U18903 ( .A(n24056), .B(n24055), .Y(n24057) );
  NAND2XL U18904 ( .A(n24052), .B(n24106), .Y(n24055) );
  AOI21XL U18905 ( .A0(n24051), .A1(n24105), .B0(n24108), .Y(n24056) );
  MXI2XL U18906 ( .A(Q3[17]), .B(n23999), .S0(n24128), .Y(n3553) );
  XOR2XL U18907 ( .A(n23998), .B(n23997), .Y(n23999) );
  NAND2XL U18908 ( .A(n23996), .B(n24048), .Y(n23997) );
  AOI21XL U18909 ( .A0(n24051), .A1(n23993), .B0(n23992), .Y(n23998) );
  MXI2XL U18910 ( .A(Q3[16]), .B(n23948), .S0(n24128), .Y(n3554) );
  XOR2XL U18911 ( .A(n23947), .B(n23946), .Y(n23948) );
  NAND2XL U18912 ( .A(n23943), .B(n23989), .Y(n23946) );
  MXI2XL U18913 ( .A(Q3[15]), .B(n23897), .S0(n24128), .Y(n3555) );
  MXI2XL U18914 ( .A(Q3[14]), .B(n23809), .S0(n24128), .Y(n3556) );
  XOR2XL U18915 ( .A(n23808), .B(n23807), .Y(n23809) );
  NAND2XL U18916 ( .A(n23806), .B(n23881), .Y(n23807) );
  AOI21XL U18917 ( .A0(n23803), .A1(n23802), .B0(n23801), .Y(n23808) );
  MXI2XL U18918 ( .A(Q3[13]), .B(n23760), .S0(n24128), .Y(n3557) );
  XNOR2XL U18919 ( .A(n23803), .B(n23759), .Y(n23760) );
  NAND2XL U18920 ( .A(n23802), .B(n23882), .Y(n23759) );
  MXI2XL U18921 ( .A(Q3[12]), .B(n23705), .S0(n24128), .Y(n3558) );
  XOR2XL U18922 ( .A(n23704), .B(n23703), .Y(n23705) );
  NAND2XL U18923 ( .A(n23702), .B(n23751), .Y(n23703) );
  AOI21XL U18924 ( .A0(n23699), .A1(n23698), .B0(n23697), .Y(n23704) );
  MXI2XL U18925 ( .A(Q3[11]), .B(n23653), .S0(n24128), .Y(n3559) );
  XOR2XL U18926 ( .A(n23756), .B(n23652), .Y(n23653) );
  NAND2XL U18927 ( .A(n23698), .B(n23752), .Y(n23652) );
  MXI2XL U18928 ( .A(Q3[10]), .B(n23616), .S0(n24128), .Y(n3560) );
  XOR2XL U18929 ( .A(n23615), .B(n23614), .Y(n23616) );
  NAND2XL U18930 ( .A(n23613), .B(n23643), .Y(n23614) );
  AOI21XL U18931 ( .A0(n23610), .A1(n23609), .B0(n23608), .Y(n23615) );
  MXI2XL U18932 ( .A(Q3[9]), .B(n23560), .S0(n23559), .Y(n3561) );
  XNOR2XL U18933 ( .A(n23610), .B(n23558), .Y(n23560) );
  NAND2XL U18934 ( .A(n23609), .B(n23644), .Y(n23558) );
  MXI2XL U18935 ( .A(Q3[8]), .B(n23513), .S0(n23559), .Y(n3562) );
  XNOR2XL U18936 ( .A(n23512), .B(n23511), .Y(n23513) );
  NAND2XL U18937 ( .A(n23510), .B(n23551), .Y(n23511) );
  MXI2XL U18938 ( .A(Q3[7]), .B(n23463), .S0(n23559), .Y(n3563) );
  XOR2XL U18939 ( .A(n23649), .B(n23462), .Y(n23463) );
  NAND2XL U18940 ( .A(n23461), .B(n23552), .Y(n23462) );
  INVXL U18941 ( .A(n23550), .Y(n23461) );
  MXI2XL U18942 ( .A(Q3[6]), .B(n23410), .S0(n23559), .Y(n3564) );
  XNOR2XL U18943 ( .A(n23409), .B(n23408), .Y(n23410) );
  NAND2XL U18944 ( .A(n23407), .B(n23450), .Y(n23408) );
  MXI2XL U18945 ( .A(Q3[5]), .B(n23352), .S0(n24128), .Y(n3565) );
  XOR2XL U18946 ( .A(n23404), .B(n23351), .Y(n23352) );
  NAND2XL U18947 ( .A(n23350), .B(n23451), .Y(n23351) );
  INVXL U18948 ( .A(n23448), .Y(n23350) );
  MXI2XL U18949 ( .A(Q3[4]), .B(n23308), .S0(n24128), .Y(n3566) );
  XOR2XL U18950 ( .A(n23307), .B(n23306), .Y(n23308) );
  NAND2XL U18951 ( .A(n23305), .B(n23344), .Y(n23306) );
  AOI21XL U18952 ( .A0(n23347), .A1(n23302), .B0(n23301), .Y(n23307) );
  MXI2XL U18953 ( .A(Q3[3]), .B(n23259), .S0(n24128), .Y(n3567) );
  XNOR2XL U18954 ( .A(n23347), .B(n23258), .Y(n23259) );
  NAND2XL U18955 ( .A(n23302), .B(n23345), .Y(n23258) );
  MXI2XL U18956 ( .A(Q3[2]), .B(n23211), .S0(n23239), .Y(n3568) );
  XNOR2XL U18957 ( .A(n23210), .B(n23209), .Y(n23211) );
  NAND2XL U18958 ( .A(n23208), .B(n23250), .Y(n23209) );
  MXI2XL U18959 ( .A(Q3[1]), .B(n23158), .S0(n23239), .Y(n3569) );
  XOR2XL U18960 ( .A(n23205), .B(n23157), .Y(n23158) );
  NAND2XL U18961 ( .A(n23156), .B(n23251), .Y(n23157) );
  INVXL U18962 ( .A(n23249), .Y(n23156) );
  MXI2XL U18963 ( .A(Q3[0]), .B(n22734), .S0(n23239), .Y(n3570) );
  NAND2XL U18964 ( .A(n22729), .B(n23151), .Y(n22733) );
  INVXL U18965 ( .A(n23152), .Y(n22729) );
  XOR2XL U18966 ( .A(n28916), .B(U0_pipe13[27]), .Y(n27048) );
  XOR2XL U18967 ( .A(n27045), .B(n27003), .Y(n27004) );
  NAND2XL U18968 ( .A(n27002), .B(n27043), .Y(n27003) );
  INVXL U18969 ( .A(n27044), .Y(n27002) );
  MXI2XL U18970 ( .A(Q3[51]), .B(n26961), .S0(n24128), .Y(n3573) );
  XNOR2XL U18971 ( .A(n26999), .B(n26960), .Y(n26961) );
  NAND2XL U18972 ( .A(n26957), .B(n26997), .Y(n26960) );
  MXI2XL U18973 ( .A(Q3[50]), .B(n26921), .S0(n24128), .Y(n3574) );
  XOR2XL U18974 ( .A(n26956), .B(n26920), .Y(n26921) );
  NAND2XL U18975 ( .A(n26919), .B(n26954), .Y(n26920) );
  INVXL U18976 ( .A(n26955), .Y(n26919) );
  MXI2XL U18977 ( .A(Q3[49]), .B(n26879), .S0(n23239), .Y(n3575) );
  XNOR2XL U18978 ( .A(n26916), .B(n26878), .Y(n26879) );
  NAND2XL U18979 ( .A(n26875), .B(n26914), .Y(n26878) );
  MXI2XL U18980 ( .A(Q3[48]), .B(n26834), .S0(n23239), .Y(n3576) );
  XOR2XL U18981 ( .A(n26874), .B(n26833), .Y(n26834) );
  NAND2XL U18982 ( .A(n26832), .B(n26872), .Y(n26833) );
  INVXL U18983 ( .A(n26873), .Y(n26832) );
  MXI2XL U18984 ( .A(Q3[47]), .B(n26778), .S0(n23239), .Y(n3577) );
  XNOR2XL U18985 ( .A(n26829), .B(n26777), .Y(n26778) );
  NAND2XL U18986 ( .A(n26774), .B(n26827), .Y(n26777) );
  MXI2XL U18987 ( .A(Q3[46]), .B(n26719), .S0(n23239), .Y(n3578) );
  XOR2XL U18988 ( .A(n26718), .B(n26717), .Y(n26719) );
  NAND2XL U18989 ( .A(n26714), .B(n26768), .Y(n26717) );
  AOI21XL U18990 ( .A0(n26713), .A1(n26767), .B0(n26770), .Y(n26718) );
  MXI2XL U18991 ( .A(Q3[45]), .B(n26663), .S0(n24128), .Y(n3579) );
  XOR2XL U18992 ( .A(n26662), .B(n26661), .Y(n26663) );
  NAND2XL U18993 ( .A(n26660), .B(n26710), .Y(n26661) );
  AOI21XL U18994 ( .A0(n26713), .A1(n26657), .B0(n26656), .Y(n26662) );
  MXI2XL U18995 ( .A(Q3[44]), .B(n26618), .S0(n23239), .Y(n3580) );
  XOR2XL U18996 ( .A(n26617), .B(n26616), .Y(n26618) );
  NAND2XL U18997 ( .A(n26613), .B(n26653), .Y(n26616) );
  AOI21XL U18998 ( .A0(n26713), .A1(n26538), .B0(n26655), .Y(n26617) );
  MXI2XL U18999 ( .A(Q3[43]), .B(n26542), .S0(n23239), .Y(n3581) );
  XNOR2XL U19000 ( .A(n26713), .B(n26541), .Y(n26542) );
  NAND2XL U19001 ( .A(n26538), .B(n26612), .Y(n26541) );
  MXI2XL U19002 ( .A(Q3[42]), .B(n26474), .S0(n23239), .Y(n3582) );
  XOR2XL U19003 ( .A(n26473), .B(n26472), .Y(n26474) );
  NAND2XL U19004 ( .A(n26471), .B(n26526), .Y(n26472) );
  AOI21XL U19005 ( .A0(n26468), .A1(n26467), .B0(n26466), .Y(n26473) );
  MXI2XL U19006 ( .A(Q3[41]), .B(n26421), .S0(n24128), .Y(n3583) );
  XNOR2XL U19007 ( .A(n26468), .B(n26420), .Y(n26421) );
  NAND2XL U19008 ( .A(n26467), .B(n26527), .Y(n26420) );
  MXI2XL U19009 ( .A(Q3[40]), .B(n26370), .S0(n24128), .Y(n3584) );
  XOR2XL U19010 ( .A(n26369), .B(n26368), .Y(n26370) );
  NAND2XL U19011 ( .A(n26367), .B(n26412), .Y(n26368) );
  AOI21XL U19012 ( .A0(n26364), .A1(n26363), .B0(n26362), .Y(n26369) );
  MXI2XL U19013 ( .A(Q3[39]), .B(n26310), .S0(n23239), .Y(n3585) );
  NAND2XL U19014 ( .A(n26363), .B(n26413), .Y(n26309) );
  MXI2XL U19015 ( .A(Q3[38]), .B(n26277), .S0(n23239), .Y(n3586) );
  XOR2XL U19016 ( .A(n26276), .B(n26275), .Y(n26277) );
  NAND2XL U19017 ( .A(n26274), .B(n26300), .Y(n26275) );
  AOI21XL U19018 ( .A0(n26271), .A1(n26270), .B0(n26269), .Y(n26276) );
  MXI2XL U19019 ( .A(Q3[37]), .B(n26224), .S0(n24128), .Y(n3587) );
  XNOR2XL U19020 ( .A(n26271), .B(n26223), .Y(n26224) );
  NAND2XL U19021 ( .A(n26270), .B(n26301), .Y(n26223) );
  MXI2XL U19022 ( .A(Q3[36]), .B(n26181), .S0(n23239), .Y(n3588) );
  XNOR2XL U19023 ( .A(n26180), .B(n26179), .Y(n26181) );
  NAND2XL U19024 ( .A(n26178), .B(n26216), .Y(n26179) );
  MXI2XL U19025 ( .A(Q3[35]), .B(n26125), .S0(n24128), .Y(n3589) );
  XOR2XL U19026 ( .A(n26306), .B(n26124), .Y(n26125) );
  NAND2XL U19027 ( .A(n26123), .B(n26217), .Y(n26124) );
  INVXL U19028 ( .A(n26215), .Y(n26123) );
  MXI2XL U19029 ( .A(Q3[34]), .B(n26071), .S0(n24128), .Y(n3590) );
  XNOR2XL U19030 ( .A(n26070), .B(n26069), .Y(n26071) );
  NAND2XL U19031 ( .A(n26068), .B(n26112), .Y(n26069) );
  MXI2XL U19032 ( .A(Q3[33]), .B(n26019), .S0(n23239), .Y(n3591) );
  XOR2XL U19033 ( .A(n26065), .B(n26018), .Y(n26019) );
  NAND2XL U19034 ( .A(n26017), .B(n26113), .Y(n26018) );
  INVXL U19035 ( .A(n26110), .Y(n26017) );
  MXI2XL U19036 ( .A(Q3[32]), .B(n25974), .S0(n24128), .Y(n3592) );
  XOR2XL U19037 ( .A(n25973), .B(n25972), .Y(n25974) );
  NAND2XL U19038 ( .A(n25971), .B(n26011), .Y(n25972) );
  AOI21XL U19039 ( .A0(n26014), .A1(n25968), .B0(n25967), .Y(n25973) );
  MXI2XL U19040 ( .A(Q3[31]), .B(n25924), .S0(n23239), .Y(n3593) );
  XNOR2XL U19041 ( .A(n26014), .B(n25923), .Y(n25924) );
  NAND2XL U19042 ( .A(n25968), .B(n26012), .Y(n25923) );
  MXI2XL U19043 ( .A(Q3[30]), .B(n25878), .S0(n23239), .Y(n3594) );
  XNOR2XL U19044 ( .A(n25877), .B(n25876), .Y(n25878) );
  NAND2XL U19045 ( .A(n25875), .B(n25915), .Y(n25876) );
  MXI2XL U19046 ( .A(Q3[29]), .B(n25828), .S0(n24128), .Y(n3595) );
  XOR2XL U19047 ( .A(n25872), .B(n25827), .Y(n25828) );
  NAND2XL U19048 ( .A(n25826), .B(n25916), .Y(n25827) );
  INVXL U19049 ( .A(n25914), .Y(n25826) );
  MXI2XL U19050 ( .A(Q3[28]), .B(n25456), .S0(n23239), .Y(n3596) );
  NAND2XL U19051 ( .A(n25451), .B(n25821), .Y(n25455) );
  INVXL U19052 ( .A(n25822), .Y(n25451) );
  XOR2XL U19053 ( .A(n28692), .B(n28996), .Y(n24393) );
  XOR2XL U19054 ( .A(n24390), .B(n24368), .Y(n24369) );
  NAND2XL U19055 ( .A(n24367), .B(n24388), .Y(n24368) );
  INVXL U19056 ( .A(n24389), .Y(n24367) );
  MXI2XL U19057 ( .A(Q2[23]), .B(n24326), .S0(n23239), .Y(n3599) );
  XNOR2XL U19058 ( .A(n24364), .B(n24325), .Y(n24326) );
  NAND2XL U19059 ( .A(n24322), .B(n24362), .Y(n24325) );
  MXI2XL U19060 ( .A(Q2[22]), .B(n24269), .S0(n23239), .Y(n3600) );
  XOR2XL U19061 ( .A(n24321), .B(n24268), .Y(n24269) );
  NAND2XL U19062 ( .A(n24267), .B(n24319), .Y(n24268) );
  INVXL U19063 ( .A(n24320), .Y(n24267) );
  MXI2XL U19064 ( .A(Q2[21]), .B(n24227), .S0(n23239), .Y(n3601) );
  XNOR2XL U19065 ( .A(n24264), .B(n24226), .Y(n24227) );
  NAND2XL U19066 ( .A(n24223), .B(n24262), .Y(n24226) );
  MXI2XL U19067 ( .A(Q2[20]), .B(n24182), .S0(n23239), .Y(n3602) );
  XOR2XL U19068 ( .A(n24222), .B(n24181), .Y(n24182) );
  NAND2XL U19069 ( .A(n24180), .B(n24220), .Y(n24181) );
  INVXL U19070 ( .A(n24221), .Y(n24180) );
  MXI2XL U19071 ( .A(Q2[19]), .B(n24153), .S0(n23239), .Y(n3603) );
  XNOR2XL U19072 ( .A(n24177), .B(n24152), .Y(n24153) );
  NAND2XL U19073 ( .A(n24149), .B(n24175), .Y(n24152) );
  MXI2XL U19074 ( .A(Q2[18]), .B(n24068), .S0(n24128), .Y(n3604) );
  XOR2XL U19075 ( .A(n24067), .B(n24066), .Y(n24068) );
  NAND2XL U19076 ( .A(n24063), .B(n24143), .Y(n24066) );
  AOI21XL U19077 ( .A0(n24062), .A1(n24142), .B0(n24145), .Y(n24067) );
  MXI2XL U19078 ( .A(Q2[17]), .B(n24035), .S0(n24128), .Y(n3605) );
  XOR2XL U19079 ( .A(n24034), .B(n24033), .Y(n24035) );
  NAND2XL U19080 ( .A(n24032), .B(n24059), .Y(n24033) );
  AOI21XL U19081 ( .A0(n24062), .A1(n24029), .B0(n24028), .Y(n24034) );
  MXI2XL U19082 ( .A(Q2[16]), .B(n23958), .S0(n24128), .Y(n3606) );
  XOR2XL U19083 ( .A(n23957), .B(n23956), .Y(n23958) );
  NAND2XL U19084 ( .A(n23953), .B(n24025), .Y(n23956) );
  AOI21XL U19085 ( .A0(n24062), .A1(n24024), .B0(n24027), .Y(n23957) );
  MXI2XL U19086 ( .A(Q2[15]), .B(n23905), .S0(n23239), .Y(n3607) );
  XOR2XL U19087 ( .A(n23904), .B(n23903), .Y(n23905) );
  NAND2XL U19088 ( .A(n23902), .B(n23950), .Y(n23903) );
  AOI21XL U19089 ( .A0(n24062), .A1(n23899), .B0(n23898), .Y(n23904) );
  MXI2XL U19090 ( .A(Q2[14]), .B(n23866), .S0(n23239), .Y(n3608) );
  MXI2XL U19091 ( .A(Q2[13]), .B(n23787), .S0(n23239), .Y(n3609) );
  XOR2XL U19092 ( .A(n23786), .B(n23785), .Y(n23787) );
  NAND2XL U19093 ( .A(n23784), .B(n23851), .Y(n23785) );
  AOI21XL U19094 ( .A0(n23781), .A1(n23780), .B0(n23779), .Y(n23786) );
  MXI2XL U19095 ( .A(Q2[12]), .B(n23716), .S0(n23239), .Y(n3610) );
  XNOR2XL U19096 ( .A(n23781), .B(n23715), .Y(n23716) );
  NAND2XL U19097 ( .A(n23780), .B(n23852), .Y(n23715) );
  MXI2XL U19098 ( .A(Q2[11]), .B(n23680), .S0(n23239), .Y(n3611) );
  XOR2XL U19099 ( .A(n23679), .B(n23678), .Y(n23680) );
  NAND2XL U19100 ( .A(n23677), .B(n23707), .Y(n23678) );
  AOI21XL U19101 ( .A0(n23674), .A1(n23673), .B0(n23672), .Y(n23679) );
  MXI2XL U19102 ( .A(Q2[10]), .B(n23629), .S0(n23239), .Y(n3612) );
  XOR2XL U19103 ( .A(n23712), .B(n23628), .Y(n23629) );
  NAND2XL U19104 ( .A(n23673), .B(n23708), .Y(n23628) );
  MXI2XL U19105 ( .A(Q2[9]), .B(n23540), .S0(n23559), .Y(n3613) );
  XOR2XL U19106 ( .A(n23539), .B(n23538), .Y(n23540) );
  NAND2XL U19107 ( .A(n23537), .B(n23619), .Y(n23538) );
  MXI2XL U19108 ( .A(Q2[8]), .B(n23497), .S0(n23559), .Y(n3614) );
  XNOR2XL U19109 ( .A(n23534), .B(n23496), .Y(n23497) );
  NAND2XL U19110 ( .A(n23533), .B(n23620), .Y(n23496) );
  MXI2XL U19111 ( .A(Q2[7]), .B(n23469), .S0(n23559), .Y(n3615) );
  XNOR2XL U19112 ( .A(n23468), .B(n23467), .Y(n23469) );
  NAND2XL U19113 ( .A(n23466), .B(n23489), .Y(n23467) );
  MXI2XL U19114 ( .A(Q2[6]), .B(n23387), .S0(n24128), .Y(n3616) );
  XOR2XL U19115 ( .A(n23625), .B(n23386), .Y(n23387) );
  NAND2XL U19116 ( .A(n23385), .B(n23490), .Y(n23386) );
  INVXL U19117 ( .A(n23488), .Y(n23385) );
  MXI2XL U19118 ( .A(Q2[5]), .B(n23335), .S0(n24128), .Y(n3617) );
  XNOR2XL U19119 ( .A(n23334), .B(n23333), .Y(n23335) );
  NAND2XL U19120 ( .A(n23332), .B(n23374), .Y(n23333) );
  MXI2XL U19121 ( .A(Q2[4]), .B(n23290), .S0(n24128), .Y(n3618) );
  XOR2XL U19122 ( .A(n23329), .B(n23289), .Y(n23290) );
  NAND2XL U19123 ( .A(n23288), .B(n23375), .Y(n23289) );
  INVXL U19124 ( .A(n23372), .Y(n23288) );
  MXI2XL U19125 ( .A(Q2[3]), .B(n23267), .S0(n23239), .Y(n3619) );
  AOI21XL U19126 ( .A0(n23285), .A1(n23261), .B0(n23260), .Y(n23266) );
  MXI2XL U19127 ( .A(Q2[2]), .B(n23222), .S0(n23239), .Y(n3620) );
  XNOR2XL U19128 ( .A(n23285), .B(n23221), .Y(n23222) );
  NAND2XL U19129 ( .A(n23261), .B(n23283), .Y(n23221) );
  MXI2XL U19130 ( .A(Q2[1]), .B(n23165), .S0(n23239), .Y(n3621) );
  XNOR2XL U19131 ( .A(n23164), .B(n23163), .Y(n23165) );
  NAND2XL U19132 ( .A(n23162), .B(n23213), .Y(n23163) );
  MXI2XL U19133 ( .A(Q2[0]), .B(n22107), .S0(n23239), .Y(n3622) );
  XOR2XL U19134 ( .A(n23159), .B(n22106), .Y(n22107) );
  NAND2XL U19135 ( .A(n22105), .B(n23214), .Y(n22106) );
  INVXL U19136 ( .A(n23212), .Y(n22105) );
  XOR2XL U19137 ( .A(n28915), .B(U0_pipe3[27]), .Y(n27055) );
  XOR2XL U19138 ( .A(n27052), .B(n27011), .Y(n27012) );
  NAND2XL U19139 ( .A(n27010), .B(n27050), .Y(n27011) );
  INVXL U19140 ( .A(n27051), .Y(n27010) );
  MXI2XL U19141 ( .A(Q2[51]), .B(n26969), .S0(n23239), .Y(n3625) );
  XNOR2XL U19142 ( .A(n27007), .B(n26968), .Y(n26969) );
  NAND2XL U19143 ( .A(n26965), .B(n27005), .Y(n26968) );
  MXI2XL U19144 ( .A(Q2[50]), .B(n26945), .S0(n24128), .Y(n3626) );
  XOR2XL U19145 ( .A(n26964), .B(n26944), .Y(n26945) );
  NAND2XL U19146 ( .A(n26943), .B(n26962), .Y(n26944) );
  INVXL U19147 ( .A(n26963), .Y(n26943) );
  MXI2XL U19148 ( .A(Q2[49]), .B(n26903), .S0(n24128), .Y(n3627) );
  XNOR2XL U19149 ( .A(n26940), .B(n26902), .Y(n26903) );
  NAND2XL U19150 ( .A(n26899), .B(n26938), .Y(n26902) );
  MXI2XL U19151 ( .A(Q2[48]), .B(n26858), .S0(n24128), .Y(n3628) );
  XOR2XL U19152 ( .A(n26898), .B(n26857), .Y(n26858) );
  NAND2XL U19153 ( .A(n26856), .B(n26896), .Y(n26857) );
  INVXL U19154 ( .A(n26897), .Y(n26856) );
  MXI2XL U19155 ( .A(Q2[47]), .B(n26814), .S0(n23239), .Y(n3629) );
  XNOR2XL U19156 ( .A(n26853), .B(n26813), .Y(n26814) );
  NAND2XL U19157 ( .A(n26810), .B(n26851), .Y(n26813) );
  MXI2XL U19158 ( .A(Q2[46]), .B(n26730), .S0(n24128), .Y(n3630) );
  XOR2XL U19159 ( .A(n26729), .B(n26728), .Y(n26730) );
  NAND2XL U19160 ( .A(n26725), .B(n26804), .Y(n26728) );
  AOI21XL U19161 ( .A0(n26724), .A1(n26803), .B0(n26806), .Y(n26729) );
  MXI2XL U19162 ( .A(Q2[45]), .B(n26697), .S0(n23239), .Y(n3631) );
  NAND2XL U19163 ( .A(n26694), .B(n26721), .Y(n26695) );
  AOI21XL U19164 ( .A0(n26724), .A1(n26691), .B0(n26690), .Y(n26696) );
  MXI2XL U19165 ( .A(Q2[44]), .B(n26642), .S0(n24128), .Y(n3632) );
  XOR2XL U19166 ( .A(n26641), .B(n26640), .Y(n26642) );
  NAND2XL U19167 ( .A(n26637), .B(n26687), .Y(n26640) );
  AOI21XL U19168 ( .A0(n26724), .A1(n26558), .B0(n26689), .Y(n26641) );
  MXI2XL U19169 ( .A(Q2[43]), .B(n26562), .S0(n23239), .Y(n3633) );
  XNOR2XL U19170 ( .A(n26724), .B(n26561), .Y(n26562) );
  NAND2XL U19171 ( .A(n26558), .B(n26636), .Y(n26561) );
  MXI2XL U19172 ( .A(Q2[42]), .B(n26483), .S0(n24128), .Y(n3634) );
  XOR2XL U19173 ( .A(n26482), .B(n26481), .Y(n26483) );
  NAND2XL U19174 ( .A(n26480), .B(n26546), .Y(n26481) );
  AOI21XL U19175 ( .A0(n26477), .A1(n26476), .B0(n26475), .Y(n26482) );
  MXI2XL U19176 ( .A(Q2[41]), .B(n26452), .S0(n24128), .Y(n3635) );
  XNOR2XL U19177 ( .A(n26477), .B(n26451), .Y(n26452) );
  NAND2XL U19178 ( .A(n26476), .B(n26547), .Y(n26451) );
  OAI211XL U19179 ( .A0(n5836), .A1(n15985), .B0(n15984), .C0(n15983), .Y(
        n15986) );
  AOI22XL U19180 ( .A0(B7_q[0]), .A1(n15982), .B0(B6_q[0]), .B1(n15958), .Y(
        n15984) );
  OAI211XL U19181 ( .A0(n15495), .A1(n15578), .B0(n15577), .C0(n15576), .Y(
        n15579) );
  AOI21XL U19182 ( .A0(B4_q[0]), .A1(n15557), .B0(n5924), .Y(n15576) );
  AOI22XL U19183 ( .A0(B5_q[0]), .A1(n16165), .B0(B7_q[0]), .B1(n16128), .Y(
        n15577) );
  NAND4XL U19184 ( .A(n15939), .B(n15938), .C(n5909), .D(n15937), .Y(n15940)
         );
  NAND2XL U19185 ( .A(B5_q[10]), .B(n15963), .Y(n15939) );
  NAND2XL U19186 ( .A(B4_q[10]), .B(n5925), .Y(n15938) );
  NAND4XL U19187 ( .A(n15733), .B(n15732), .C(n5800), .D(n15731), .Y(n15734)
         );
  NAND2XL U19188 ( .A(B4_q[10]), .B(n15687), .Y(n15733) );
  NAND2XL U19189 ( .A(B6_q[10]), .B(n16293), .Y(n15732) );
  NAND4XL U19190 ( .A(n15541), .B(n15540), .C(n5800), .D(n15539), .Y(n15542)
         );
  NAND2XL U19191 ( .A(B4_q[10]), .B(n15557), .Y(n15541) );
  NAND2XL U19192 ( .A(B6_q[10]), .B(n16161), .Y(n15540) );
  NAND4XL U19193 ( .A(n15339), .B(n15338), .C(n5800), .D(n15337), .Y(n15340)
         );
  NAND2XL U19194 ( .A(B7_q[10]), .B(n16569), .Y(n15339) );
  NAND2XL U19195 ( .A(B4_q[10]), .B(n7126), .Y(n15338) );
  NAND4XL U19196 ( .A(n15935), .B(n15934), .C(n5908), .D(n15933), .Y(n15936)
         );
  NAND2XL U19197 ( .A(B4_q[11]), .B(n5925), .Y(n15935) );
  NAND2XL U19198 ( .A(B5_q[11]), .B(n15963), .Y(n15934) );
  NAND4XL U19199 ( .A(n15729), .B(n15728), .C(R7_valid), .D(n15727), .Y(n15730) );
  NAND2XL U19200 ( .A(B4_q[11]), .B(n15687), .Y(n15729) );
  NAND2XL U19201 ( .A(B7_q[11]), .B(n16325), .Y(n15728) );
  NAND4XL U19202 ( .A(n15332), .B(n15331), .C(n5915), .D(n15330), .Y(n15333)
         );
  NAND2XL U19203 ( .A(B6_q[11]), .B(n16570), .Y(n15332) );
  NAND2XL U19204 ( .A(B5_q[11]), .B(n16375), .Y(n15331) );
  NAND4XL U19205 ( .A(n15931), .B(n15930), .C(n5800), .D(n15929), .Y(n15932)
         );
  NAND2XL U19206 ( .A(B4_q[12]), .B(n5925), .Y(n15931) );
  NAND2XL U19207 ( .A(B7_q[12]), .B(n5930), .Y(n15930) );
  NAND4XL U19208 ( .A(n15725), .B(n15724), .C(n5915), .D(n15723), .Y(n15726)
         );
  NAND2XL U19209 ( .A(B4_q[12]), .B(n15687), .Y(n15725) );
  NAND2XL U19210 ( .A(B7_q[12]), .B(n16325), .Y(n15724) );
  NAND4XL U19211 ( .A(n15533), .B(n15532), .C(n6880), .D(n15531), .Y(n15534)
         );
  NAND2XL U19212 ( .A(B6_q[12]), .B(n16161), .Y(n15533) );
  NAND2XL U19213 ( .A(B4_q[12]), .B(n15557), .Y(n15532) );
  NAND4XL U19214 ( .A(n15324), .B(n15323), .C(n5800), .D(n15322), .Y(n15325)
         );
  NAND2XL U19215 ( .A(B5_q[12]), .B(n16375), .Y(n15324) );
  NAND2XL U19216 ( .A(B4_q[12]), .B(n7126), .Y(n15323) );
  OAI211XL U19217 ( .A0(n15967), .A1(n15927), .B0(n15926), .C0(n15925), .Y(
        n15928) );
  AOI22XL U19218 ( .A0(B5_q[13]), .A1(n15963), .B0(B6_q[13]), .B1(n15958), .Y(
        n15926) );
  OAI211XL U19219 ( .A0(n5841), .A1(n15927), .B0(n15529), .C0(n15528), .Y(
        n15530) );
  AOI22XL U19220 ( .A0(B5_q[13]), .A1(n16165), .B0(B6_q[13]), .B1(n16143), .Y(
        n15529) );
  AOI21XL U19221 ( .A0(B4_q[13]), .A1(n5933), .B0(n28985), .Y(n15528) );
  OAI211XL U19222 ( .A0(n15316), .A1(n5914), .B0(n15315), .C0(n15314), .Y(
        n15317) );
  AOI21XL U19223 ( .A0(B7_q[13]), .A1(n7127), .B0(n5924), .Y(n15314) );
  AOI22XL U19224 ( .A0(B5_q[13]), .A1(n16559), .B0(B6_q[13]), .B1(n16570), .Y(
        n15315) );
  NAND4XL U19225 ( .A(n15923), .B(n15922), .C(n5912), .D(n15921), .Y(n15924)
         );
  NAND2XL U19226 ( .A(B4_q[14]), .B(n5925), .Y(n15923) );
  NAND2XL U19227 ( .A(B7_q[14]), .B(n15982), .Y(n15922) );
  NAND4XL U19228 ( .A(n15717), .B(n15716), .C(n5913), .D(n15715), .Y(n15718)
         );
  NAND2XL U19229 ( .A(B5_q[14]), .B(n15747), .Y(n15717) );
  NAND2XL U19230 ( .A(B4_q[14]), .B(n15687), .Y(n15716) );
  NAND4XL U19231 ( .A(n15526), .B(n15525), .C(n5800), .D(n15524), .Y(n15527)
         );
  NAND2XL U19232 ( .A(B4_q[14]), .B(n15557), .Y(n15526) );
  NAND2XL U19233 ( .A(B7_q[14]), .B(n16158), .Y(n15525) );
  NAND4XL U19234 ( .A(n15308), .B(n15307), .C(n5800), .D(n15306), .Y(n15309)
         );
  NAND2XL U19235 ( .A(B6_q[14]), .B(n16570), .Y(n15308) );
  NAND2XL U19236 ( .A(B4_q[14]), .B(n7126), .Y(n15307) );
  NAND4XL U19237 ( .A(n15919), .B(n15918), .C(n5800), .D(n15917), .Y(n15920)
         );
  NAND2XL U19238 ( .A(B4_q[15]), .B(n15969), .Y(n15919) );
  NAND2XL U19239 ( .A(B5_q[15]), .B(n15963), .Y(n15918) );
  NAND4XL U19240 ( .A(n15713), .B(n15712), .C(n5800), .D(n15711), .Y(n15714)
         );
  NAND2XL U19241 ( .A(B7_q[15]), .B(n16325), .Y(n15713) );
  NAND2XL U19242 ( .A(B5_q[15]), .B(n15747), .Y(n15712) );
  NAND4XL U19243 ( .A(n15301), .B(n15300), .C(n5917), .D(n15299), .Y(n15302)
         );
  NAND2XL U19244 ( .A(B4_q[15]), .B(n7126), .Y(n15301) );
  NAND2XL U19245 ( .A(B5_q[15]), .B(n16559), .Y(n15300) );
  NAND4XL U19246 ( .A(n15518), .B(n15517), .C(n5905), .D(n15516), .Y(n15519)
         );
  NAND2XL U19247 ( .A(B7_q[16]), .B(n16158), .Y(n15518) );
  NAND2XL U19248 ( .A(B4_q[16]), .B(n15557), .Y(n15517) );
  NAND4XL U19249 ( .A(n15294), .B(n15293), .C(n5800), .D(n15292), .Y(n15295)
         );
  NAND2XL U19250 ( .A(B5_q[16]), .B(n16375), .Y(n15294) );
  NAND2XL U19251 ( .A(B4_q[16]), .B(n7126), .Y(n15293) );
  NAND4XL U19252 ( .A(n15911), .B(n15910), .C(n5800), .D(n15909), .Y(n15912)
         );
  NAND2XL U19253 ( .A(B6_q[17]), .B(n15958), .Y(n15911) );
  NAND2XL U19254 ( .A(B5_q[17]), .B(n15963), .Y(n15910) );
  NAND4XL U19255 ( .A(n15705), .B(n15704), .C(n5800), .D(n15703), .Y(n15706)
         );
  NAND2XL U19256 ( .A(B6_q[17]), .B(n5926), .Y(n15705) );
  NAND2XL U19257 ( .A(B5_q[17]), .B(n15747), .Y(n15704) );
  NAND4XL U19258 ( .A(n15514), .B(n15513), .C(n5907), .D(n15512), .Y(n15515)
         );
  NAND2XL U19259 ( .A(B7_q[17]), .B(n16158), .Y(n15514) );
  NAND2XL U19260 ( .A(B5_q[17]), .B(n5931), .Y(n15513) );
  NAND4XL U19261 ( .A(n15286), .B(n15285), .C(n5907), .D(n15284), .Y(n15287)
         );
  NAND2XL U19262 ( .A(B4_q[17]), .B(n7126), .Y(n15286) );
  NAND2XL U19263 ( .A(B5_q[17]), .B(n16559), .Y(n15285) );
  OAI211XL U19264 ( .A0(n15967), .A1(n15907), .B0(n15906), .C0(n15905), .Y(
        n15908) );
  AOI21XL U19265 ( .A0(B5_q[18]), .A1(n15963), .B0(n16564), .Y(n15905) );
  AOI22XL U19266 ( .A0(B6_q[18]), .A1(n15958), .B0(B4_q[18]), .B1(n5925), .Y(
        n15906) );
  OAI211XL U19267 ( .A0(n5806), .A1(n15701), .B0(n15510), .C0(n15509), .Y(
        n15511) );
  AOI22XL U19268 ( .A0(B6_q[18]), .A1(n16143), .B0(B7_q[18]), .B1(n16128), .Y(
        n15510) );
  AOI21XL U19269 ( .A0(B4_q[18]), .A1(n5933), .B0(n28985), .Y(n15509) );
  OAI211XL U19270 ( .A0(n5799), .A1(n15701), .B0(n15279), .C0(n15278), .Y(
        n15280) );
  AOI21XL U19271 ( .A0(B4_q[18]), .A1(n7126), .B0(n16496), .Y(n15278) );
  AOI22XL U19272 ( .A0(B7_q[18]), .A1(n7127), .B0(B6_q[18]), .B1(n16570), .Y(
        n15279) );
  NAND4XL U19273 ( .A(n15903), .B(n15902), .C(n5905), .D(n15901), .Y(n15904)
         );
  NAND2XL U19274 ( .A(B4_q[19]), .B(n5925), .Y(n15903) );
  NAND2XL U19275 ( .A(B5_q[19]), .B(n15963), .Y(n15902) );
  NAND4XL U19276 ( .A(n15507), .B(n15506), .C(n5905), .D(n15505), .Y(n15508)
         );
  NAND2XL U19277 ( .A(B6_q[19]), .B(n15431), .Y(n15507) );
  NAND2XL U19278 ( .A(B4_q[19]), .B(n15557), .Y(n15506) );
  NAND4XL U19279 ( .A(n15272), .B(n15271), .C(n5800), .D(n15270), .Y(n15273)
         );
  NAND2XL U19280 ( .A(B7_q[19]), .B(n16569), .Y(n15272) );
  NAND2XL U19281 ( .A(B4_q[19]), .B(n7126), .Y(n15271) );
  OAI211XL U19282 ( .A0(n5836), .A1(n15980), .B0(n15979), .C0(n15978), .Y(
        n15981) );
  AOI21XL U19283 ( .A0(B4_q[1]), .A1(n5925), .B0(n5924), .Y(n15978) );
  AOI22XL U19284 ( .A0(B7_q[1]), .A1(n15982), .B0(B6_q[1]), .B1(n15958), .Y(
        n15979) );
  OAI211XL U19285 ( .A0(n15980), .A1(n5813), .B0(n15768), .C0(n15767), .Y(
        n15769) );
  AOI22XL U19286 ( .A0(B7_q[1]), .A1(n16325), .B0(B6_q[1]), .B1(n16354), .Y(
        n15768) );
  AOI21XL U19287 ( .A0(B4_q[1]), .A1(n15687), .B0(n28985), .Y(n15767) );
  OAI211XL U19288 ( .A0(n5841), .A1(n15574), .B0(n15573), .C0(n15572), .Y(
        n15575) );
  AOI21XL U19289 ( .A0(B5_q[1]), .A1(n16165), .B0(n5924), .Y(n15572) );
  AOI22XL U19290 ( .A0(B6_q[1]), .A1(n16143), .B0(B4_q[1]), .B1(n15557), .Y(
        n15573) );
  OAI211XL U19291 ( .A0(n5836), .A1(n15899), .B0(n15898), .C0(n15897), .Y(
        n15900) );
  AOI22XL U19292 ( .A0(B7_q[20]), .A1(n15982), .B0(B4_q[20]), .B1(n5925), .Y(
        n15898) );
  OAI211XL U19293 ( .A0(n5813), .A1(n15899), .B0(n15693), .C0(n15692), .Y(
        n15694) );
  AOI21XL U19294 ( .A0(B4_q[20]), .A1(n15687), .B0(n5924), .Y(n15692) );
  AOI22XL U19295 ( .A0(B7_q[20]), .A1(n16325), .B0(B6_q[20]), .B1(n16354), .Y(
        n15693) );
  OAI211XL U19296 ( .A0(n15495), .A1(n15503), .B0(n15502), .C0(n15501), .Y(
        n15504) );
  AOI22XL U19297 ( .A0(B7_q[20]), .A1(n16128), .B0(B5_q[20]), .B1(n16165), .Y(
        n15502) );
  AOI21XL U19298 ( .A0(B4_q[20]), .A1(n5933), .B0(n28985), .Y(n15501) );
  OAI211XL U19299 ( .A0(n15264), .A1(n5914), .B0(n15263), .C0(n15262), .Y(
        n15265) );
  AOI21XL U19300 ( .A0(B5_q[20]), .A1(n16559), .B0(n28985), .Y(n15262) );
  AOI22XL U19301 ( .A0(B7_q[20]), .A1(n7127), .B0(B6_q[20]), .B1(n16570), .Y(
        n15263) );
  NAND4XL U19302 ( .A(n15895), .B(n15894), .C(n5917), .D(n15893), .Y(n15896)
         );
  NAND2XL U19303 ( .A(B6_q[21]), .B(n15958), .Y(n15895) );
  NAND2XL U19304 ( .A(B5_q[21]), .B(n15963), .Y(n15894) );
  NAND4XL U19305 ( .A(n15690), .B(n15689), .C(n5913), .D(n15688), .Y(n15691)
         );
  NAND2XL U19306 ( .A(B4_q[21]), .B(n15687), .Y(n15690) );
  NAND2XL U19307 ( .A(B5_q[21]), .B(n15747), .Y(n15689) );
  NAND4XL U19308 ( .A(n15499), .B(n15498), .C(n5909), .D(n15497), .Y(n15500)
         );
  NAND2XL U19309 ( .A(B7_q[21]), .B(n16158), .Y(n15499) );
  NAND2XL U19310 ( .A(B4_q[21]), .B(n5933), .Y(n15498) );
  NAND4XL U19311 ( .A(n15256), .B(n15255), .C(n5908), .D(n15254), .Y(n15257)
         );
  NAND2XL U19312 ( .A(B6_q[21]), .B(n16570), .Y(n15256) );
  NAND2XL U19313 ( .A(B4_q[21]), .B(n7126), .Y(n15255) );
  OAI211XL U19314 ( .A0(n5836), .A1(n15891), .B0(n15890), .C0(n15889), .Y(
        n15892) );
  AOI21XL U19315 ( .A0(B4_q[22]), .A1(n15969), .B0(n5924), .Y(n15889) );
  AOI22XL U19316 ( .A0(B6_q[22]), .A1(n15958), .B0(B7_q[22]), .B1(n15982), .Y(
        n15890) );
  OAI211XL U19317 ( .A0(n15633), .A1(n15685), .B0(n15684), .C0(n15683), .Y(
        n15686) );
  AOI21XL U19318 ( .A0(B4_q[22]), .A1(n15687), .B0(n5924), .Y(n15683) );
  AOI22XL U19319 ( .A0(B7_q[22]), .A1(n16325), .B0(B5_q[22]), .B1(n16344), .Y(
        n15684) );
  OAI211XL U19320 ( .A0(n15495), .A1(n15685), .B0(n15494), .C0(n15493), .Y(
        n15496) );
  AOI21XL U19321 ( .A0(B4_q[22]), .A1(n5933), .B0(n5924), .Y(n15493) );
  AOI22XL U19322 ( .A0(B7_q[22]), .A1(n16128), .B0(B5_q[22]), .B1(n16165), .Y(
        n15494) );
  OAI211XL U19323 ( .A0(n15248), .A1(n5914), .B0(n15247), .C0(n15246), .Y(
        n15249) );
  AOI21XL U19324 ( .A0(B5_q[22]), .A1(n16559), .B0(n5924), .Y(n15246) );
  AOI22XL U19325 ( .A0(B7_q[22]), .A1(n7127), .B0(B6_q[22]), .B1(n16570), .Y(
        n15247) );
  NAND4XL U19326 ( .A(n15887), .B(n15886), .C(n5905), .D(n15885), .Y(n15888)
         );
  NAND2XL U19327 ( .A(B7_q[23]), .B(n5930), .Y(n15887) );
  NAND2XL U19328 ( .A(B4_q[23]), .B(n5925), .Y(n15886) );
  NAND4XL U19329 ( .A(n15681), .B(n15680), .C(n5908), .D(n15679), .Y(n15682)
         );
  NAND2XL U19330 ( .A(B4_q[23]), .B(n16277), .Y(n15681) );
  NAND2XL U19331 ( .A(B6_q[23]), .B(n16293), .Y(n15680) );
  NAND4XL U19332 ( .A(n15491), .B(n15490), .C(n5909), .D(n15489), .Y(n15492)
         );
  NAND2XL U19333 ( .A(B4_q[23]), .B(n5933), .Y(n15491) );
  NAND2XL U19334 ( .A(B6_q[23]), .B(n16143), .Y(n15490) );
  NAND4XL U19335 ( .A(n15241), .B(n15240), .C(R7_valid), .D(n15239), .Y(n15242) );
  NAND2XL U19336 ( .A(B5_q[23]), .B(n16375), .Y(n15241) );
  NAND2XL U19337 ( .A(B4_q[23]), .B(n7126), .Y(n15240) );
  OAI211XL U19338 ( .A0(n5836), .A1(n15883), .B0(n15882), .C0(n15881), .Y(
        n15884) );
  AOI21XL U19339 ( .A0(B4_q[24]), .A1(n15969), .B0(n5924), .Y(n15881) );
  AOI22XL U19340 ( .A0(B7_q[24]), .A1(n15982), .B0(B6_q[24]), .B1(n15958), .Y(
        n15882) );
  OAI211XL U19341 ( .A0(n5813), .A1(n15883), .B0(n15677), .C0(n15676), .Y(
        n15678) );
  AOI21XL U19342 ( .A0(B4_q[24]), .A1(n15687), .B0(n5924), .Y(n15676) );
  AOI22XL U19343 ( .A0(B7_q[24]), .A1(n16325), .B0(B6_q[24]), .B1(n5926), .Y(
        n15677) );
  OAI211XL U19344 ( .A0(n5806), .A1(n15883), .B0(n15487), .C0(n15486), .Y(
        n15488) );
  AOI21XL U19345 ( .A0(B6_q[24]), .A1(n16161), .B0(n5807), .Y(n15486) );
  AOI22XL U19346 ( .A0(B7_q[24]), .A1(n16128), .B0(B4_q[24]), .B1(n15557), .Y(
        n15487) );
  OAI211XL U19347 ( .A0(n5799), .A1(n15883), .B0(n15234), .C0(n15233), .Y(
        n15235) );
  AOI21XL U19348 ( .A0(B6_q[24]), .A1(n16570), .B0(n28985), .Y(n15233) );
  AOI22XL U19349 ( .A0(B4_q[24]), .A1(n7126), .B0(B7_q[24]), .B1(n7127), .Y(
        n15234) );
  OAI211XL U19350 ( .A0(n5836), .A1(n15879), .B0(n15878), .C0(n15877), .Y(
        n15880) );
  AOI21XL U19351 ( .A0(B4_q[25]), .A1(n5925), .B0(n16470), .Y(n15877) );
  AOI22XL U19352 ( .A0(B6_q[25]), .A1(n15958), .B0(B7_q[25]), .B1(n15982), .Y(
        n15878) );
  OAI211XL U19353 ( .A0(n5813), .A1(n15879), .B0(n15674), .C0(n15673), .Y(
        n15675) );
  AOI21XL U19354 ( .A0(B7_q[25]), .A1(n16325), .B0(n5924), .Y(n15673) );
  AOI22XL U19355 ( .A0(B6_q[25]), .A1(n5926), .B0(B4_q[25]), .B1(n15687), .Y(
        n15674) );
  OAI211XL U19356 ( .A0(n5841), .A1(n15484), .B0(n15483), .C0(n15482), .Y(
        n15485) );
  AOI22XL U19357 ( .A0(B6_q[25]), .A1(n16143), .B0(B4_q[25]), .B1(n15557), .Y(
        n15483) );
  OAI211XL U19358 ( .A0(n5799), .A1(n15879), .B0(n15227), .C0(n15226), .Y(
        n15228) );
  AOI21XL U19359 ( .A0(B7_q[25]), .A1(n7127), .B0(n28985), .Y(n15226) );
  AOI22XL U19360 ( .A0(B4_q[25]), .A1(n7126), .B0(B6_q[25]), .B1(n16570), .Y(
        n15227) );
  OAI211XL U19361 ( .A0(n5836), .A1(n15875), .B0(n15874), .C0(n15873), .Y(
        n15876) );
  AOI21XL U19362 ( .A0(B6_q[26]), .A1(n15958), .B0(n5924), .Y(n15873) );
  AOI22XL U19363 ( .A0(B4_q[26]), .A1(n5925), .B0(B7_q[26]), .B1(n5930), .Y(
        n15874) );
  OAI211XL U19364 ( .A0(n5813), .A1(n15875), .B0(n15671), .C0(n15670), .Y(
        n15672) );
  AOI21XL U19365 ( .A0(B6_q[26]), .A1(n5926), .B0(n5924), .Y(n15670) );
  AOI22XL U19366 ( .A0(B4_q[26]), .A1(n15687), .B0(B7_q[26]), .B1(n16325), .Y(
        n15671) );
  OAI211XL U19367 ( .A0(n5841), .A1(n15480), .B0(n15479), .C0(n15478), .Y(
        n15481) );
  AOI22XL U19368 ( .A0(B6_q[26]), .A1(n16143), .B0(B4_q[26]), .B1(n15557), .Y(
        n15479) );
  AOI21XL U19369 ( .A0(B5_q[26]), .A1(n5931), .B0(n28985), .Y(n15478) );
  OAI211XL U19370 ( .A0(n5799), .A1(n15875), .B0(n15021), .C0(n15020), .Y(
        n15022) );
  AOI21XL U19371 ( .A0(B7_q[26]), .A1(n16569), .B0(n16496), .Y(n15020) );
  AOI22XL U19372 ( .A0(B4_q[26]), .A1(n7126), .B0(B6_q[26]), .B1(n16570), .Y(
        n15021) );
  NAND4XL U19373 ( .A(n15476), .B(n15475), .C(n5915), .D(n15474), .Y(n15477)
         );
  NAND2XL U19374 ( .A(B5_q[27]), .B(n16165), .Y(n15476) );
  NAND2XL U19375 ( .A(B4_q[27]), .B(n15557), .Y(n15475) );
  NAND4XL U19376 ( .A(n15001), .B(n15000), .C(R7_valid), .D(n14999), .Y(n15002) );
  NAND2XL U19377 ( .A(B7_q[27]), .B(n7127), .Y(n15001) );
  NAND2XL U19378 ( .A(B4_q[27]), .B(n7126), .Y(n15000) );
  OAI211XL U19379 ( .A0(n5836), .A1(n15867), .B0(n15866), .C0(n15865), .Y(
        n15868) );
  AOI21XL U19380 ( .A0(B4_q[28]), .A1(n5925), .B0(n5924), .Y(n15865) );
  AOI22XL U19381 ( .A0(B7_q[28]), .A1(n15982), .B0(B6_q[28]), .B1(n15958), .Y(
        n15866) );
  OAI211XL U19382 ( .A0(n5841), .A1(n15664), .B0(n15472), .C0(n15471), .Y(
        n15473) );
  AOI22XL U19383 ( .A0(B6_q[28]), .A1(n16143), .B0(B5_q[28]), .B1(n16165), .Y(
        n15472) );
  AOI21XL U19384 ( .A0(B4_q[28]), .A1(n5933), .B0(n28985), .Y(n15471) );
  OAI211XL U19385 ( .A0(n15036), .A1(n5914), .B0(n15035), .C0(n15034), .Y(
        n15037) );
  AOI21XL U19386 ( .A0(B5_q[28]), .A1(n16375), .B0(n16496), .Y(n15034) );
  AOI22XL U19387 ( .A0(B7_q[28]), .A1(n7127), .B0(B6_q[28]), .B1(n16570), .Y(
        n15035) );
  NAND4XL U19388 ( .A(n15469), .B(n15468), .C(n5909), .D(n15467), .Y(n15470)
         );
  NAND2XL U19389 ( .A(B6_q[29]), .B(n16143), .Y(n15469) );
  NAND2XL U19390 ( .A(B4_q[29]), .B(n5933), .Y(n15468) );
  NAND4XL U19391 ( .A(n15373), .B(n15372), .C(n5913), .D(n15371), .Y(n15374)
         );
  NAND2XL U19392 ( .A(B5_q[29]), .B(n16375), .Y(n15373) );
  NAND2XL U19393 ( .A(B4_q[29]), .B(n7126), .Y(n15372) );
  NAND4XL U19394 ( .A(n15976), .B(n15975), .C(n5906), .D(n15974), .Y(n15977)
         );
  NAND2XL U19395 ( .A(B4_q[2]), .B(n5925), .Y(n15976) );
  NAND2XL U19396 ( .A(B5_q[2]), .B(n15963), .Y(n15975) );
  NAND4XL U19397 ( .A(n15765), .B(n15764), .C(n5910), .D(n15763), .Y(n15766)
         );
  NAND2XL U19398 ( .A(B7_q[2]), .B(n16325), .Y(n15765) );
  NAND2XL U19399 ( .A(B5_q[2]), .B(n16344), .Y(n15764) );
  NAND4XL U19400 ( .A(n15570), .B(n15569), .C(n5912), .D(n15568), .Y(n15571)
         );
  NAND2XL U19401 ( .A(B6_q[2]), .B(n16143), .Y(n15570) );
  NAND2XL U19402 ( .A(B5_q[2]), .B(n16165), .Y(n15569) );
  OAI211XL U19403 ( .A0(n5799), .A1(n15855), .B0(n15359), .C0(n15358), .Y(
        n15360) );
  AOI21XL U19404 ( .A0(B6_q[31]), .A1(n16570), .B0(n16496), .Y(n15358) );
  AOI22XL U19405 ( .A0(B4_q[31]), .A1(n7126), .B0(B7_q[31]), .B1(n7127), .Y(
        n15359) );
  OAI211XL U19406 ( .A0(n5799), .A1(n15650), .B0(n15018), .C0(n15017), .Y(
        n15019) );
  AOI21XL U19407 ( .A0(B7_q[32]), .A1(n16569), .B0(n15349), .Y(n15017) );
  AOI22XL U19408 ( .A0(B4_q[32]), .A1(n7126), .B0(B6_q[32]), .B1(n16570), .Y(
        n15018) );
  OAI211XL U19409 ( .A0(n5806), .A1(n15847), .B0(n15456), .C0(n15455), .Y(
        n15457) );
  AOI22XL U19410 ( .A0(B7_q[33]), .A1(n16128), .B0(B6_q[33]), .B1(n16143), .Y(
        n15456) );
  AOI21XL U19411 ( .A0(B4_q[33]), .A1(n5933), .B0(n28985), .Y(n15455) );
  OAI211XL U19412 ( .A0(n5799), .A1(n15847), .B0(n15007), .C0(n15006), .Y(
        n15008) );
  AOI21XL U19413 ( .A0(B4_q[33]), .A1(n7126), .B0(n15349), .Y(n15006) );
  AOI22XL U19414 ( .A0(B7_q[33]), .A1(n7127), .B0(B6_q[33]), .B1(n16570), .Y(
        n15007) );
  OAI211XL U19415 ( .A0(n5836), .A1(n15843), .B0(n15842), .C0(n15841), .Y(
        n15844) );
  AOI21XL U19416 ( .A0(B4_q[34]), .A1(n5925), .B0(n16487), .Y(n15841) );
  AOI22XL U19417 ( .A0(B6_q[34]), .A1(n15958), .B0(B7_q[34]), .B1(n5930), .Y(
        n15842) );
  OAI211XL U19418 ( .A0(n15643), .A1(n15633), .B0(n15642), .C0(n15641), .Y(
        n15644) );
  AOI22XL U19419 ( .A0(B7_q[34]), .A1(n16325), .B0(B5_q[34]), .B1(n16344), .Y(
        n15642) );
  OAI211XL U19420 ( .A0(n5806), .A1(n15843), .B0(n15453), .C0(n15452), .Y(
        n15454) );
  AOI21XL U19421 ( .A0(B4_q[34]), .A1(n5933), .B0(n5924), .Y(n15452) );
  AOI22XL U19422 ( .A0(B6_q[34]), .A1(n16143), .B0(B7_q[34]), .B1(n16128), .Y(
        n15453) );
  OAI211XL U19423 ( .A0(n15015), .A1(n5914), .B0(n15014), .C0(n15013), .Y(
        n15016) );
  AOI21XL U19424 ( .A0(B5_q[34]), .A1(n16375), .B0(n5924), .Y(n15013) );
  AOI22XL U19425 ( .A0(B7_q[34]), .A1(n7127), .B0(B6_q[34]), .B1(n16570), .Y(
        n15014) );
  NAND4XL U19426 ( .A(n15839), .B(n15838), .C(n6880), .D(n15837), .Y(n15840)
         );
  NAND2XL U19427 ( .A(B7_q[35]), .B(n15982), .Y(n15839) );
  NAND2XL U19428 ( .A(B5_q[35]), .B(n15963), .Y(n15838) );
  NAND4XL U19429 ( .A(n15450), .B(n15449), .C(n5915), .D(n15448), .Y(n15451)
         );
  NAND2XL U19430 ( .A(B4_q[35]), .B(n5933), .Y(n15450) );
  NAND2XL U19431 ( .A(B5_q[35]), .B(n16165), .Y(n15449) );
  NAND4XL U19432 ( .A(n15831), .B(n15830), .C(n5915), .D(n15829), .Y(n15832)
         );
  NAND2XL U19433 ( .A(B6_q[37]), .B(n15958), .Y(n15831) );
  NAND2XL U19434 ( .A(B5_q[37]), .B(n15963), .Y(n15830) );
  NAND4XL U19435 ( .A(n15827), .B(n15826), .C(n5909), .D(n15825), .Y(n15828)
         );
  NAND2XL U19436 ( .A(B4_q[38]), .B(n5925), .Y(n15827) );
  NAND2XL U19437 ( .A(B5_q[38]), .B(n15963), .Y(n15826) );
  NAND4XL U19438 ( .A(n15438), .B(n15437), .C(n5915), .D(n15436), .Y(n15439)
         );
  NAND2XL U19439 ( .A(B4_q[38]), .B(n15557), .Y(n15438) );
  NAND2XL U19440 ( .A(B5_q[38]), .B(n16165), .Y(n15437) );
  NAND4XL U19441 ( .A(n15320), .B(n15319), .C(n5909), .D(n15318), .Y(n15321)
         );
  NAND2XL U19442 ( .A(B7_q[38]), .B(n16569), .Y(n15320) );
  NAND2XL U19443 ( .A(B4_q[38]), .B(n7126), .Y(n15319) );
  OAI211XL U19444 ( .A0(n5836), .A1(n15823), .B0(n15822), .C0(n15821), .Y(
        n15824) );
  AOI21XL U19445 ( .A0(B4_q[39]), .A1(n5925), .B0(n16496), .Y(n15821) );
  AOI22XL U19446 ( .A0(B7_q[39]), .A1(n15982), .B0(B6_q[39]), .B1(n15958), .Y(
        n15822) );
  OAI211XL U19447 ( .A0(n15495), .A1(n15434), .B0(n15433), .C0(n15432), .Y(
        n15435) );
  AOI21XL U19448 ( .A0(B4_q[39]), .A1(n5933), .B0(n5924), .Y(n15432) );
  AOI22XL U19449 ( .A0(B7_q[39]), .A1(n16128), .B0(B5_q[39]), .B1(n16165), .Y(
        n15433) );
  OAI211XL U19450 ( .A0(n15312), .A1(n5914), .B0(n15311), .C0(n15310), .Y(
        n15313) );
  AOI21XL U19451 ( .A0(B6_q[39]), .A1(n16570), .B0(n5924), .Y(n15310) );
  AOI22XL U19452 ( .A0(B7_q[39]), .A1(n7127), .B0(B5_q[39]), .B1(n16559), .Y(
        n15311) );
  OAI211XL U19453 ( .A0(n5836), .A1(n15972), .B0(n15971), .C0(n15970), .Y(
        n15973) );
  AOI21XL U19454 ( .A0(B4_q[3]), .A1(n15969), .B0(n5924), .Y(n15970) );
  AOI22XL U19455 ( .A0(B6_q[3]), .A1(n15958), .B0(B7_q[3]), .B1(n15982), .Y(
        n15971) );
  OAI211XL U19456 ( .A0(n5806), .A1(n15972), .B0(n15566), .C0(n15565), .Y(
        n15567) );
  AOI21XL U19457 ( .A0(B4_q[3]), .A1(n5933), .B0(n5924), .Y(n15565) );
  AOI22XL U19458 ( .A0(B6_q[3]), .A1(n16143), .B0(B7_q[3]), .B1(n16128), .Y(
        n15566) );
  OAI211XL U19459 ( .A0(n5836), .A1(n15815), .B0(n15814), .C0(n15813), .Y(
        n15816) );
  AOI22XL U19460 ( .A0(B7_q[41]), .A1(n5930), .B0(B6_q[41]), .B1(n15958), .Y(
        n15814) );
  AOI21XL U19461 ( .A0(B4_q[41]), .A1(n5925), .B0(n28985), .Y(n15813) );
  NAND4XL U19462 ( .A(n15811), .B(n15810), .C(n5915), .D(n15809), .Y(n15812)
         );
  NAND2XL U19463 ( .A(B6_q[42]), .B(n15958), .Y(n15811) );
  NAND2XL U19464 ( .A(B5_q[42]), .B(n15963), .Y(n15810) );
  NAND4XL U19465 ( .A(n15614), .B(n15613), .C(n5909), .D(n15612), .Y(n15615)
         );
  NAND2XL U19466 ( .A(B7_q[42]), .B(n16325), .Y(n15614) );
  NAND2XL U19467 ( .A(B5_q[42]), .B(n15747), .Y(n15613) );
  NAND4XL U19468 ( .A(n15423), .B(n15422), .C(n5915), .D(n15421), .Y(n15424)
         );
  NAND2XL U19469 ( .A(B4_q[42]), .B(n15557), .Y(n15423) );
  NAND2XL U19470 ( .A(B5_q[42]), .B(n16165), .Y(n15422) );
  OAI211XL U19471 ( .A0(n5836), .A1(n15807), .B0(n15806), .C0(n15805), .Y(
        n15808) );
  AOI21XL U19472 ( .A0(B4_q[43]), .A1(n5925), .B0(n5807), .Y(n15805) );
  AOI22XL U19473 ( .A0(B6_q[43]), .A1(n15958), .B0(B7_q[43]), .B1(n5930), .Y(
        n15806) );
  OAI211XL U19474 ( .A0(n5806), .A1(n15807), .B0(n15419), .C0(n15418), .Y(
        n15420) );
  AOI21XL U19475 ( .A0(B4_q[43]), .A1(n5933), .B0(n16461), .Y(n15418) );
  AOI22XL U19476 ( .A0(B6_q[43]), .A1(n16143), .B0(B7_q[43]), .B1(n16128), .Y(
        n15419) );
  OAI211XL U19477 ( .A0(n5799), .A1(n15807), .B0(n15282), .C0(n15281), .Y(
        n15283) );
  AOI21XL U19478 ( .A0(B7_q[43]), .A1(n16569), .B0(n28985), .Y(n15281) );
  AOI22XL U19479 ( .A0(B4_q[43]), .A1(n7126), .B0(B6_q[43]), .B1(n16570), .Y(
        n15282) );
  NAND4XL U19480 ( .A(n15803), .B(n15802), .C(n5909), .D(n15801), .Y(n15804)
         );
  NAND2XL U19481 ( .A(B4_q[44]), .B(n15969), .Y(n15803) );
  NAND2XL U19482 ( .A(B5_q[44]), .B(n15963), .Y(n15802) );
  NAND4XL U19483 ( .A(n15416), .B(n15415), .C(n5909), .D(n15414), .Y(n15417)
         );
  NAND2XL U19484 ( .A(B5_q[44]), .B(n16165), .Y(n15416) );
  NAND2XL U19485 ( .A(B7_q[44]), .B(n16158), .Y(n15415) );
  NAND4XL U19486 ( .A(n15276), .B(n15275), .C(n5915), .D(n15274), .Y(n15277)
         );
  NAND2XL U19487 ( .A(B6_q[44]), .B(n16570), .Y(n15276) );
  NAND2XL U19488 ( .A(B5_q[44]), .B(n16559), .Y(n15275) );
  NAND4XL U19489 ( .A(n15795), .B(n15794), .C(n5915), .D(n15793), .Y(n15796)
         );
  NAND2XL U19490 ( .A(B4_q[46]), .B(n15969), .Y(n15795) );
  NAND2XL U19491 ( .A(B5_q[46]), .B(n15963), .Y(n15794) );
  NAND4XL U19492 ( .A(n15599), .B(n15598), .C(n5915), .D(n15597), .Y(n15600)
         );
  NAND2XL U19493 ( .A(B6_q[46]), .B(n5926), .Y(n15599) );
  NAND2XL U19494 ( .A(B4_q[46]), .B(n16277), .Y(n15598) );
  NAND4XL U19495 ( .A(n15409), .B(n15408), .C(n5915), .D(n15407), .Y(n15410)
         );
  NAND2XL U19496 ( .A(B4_q[46]), .B(n15557), .Y(n15409) );
  NAND2XL U19497 ( .A(B5_q[46]), .B(n16165), .Y(n15408) );
  OAI211XL U19498 ( .A0(n15967), .A1(n15791), .B0(n15790), .C0(n15789), .Y(
        n15792) );
  AOI21XL U19499 ( .A0(B4_q[47]), .A1(n5925), .B0(n16487), .Y(n15789) );
  AOI22XL U19500 ( .A0(B6_q[47]), .A1(n15958), .B0(B5_q[47]), .B1(n15963), .Y(
        n15790) );
  OAI211XL U19501 ( .A0(n5813), .A1(n15595), .B0(n15594), .C0(n15593), .Y(
        n15596) );
  AOI21XL U19502 ( .A0(B4_q[47]), .A1(n16277), .B0(n16496), .Y(n15593) );
  AOI22XL U19503 ( .A0(B7_q[47]), .A1(n16325), .B0(B6_q[47]), .B1(n16354), .Y(
        n15594) );
  OAI211XL U19504 ( .A0(n5841), .A1(n15791), .B0(n15405), .C0(n15404), .Y(
        n15406) );
  AOI21XL U19505 ( .A0(B4_q[47]), .A1(n5933), .B0(n5924), .Y(n15404) );
  AOI22XL U19506 ( .A0(B6_q[47]), .A1(n16143), .B0(B5_q[47]), .B1(n16165), .Y(
        n15405) );
  OAI211XL U19507 ( .A0(n5836), .A1(n15787), .B0(n15786), .C0(n15785), .Y(
        n15788) );
  AOI21XL U19508 ( .A0(B6_q[48]), .A1(n15958), .B0(n16461), .Y(n15785) );
  AOI22XL U19509 ( .A0(B4_q[48]), .A1(n5925), .B0(B7_q[48]), .B1(n15982), .Y(
        n15786) );
  OAI211XL U19510 ( .A0(n5813), .A1(n15787), .B0(n15591), .C0(n15590), .Y(
        n15592) );
  AOI21XL U19511 ( .A0(B6_q[48]), .A1(n5926), .B0(n16501), .Y(n15590) );
  AOI22XL U19512 ( .A0(B4_q[48]), .A1(n15687), .B0(B7_q[48]), .B1(n16325), .Y(
        n15591) );
  OAI211XL U19513 ( .A0(n5841), .A1(n15402), .B0(n15401), .C0(n15400), .Y(
        n15403) );
  AOI21XL U19514 ( .A0(B5_q[48]), .A1(n16165), .B0(n16564), .Y(n15400) );
  AOI22XL U19515 ( .A0(B4_q[48]), .A1(n15557), .B0(B6_q[48]), .B1(n16143), .Y(
        n15401) );
  OAI211XL U19516 ( .A0(n5799), .A1(n15787), .B0(n15244), .C0(n15243), .Y(
        n15245) );
  AOI21XL U19517 ( .A0(B7_q[48]), .A1(n7127), .B0(n15349), .Y(n15243) );
  AOI22XL U19518 ( .A0(B4_q[48]), .A1(n7126), .B0(B6_q[48]), .B1(n16570), .Y(
        n15244) );
  OAI211XL U19519 ( .A0(n5836), .A1(n15783), .B0(n15782), .C0(n15781), .Y(
        n15784) );
  AOI21XL U19520 ( .A0(B4_q[49]), .A1(n5925), .B0(n16461), .Y(n15781) );
  AOI22XL U19521 ( .A0(B7_q[49]), .A1(n15982), .B0(B6_q[49]), .B1(n15958), .Y(
        n15782) );
  OAI211XL U19522 ( .A0(n5813), .A1(n15783), .B0(n15588), .C0(n15587), .Y(
        n15589) );
  AOI21XL U19523 ( .A0(B7_q[49]), .A1(n16325), .B0(n16501), .Y(n15587) );
  AOI22XL U19524 ( .A0(B6_q[49]), .A1(n16293), .B0(B4_q[49]), .B1(n15687), .Y(
        n15588) );
  OAI211XL U19525 ( .A0(n5841), .A1(n15398), .B0(n15397), .C0(n15396), .Y(
        n15399) );
  AOI22XL U19526 ( .A0(B6_q[49]), .A1(n16143), .B0(B4_q[49]), .B1(n15557), .Y(
        n15397) );
  OAI211XL U19527 ( .A0(n5799), .A1(n15783), .B0(n15237), .C0(n15236), .Y(
        n15238) );
  AOI21XL U19528 ( .A0(B4_q[49]), .A1(n7126), .B0(n28985), .Y(n15236) );
  AOI22XL U19529 ( .A0(B7_q[49]), .A1(n7127), .B0(B6_q[49]), .B1(n16570), .Y(
        n15237) );
  OAI211XL U19530 ( .A0(n5813), .A1(n15758), .B0(n15757), .C0(n15756), .Y(
        n15759) );
  AOI21XL U19531 ( .A0(B7_q[4]), .A1(n16325), .B0(n16470), .Y(n15756) );
  AOI22XL U19532 ( .A0(B6_q[4]), .A1(n16354), .B0(B4_q[4]), .B1(n15687), .Y(
        n15757) );
  OAI211XL U19533 ( .A0(n5841), .A1(n15966), .B0(n15563), .C0(n15562), .Y(
        n15564) );
  AOI21XL U19534 ( .A0(B5_q[4]), .A1(n5931), .B0(n5924), .Y(n15562) );
  AOI22XL U19535 ( .A0(B6_q[4]), .A1(n16143), .B0(B4_q[4]), .B1(n15557), .Y(
        n15563) );
  NAND4XL U19536 ( .A(n15779), .B(n15778), .C(n5915), .D(n15777), .Y(n15780)
         );
  NAND2XL U19537 ( .A(B7_q[50]), .B(n15982), .Y(n15779) );
  NAND2XL U19538 ( .A(B5_q[50]), .B(n15963), .Y(n15778) );
  NAND4XL U19539 ( .A(n15585), .B(n15584), .C(n5909), .D(n15583), .Y(n15586)
         );
  NAND2XL U19540 ( .A(B6_q[50]), .B(n16293), .Y(n15585) );
  NAND2XL U19541 ( .A(B5_q[50]), .B(n15747), .Y(n15584) );
  NAND4XL U19542 ( .A(n15394), .B(n15393), .C(n5915), .D(n15392), .Y(n15395)
         );
  NAND2XL U19543 ( .A(B6_q[50]), .B(n16161), .Y(n15394) );
  NAND2XL U19544 ( .A(B5_q[50]), .B(n16165), .Y(n15393) );
  NAND4XL U19545 ( .A(n15231), .B(n15230), .C(n5915), .D(n15229), .Y(n15232)
         );
  NAND2XL U19546 ( .A(B4_q[50]), .B(n7126), .Y(n15231) );
  NAND2XL U19547 ( .A(B5_q[50]), .B(n16375), .Y(n15230) );
  OAI211XL U19548 ( .A0(n5836), .A1(n15775), .B0(n15774), .C0(n15773), .Y(
        n15776) );
  AOI21XL U19549 ( .A0(B4_q[51]), .A1(n5925), .B0(n16501), .Y(n15773) );
  AOI22XL U19550 ( .A0(B6_q[51]), .A1(n15958), .B0(B7_q[51]), .B1(n5930), .Y(
        n15774) );
  OAI211XL U19551 ( .A0(n5813), .A1(n15775), .B0(n15581), .C0(n15580), .Y(
        n15582) );
  AOI21XL U19552 ( .A0(B4_q[51]), .A1(n15687), .B0(n16501), .Y(n15580) );
  AOI22XL U19553 ( .A0(B6_q[51]), .A1(n16293), .B0(B7_q[51]), .B1(n16325), .Y(
        n15581) );
  OAI211XL U19554 ( .A0(n5806), .A1(n15775), .B0(n15390), .C0(n15389), .Y(
        n15391) );
  AOI21XL U19555 ( .A0(B4_q[51]), .A1(n5933), .B0(n16461), .Y(n15389) );
  AOI22XL U19556 ( .A0(B6_q[51]), .A1(n16143), .B0(B7_q[51]), .B1(n16128), .Y(
        n15390) );
  OAI211XL U19557 ( .A0(n5799), .A1(n15775), .B0(n15224), .C0(n15223), .Y(
        n15225) );
  AOI21XL U19558 ( .A0(B7_q[51]), .A1(n7127), .B0(n5924), .Y(n15223) );
  AOI22XL U19559 ( .A0(B4_q[51]), .A1(n7126), .B0(B6_q[51]), .B1(n16570), .Y(
        n15224) );
  NAND4XL U19560 ( .A(n15961), .B(n15960), .C(n5909), .D(n15959), .Y(n15962)
         );
  NAND2XL U19561 ( .A(B6_q[5]), .B(n15958), .Y(n15961) );
  NAND2XL U19562 ( .A(B5_q[5]), .B(n15963), .Y(n15960) );
  NAND4XL U19563 ( .A(n15560), .B(n15559), .C(n5909), .D(n15558), .Y(n15561)
         );
  NAND2XL U19564 ( .A(B7_q[5]), .B(n16158), .Y(n15560) );
  NAND2XL U19565 ( .A(B5_q[5]), .B(n16165), .Y(n15559) );
  NAND4XL U19566 ( .A(n15956), .B(n15955), .C(n5909), .D(n15954), .Y(n15957)
         );
  NAND2XL U19567 ( .A(B6_q[6]), .B(n15958), .Y(n15956) );
  NAND2XL U19568 ( .A(B5_q[6]), .B(n15963), .Y(n15955) );
  NAND4XL U19569 ( .A(n15750), .B(n15749), .C(n5909), .D(n15748), .Y(n15751)
         );
  NAND2XL U19570 ( .A(B6_q[6]), .B(n16293), .Y(n15750) );
  NAND2XL U19571 ( .A(B5_q[6]), .B(n15747), .Y(n15749) );
  NAND4XL U19572 ( .A(n15555), .B(n15554), .C(n5909), .D(n15553), .Y(n15556)
         );
  NAND2XL U19573 ( .A(B7_q[6]), .B(n16158), .Y(n15555) );
  NAND2XL U19574 ( .A(B5_q[6]), .B(n16165), .Y(n15554) );
  OAI211XL U19575 ( .A0(n15967), .A1(n15952), .B0(n15951), .C0(n15950), .Y(
        n15953) );
  AOI21XL U19576 ( .A0(B4_q[7]), .A1(n5925), .B0(n5924), .Y(n15950) );
  AOI22XL U19577 ( .A0(B6_q[7]), .A1(n15958), .B0(B5_q[7]), .B1(n15963), .Y(
        n15951) );
  OAI211XL U19578 ( .A0(n5813), .A1(n15745), .B0(n15744), .C0(n15743), .Y(
        n15746) );
  AOI21XL U19579 ( .A0(B4_q[7]), .A1(n15687), .B0(n16470), .Y(n15743) );
  AOI22XL U19580 ( .A0(B7_q[7]), .A1(n16325), .B0(B6_q[7]), .B1(n16354), .Y(
        n15744) );
  OAI211XL U19581 ( .A0(n5841), .A1(n15952), .B0(n15551), .C0(n15550), .Y(
        n15552) );
  AOI21XL U19582 ( .A0(B4_q[7]), .A1(n5933), .B0(n5924), .Y(n15550) );
  AOI22XL U19583 ( .A0(B6_q[7]), .A1(n16143), .B0(B5_q[7]), .B1(n16165), .Y(
        n15551) );
  OAI211XL U19584 ( .A0(n15948), .A1(n15947), .B0(n15946), .C0(n15945), .Y(
        n15949) );
  AOI21XL U19585 ( .A0(B4_q[8]), .A1(n5925), .B0(n5924), .Y(n15945) );
  AOI22XL U19586 ( .A0(B7_q[8]), .A1(n15982), .B0(B5_q[8]), .B1(n15963), .Y(
        n15946) );
  OAI211XL U19587 ( .A0(n5813), .A1(n15741), .B0(n15740), .C0(n15739), .Y(
        n15742) );
  AOI21XL U19588 ( .A0(B4_q[8]), .A1(n16277), .B0(n5924), .Y(n15739) );
  AOI22XL U19589 ( .A0(B6_q[8]), .A1(n16293), .B0(B7_q[8]), .B1(n16325), .Y(
        n15740) );
  OAI211XL U19590 ( .A0(n15495), .A1(n15947), .B0(n15548), .C0(n15547), .Y(
        n15549) );
  AOI21XL U19591 ( .A0(B4_q[8]), .A1(n15557), .B0(n5924), .Y(n15547) );
  AOI22XL U19592 ( .A0(B7_q[8]), .A1(n16158), .B0(B5_q[8]), .B1(n16165), .Y(
        n15548) );
  OAI211XL U19593 ( .A0(n15347), .A1(n5914), .B0(n15346), .C0(n15345), .Y(
        n15348) );
  AOI21XL U19594 ( .A0(B5_q[8]), .A1(n16559), .B0(n5924), .Y(n15345) );
  AOI22XL U19595 ( .A0(B7_q[8]), .A1(n7127), .B0(B6_q[8]), .B1(n16570), .Y(
        n15346) );
  NAND4XL U19596 ( .A(n15943), .B(n15942), .C(n5909), .D(n15941), .Y(n15944)
         );
  NAND2XL U19597 ( .A(B5_q[9]), .B(n15963), .Y(n15943) );
  NAND2XL U19598 ( .A(B7_q[9]), .B(n15982), .Y(n15942) );
  NAND4XL U19599 ( .A(n15737), .B(n15736), .C(n5915), .D(n15735), .Y(n15738)
         );
  NAND2XL U19600 ( .A(B6_q[9]), .B(n16293), .Y(n15737) );
  NAND2XL U19601 ( .A(B5_q[9]), .B(n15747), .Y(n15736) );
  NAND4XL U19602 ( .A(n15545), .B(n15544), .C(n5909), .D(n15543), .Y(n15546)
         );
  NAND2XL U19603 ( .A(B5_q[9]), .B(n5931), .Y(n15545) );
  NAND2XL U19604 ( .A(B7_q[9]), .B(n16158), .Y(n15544) );
  NAND4XL U19605 ( .A(n15343), .B(n15342), .C(n5915), .D(n15341), .Y(n15344)
         );
  NAND2XL U19606 ( .A(B4_q[9]), .B(n7126), .Y(n15343) );
  NAND2XL U19607 ( .A(B5_q[9]), .B(n16559), .Y(n15342) );
  MXI2XL U19608 ( .A(Q6[41]), .B(n21117), .S0(n24128), .Y(n3844) );
  XNOR2XL U19609 ( .A(n21168), .B(n21116), .Y(n21117) );
  NAND2XL U19610 ( .A(n21167), .B(n21220), .Y(n21116) );
  MXI2XL U19611 ( .A(Q6[42]), .B(n21174), .S0(n23239), .Y(n3845) );
  XOR2XL U19612 ( .A(n21173), .B(n21172), .Y(n21174) );
  NAND2XL U19613 ( .A(n21171), .B(n21219), .Y(n21172) );
  AOI21XL U19614 ( .A0(n21168), .A1(n21167), .B0(n21166), .Y(n21173) );
  MXI2XL U19615 ( .A(Q6[43]), .B(n21235), .S0(n23239), .Y(n3846) );
  XNOR2XL U19616 ( .A(n21384), .B(n21234), .Y(n21235) );
  NAND2XL U19617 ( .A(n21231), .B(n21297), .Y(n21234) );
  MXI2XL U19618 ( .A(Q6[44]), .B(n21303), .S0(n24128), .Y(n3847) );
  XOR2XL U19619 ( .A(n21302), .B(n21301), .Y(n21303) );
  NAND2XL U19620 ( .A(n21298), .B(n21326), .Y(n21301) );
  AOI21XL U19621 ( .A0(n21384), .A1(n21231), .B0(n21328), .Y(n21302) );
  MXI2XL U19622 ( .A(Q6[45]), .B(n21336), .S0(n23239), .Y(n3848) );
  XOR2XL U19623 ( .A(n21335), .B(n21334), .Y(n21336) );
  NAND2XL U19624 ( .A(n21333), .B(n21381), .Y(n21334) );
  AOI21XL U19625 ( .A0(n21384), .A1(n21330), .B0(n21329), .Y(n21335) );
  MXI2XL U19626 ( .A(Q6[46]), .B(n21390), .S0(n23239), .Y(n3849) );
  NAND2XL U19627 ( .A(n21385), .B(n21442), .Y(n21388) );
  AOI21XL U19628 ( .A0(n21384), .A1(n21441), .B0(n21444), .Y(n21389) );
  MXI2XL U19629 ( .A(Q6[47]), .B(n21452), .S0(n24128), .Y(n3850) );
  XNOR2XL U19630 ( .A(n21512), .B(n21451), .Y(n21452) );
  NAND2XL U19631 ( .A(n21448), .B(n21510), .Y(n21451) );
  MXI2XL U19632 ( .A(Q6[48]), .B(n21517), .S0(n23239), .Y(n3851) );
  XOR2XL U19633 ( .A(n21562), .B(n21516), .Y(n21517) );
  NAND2XL U19634 ( .A(n21515), .B(n21560), .Y(n21516) );
  INVXL U19635 ( .A(n21561), .Y(n21515) );
  MXI2XL U19636 ( .A(Q6[49]), .B(n21567), .S0(n24128), .Y(n3852) );
  XNOR2XL U19637 ( .A(n21606), .B(n21566), .Y(n21567) );
  NAND2XL U19638 ( .A(n21563), .B(n21604), .Y(n21566) );
  MXI2XL U19639 ( .A(Q6[50]), .B(n21611), .S0(n24128), .Y(n3853) );
  XOR2XL U19640 ( .A(n21632), .B(n21610), .Y(n21611) );
  NAND2XL U19641 ( .A(n21609), .B(n21630), .Y(n21610) );
  INVXL U19642 ( .A(n21631), .Y(n21609) );
  MXI2XL U19643 ( .A(Q6[51]), .B(n21637), .S0(n23239), .Y(n3854) );
  XNOR2XL U19644 ( .A(n21670), .B(n21636), .Y(n21637) );
  NAND2XL U19645 ( .A(n21633), .B(n21668), .Y(n21636) );
  XOR2XL U19646 ( .A(n21711), .B(n21674), .Y(n21675) );
  NAND2XL U19647 ( .A(n21673), .B(n21709), .Y(n21674) );
  INVXL U19648 ( .A(n21710), .Y(n21673) );
  XOR2XL U19649 ( .A(n28913), .B(U1_pipe3[27]), .Y(n21714) );
  MXI2XL U19650 ( .A(Q6[0]), .B(n16939), .S0(n23239), .Y(n3857) );
  XOR2XL U19651 ( .A(n17758), .B(n16938), .Y(n16939) );
  NAND2XL U19652 ( .A(n16937), .B(n17799), .Y(n16938) );
  INVXL U19653 ( .A(n17797), .Y(n16937) );
  MXI2XL U19654 ( .A(Q6[1]), .B(n17764), .S0(n23239), .Y(n3858) );
  XNOR2XL U19655 ( .A(n17763), .B(n17762), .Y(n17764) );
  NAND2XL U19656 ( .A(n17761), .B(n17798), .Y(n17762) );
  MXI2XL U19657 ( .A(Q6[2]), .B(n17807), .S0(n23239), .Y(n3859) );
  XNOR2XL U19658 ( .A(n17927), .B(n17806), .Y(n17807) );
  NAND2XL U19659 ( .A(n17851), .B(n17925), .Y(n17806) );
  MXI2XL U19660 ( .A(Q6[3]), .B(n17857), .S0(n23239), .Y(n3860) );
  XOR2XL U19661 ( .A(n17856), .B(n17855), .Y(n17857) );
  NAND2XL U19662 ( .A(n17854), .B(n17924), .Y(n17855) );
  AOI21XL U19663 ( .A0(n17927), .A1(n17851), .B0(n17850), .Y(n17856) );
  MXI2XL U19664 ( .A(Q6[4]), .B(n17932), .S0(n24128), .Y(n3861) );
  XOR2XL U19665 ( .A(n17945), .B(n17931), .Y(n17932) );
  NAND2XL U19666 ( .A(n17930), .B(n17988), .Y(n17931) );
  INVXL U19667 ( .A(n17985), .Y(n17930) );
  MXI2XL U19668 ( .A(Q6[5]), .B(n17951), .S0(n24128), .Y(n3862) );
  XNOR2XL U19669 ( .A(n17950), .B(n17949), .Y(n17951) );
  NAND2XL U19670 ( .A(n17948), .B(n17987), .Y(n17949) );
  MXI2XL U19671 ( .A(Q6[6]), .B(n18000), .S0(n23239), .Y(n3863) );
  XOR2XL U19672 ( .A(n18239), .B(n17999), .Y(n18000) );
  NAND2XL U19673 ( .A(n17998), .B(n18102), .Y(n17999) );
  INVXL U19674 ( .A(n18100), .Y(n17998) );
  MXI2XL U19675 ( .A(Q6[7]), .B(n18091), .S0(U1_valid[1]), .Y(n3864) );
  MXI2XL U19676 ( .A(Q6[8]), .B(n18109), .S0(U1_valid[1]), .Y(n3865) );
  XNOR2XL U19677 ( .A(n18150), .B(n18108), .Y(n18109) );
  NAND2XL U19678 ( .A(n18149), .B(n18234), .Y(n18108) );
  MXI2XL U19679 ( .A(Q6[9]), .B(n18156), .S0(U1_valid[1]), .Y(n3866) );
  XOR2XL U19680 ( .A(n18155), .B(n18154), .Y(n18156) );
  NAND2XL U19681 ( .A(n18153), .B(n18233), .Y(n18154) );
  AOI21XL U19682 ( .A0(n18150), .A1(n18149), .B0(n18148), .Y(n18155) );
  MXI2XL U19683 ( .A(Q6[10]), .B(n18243), .S0(n18351), .Y(n3867) );
  XOR2XL U19684 ( .A(n18325), .B(n18242), .Y(n18243) );
  NAND2XL U19685 ( .A(n18273), .B(n18321), .Y(n18242) );
  MXI2XL U19686 ( .A(Q6[11]), .B(n18280), .S0(n18351), .Y(n3868) );
  XOR2XL U19687 ( .A(n18279), .B(n18278), .Y(n18280) );
  NAND2XL U19688 ( .A(n18277), .B(n18320), .Y(n18278) );
  MXI2XL U19689 ( .A(Q6[12]), .B(n18329), .S0(n18351), .Y(n3869) );
  XNOR2XL U19690 ( .A(n18397), .B(n18328), .Y(n18329) );
  NAND2XL U19691 ( .A(n18396), .B(n18428), .Y(n18328) );
  MXI2XL U19692 ( .A(Q6[13]), .B(n18403), .S0(n24128), .Y(n3870) );
  XOR2XL U19693 ( .A(n18402), .B(n18401), .Y(n18403) );
  NAND2XL U19694 ( .A(n18400), .B(n18427), .Y(n18401) );
  AOI21XL U19695 ( .A0(n18397), .A1(n18396), .B0(n18395), .Y(n18402) );
  MXI2XL U19696 ( .A(Q6[14]), .B(n18442), .S0(n24128), .Y(n3871) );
  XNOR2XL U19697 ( .A(n18693), .B(n18441), .Y(n18442) );
  NAND2XL U19698 ( .A(n18521), .B(n18583), .Y(n18441) );
  MXI2XL U19699 ( .A(Q6[15]), .B(n18527), .S0(n24128), .Y(n3872) );
  XOR2XL U19700 ( .A(n18526), .B(n18525), .Y(n18527) );
  NAND2XL U19701 ( .A(n18524), .B(n18582), .Y(n18525) );
  AOI21XL U19702 ( .A0(n18693), .A1(n18521), .B0(n18520), .Y(n18526) );
  MXI2XL U19703 ( .A(Q6[16]), .B(n18590), .S0(n18739), .Y(n3873) );
  XOR2XL U19704 ( .A(n18589), .B(n18588), .Y(n18590) );
  NAND2XL U19705 ( .A(n18585), .B(n18614), .Y(n18588) );
  AOI21XL U19706 ( .A0(n18693), .A1(n18613), .B0(n18616), .Y(n18589) );
  MXI2XL U19707 ( .A(Q6[17]), .B(n18624), .S0(n18739), .Y(n3874) );
  XOR2XL U19708 ( .A(n18623), .B(n18622), .Y(n18624) );
  NAND2XL U19709 ( .A(n18621), .B(n18690), .Y(n18622) );
  AOI21XL U19710 ( .A0(n18693), .A1(n18618), .B0(n18617), .Y(n18623) );
  MXI2XL U19711 ( .A(Q6[18]), .B(n18699), .S0(n18739), .Y(n3875) );
  XOR2XL U19712 ( .A(n18698), .B(n18697), .Y(n18699) );
  NAND2XL U19713 ( .A(n18694), .B(n18754), .Y(n18697) );
  AOI21XL U19714 ( .A0(n18693), .A1(n18753), .B0(n18756), .Y(n18698) );
  MXI2XL U19715 ( .A(Q6[19]), .B(n18764), .S0(n18893), .Y(n3876) );
  XNOR2XL U19716 ( .A(n18784), .B(n18763), .Y(n18764) );
  NAND2XL U19717 ( .A(n18760), .B(n18782), .Y(n18763) );
  MXI2XL U19718 ( .A(Q6[20]), .B(n18789), .S0(n18893), .Y(n3877) );
  XOR2XL U19719 ( .A(n18850), .B(n18788), .Y(n18789) );
  NAND2XL U19720 ( .A(n18787), .B(n18848), .Y(n18788) );
  INVXL U19721 ( .A(n18849), .Y(n18787) );
  MXI2XL U19722 ( .A(Q6[21]), .B(n18855), .S0(n18893), .Y(n3878) );
  XNOR2XL U19723 ( .A(n18897), .B(n18854), .Y(n18855) );
  NAND2XL U19724 ( .A(n18851), .B(n18895), .Y(n18854) );
  MXI2XL U19725 ( .A(Q6[22]), .B(n18902), .S0(U1_valid[1]), .Y(n3879) );
  NAND2XL U19726 ( .A(n18900), .B(n18935), .Y(n18901) );
  INVXL U19727 ( .A(n18936), .Y(n18900) );
  MXI2XL U19728 ( .A(Q6[23]), .B(n18942), .S0(U1_valid[1]), .Y(n3880) );
  XNOR2XL U19729 ( .A(n18973), .B(n18941), .Y(n18942) );
  NAND2XL U19730 ( .A(n18938), .B(n18971), .Y(n18941) );
  MXI2XL U19731 ( .A(Q6[24]), .B(n18978), .S0(U1_valid[1]), .Y(n3881) );
  XOR2XL U19732 ( .A(n18997), .B(n18977), .Y(n18978) );
  NAND2XL U19733 ( .A(n18976), .B(n18995), .Y(n18977) );
  INVXL U19734 ( .A(n18996), .Y(n18976) );
  XOR2XL U19735 ( .A(n28696), .B(n28992), .Y(n19000) );
  MXI2XL U19736 ( .A(Q7[28]), .B(n20187), .S0(n23239), .Y(n3883) );
  XOR2XL U19737 ( .A(n20186), .B(n20491), .Y(n20187) );
  NAND2XL U19738 ( .A(n20182), .B(n20489), .Y(n20186) );
  INVXL U19739 ( .A(n20490), .Y(n20182) );
  MXI2XL U19740 ( .A(Q7[29]), .B(n20496), .S0(n23239), .Y(n3884) );
  XOR2XL U19741 ( .A(n20533), .B(n20495), .Y(n20496) );
  NAND2XL U19742 ( .A(n20494), .B(n20581), .Y(n20495) );
  INVXL U19743 ( .A(n20579), .Y(n20494) );
  MXI2XL U19744 ( .A(Q7[30]), .B(n20539), .S0(n24128), .Y(n3885) );
  XNOR2XL U19745 ( .A(n20538), .B(n20537), .Y(n20539) );
  NAND2XL U19746 ( .A(n20536), .B(n20580), .Y(n20537) );
  MXI2XL U19747 ( .A(Q7[31]), .B(n20589), .S0(n23239), .Y(n3886) );
  XNOR2XL U19748 ( .A(n20678), .B(n20588), .Y(n20589) );
  NAND2XL U19749 ( .A(n20630), .B(n20676), .Y(n20588) );
  MXI2XL U19750 ( .A(Q7[32]), .B(n20636), .S0(n24128), .Y(n3887) );
  XOR2XL U19751 ( .A(n20635), .B(n20634), .Y(n20636) );
  NAND2XL U19752 ( .A(n20633), .B(n20675), .Y(n20634) );
  AOI21XL U19753 ( .A0(n20678), .A1(n20630), .B0(n20629), .Y(n20635) );
  MXI2XL U19754 ( .A(Q7[33]), .B(n20683), .S0(n23239), .Y(n3888) );
  XOR2XL U19755 ( .A(n20726), .B(n20682), .Y(n20683) );
  NAND2XL U19756 ( .A(n20681), .B(n20783), .Y(n20682) );
  INVXL U19757 ( .A(n20780), .Y(n20681) );
  MXI2XL U19758 ( .A(Q7[34]), .B(n20732), .S0(n24128), .Y(n3889) );
  XNOR2XL U19759 ( .A(n20731), .B(n20730), .Y(n20732) );
  NAND2XL U19760 ( .A(n20729), .B(n20782), .Y(n20730) );
  MXI2XL U19761 ( .A(Q7[35]), .B(n20795), .S0(n24128), .Y(n3890) );
  XOR2XL U19762 ( .A(n20973), .B(n20794), .Y(n20795) );
  NAND2XL U19763 ( .A(n20793), .B(n20881), .Y(n20794) );
  INVXL U19764 ( .A(n20879), .Y(n20793) );
  MXI2XL U19765 ( .A(Q7[36]), .B(n20841), .S0(n24128), .Y(n3891) );
  XNOR2XL U19766 ( .A(n20840), .B(n20839), .Y(n20841) );
  NAND2XL U19767 ( .A(n20838), .B(n20880), .Y(n20839) );
  MXI2XL U19768 ( .A(Q7[37]), .B(n20888), .S0(n23239), .Y(n3892) );
  XNOR2XL U19769 ( .A(n20934), .B(n20887), .Y(n20888) );
  NAND2XL U19770 ( .A(n20933), .B(n20968), .Y(n20887) );
  MXI2XL U19771 ( .A(Q7[38]), .B(n20940), .S0(n24128), .Y(n3893) );
  XOR2XL U19772 ( .A(n20939), .B(n20938), .Y(n20940) );
  NAND2XL U19773 ( .A(n20937), .B(n20967), .Y(n20938) );
  AOI21XL U19774 ( .A0(n20934), .A1(n20933), .B0(n20932), .Y(n20939) );
  MXI2XL U19775 ( .A(Q7[39]), .B(n20977), .S0(n24128), .Y(n3894) );
  NAND2XL U19776 ( .A(n21026), .B(n21078), .Y(n20976) );
  MXI2XL U19777 ( .A(Q7[40]), .B(n21033), .S0(n23239), .Y(n3895) );
  XOR2XL U19778 ( .A(n21032), .B(n21031), .Y(n21033) );
  NAND2XL U19779 ( .A(n21030), .B(n21077), .Y(n21031) );
  AOI21XL U19780 ( .A0(n21027), .A1(n21026), .B0(n21025), .Y(n21032) );
  MXI2XL U19781 ( .A(Q7[41]), .B(n21086), .S0(n24128), .Y(n3896) );
  XNOR2XL U19782 ( .A(n21131), .B(n21085), .Y(n21086) );
  NAND2XL U19783 ( .A(n21130), .B(n21200), .Y(n21085) );
  MXI2XL U19784 ( .A(Q7[42]), .B(n21137), .S0(n23239), .Y(n3897) );
  XOR2XL U19785 ( .A(n21136), .B(n21135), .Y(n21137) );
  NAND2XL U19786 ( .A(n21134), .B(n21199), .Y(n21135) );
  AOI21XL U19787 ( .A0(n21131), .A1(n21130), .B0(n21129), .Y(n21136) );
  MXI2XL U19788 ( .A(Q7[43]), .B(n21215), .S0(n24128), .Y(n3898) );
  XNOR2XL U19789 ( .A(n21373), .B(n21214), .Y(n21215) );
  NAND2XL U19790 ( .A(n21211), .B(n21273), .Y(n21214) );
  MXI2XL U19791 ( .A(Q7[44]), .B(n21279), .S0(n23239), .Y(n3899) );
  XOR2XL U19792 ( .A(n21278), .B(n21277), .Y(n21279) );
  NAND2XL U19793 ( .A(n21274), .B(n21315), .Y(n21277) );
  AOI21XL U19794 ( .A0(n21373), .A1(n21211), .B0(n21317), .Y(n21278) );
  MXI2XL U19795 ( .A(Q7[45]), .B(n21325), .S0(n24128), .Y(n3900) );
  XOR2XL U19796 ( .A(n21324), .B(n21323), .Y(n21325) );
  NAND2XL U19797 ( .A(n21322), .B(n21370), .Y(n21323) );
  AOI21XL U19798 ( .A0(n21373), .A1(n21319), .B0(n21318), .Y(n21324) );
  MXI2XL U19799 ( .A(Q7[46]), .B(n21379), .S0(n24128), .Y(n3901) );
  XOR2XL U19800 ( .A(n21378), .B(n21377), .Y(n21379) );
  NAND2XL U19801 ( .A(n21374), .B(n21430), .Y(n21377) );
  AOI21XL U19802 ( .A0(n21373), .A1(n21429), .B0(n21432), .Y(n21378) );
  MXI2XL U19803 ( .A(Q7[47]), .B(n21440), .S0(n23239), .Y(n3902) );
  XNOR2XL U19804 ( .A(n21488), .B(n21439), .Y(n21440) );
  NAND2XL U19805 ( .A(n21436), .B(n21486), .Y(n21439) );
  MXI2XL U19806 ( .A(Q7[48]), .B(n21493), .S0(n23239), .Y(n3903) );
  XOR2XL U19807 ( .A(n21538), .B(n21492), .Y(n21493) );
  NAND2XL U19808 ( .A(n21491), .B(n21536), .Y(n21492) );
  INVXL U19809 ( .A(n21537), .Y(n21491) );
  MXI2XL U19810 ( .A(Q7[49]), .B(n21543), .S0(n24128), .Y(n3904) );
  XNOR2XL U19811 ( .A(n21582), .B(n21542), .Y(n21543) );
  NAND2XL U19812 ( .A(n21539), .B(n21580), .Y(n21542) );
  MXI2XL U19813 ( .A(Q7[50]), .B(n21587), .S0(n23239), .Y(n3905) );
  XOR2XL U19814 ( .A(n21624), .B(n21586), .Y(n21587) );
  NAND2XL U19815 ( .A(n21585), .B(n21622), .Y(n21586) );
  INVXL U19816 ( .A(n21623), .Y(n21585) );
  MXI2XL U19817 ( .A(Q7[51]), .B(n21629), .S0(n24128), .Y(n3906) );
  XNOR2XL U19818 ( .A(n21662), .B(n21628), .Y(n21629) );
  NAND2XL U19819 ( .A(n21625), .B(n21660), .Y(n21628) );
  XOR2XL U19820 ( .A(n21704), .B(n21666), .Y(n21667) );
  NAND2XL U19821 ( .A(n21665), .B(n21702), .Y(n21666) );
  INVXL U19822 ( .A(n21703), .Y(n21665) );
  XOR2XL U19823 ( .A(n28918), .B(U1_pipe13[27]), .Y(n21707) );
  MXI2XL U19824 ( .A(Q7[0]), .B(n17453), .S0(n23239), .Y(n3909) );
  NAND2XL U19825 ( .A(n17448), .B(n17772), .Y(n17452) );
  INVXL U19826 ( .A(n17773), .Y(n17448) );
  MXI2XL U19827 ( .A(Q7[1]), .B(n17779), .S0(n24128), .Y(n3910) );
  XOR2XL U19828 ( .A(n17819), .B(n17778), .Y(n17779) );
  NAND2XL U19829 ( .A(n17777), .B(n17868), .Y(n17778) );
  INVXL U19830 ( .A(n17866), .Y(n17777) );
  MXI2XL U19831 ( .A(Q7[2]), .B(n17825), .S0(n24128), .Y(n3911) );
  XNOR2XL U19832 ( .A(n17824), .B(n17823), .Y(n17825) );
  NAND2XL U19833 ( .A(n17822), .B(n17867), .Y(n17823) );
  MXI2XL U19834 ( .A(Q7[3]), .B(n17876), .S0(n23239), .Y(n3912) );
  XNOR2XL U19835 ( .A(n17963), .B(n17875), .Y(n17876) );
  NAND2XL U19836 ( .A(n17916), .B(n17961), .Y(n17875) );
  MXI2XL U19837 ( .A(Q7[4]), .B(n17922), .S0(n23239), .Y(n3913) );
  XOR2XL U19838 ( .A(n17921), .B(n17920), .Y(n17922) );
  NAND2XL U19839 ( .A(n17919), .B(n17960), .Y(n17920) );
  AOI21XL U19840 ( .A0(n17963), .A1(n17916), .B0(n17915), .Y(n17921) );
  MXI2XL U19841 ( .A(Q7[5]), .B(n17968), .S0(n24128), .Y(n3914) );
  XOR2XL U19842 ( .A(n18017), .B(n17967), .Y(n17968) );
  NAND2XL U19843 ( .A(n17966), .B(n18073), .Y(n17967) );
  INVXL U19844 ( .A(n18070), .Y(n17966) );
  MXI2XL U19845 ( .A(Q7[6]), .B(n18023), .S0(U1_valid[1]), .Y(n3915) );
  XNOR2XL U19846 ( .A(n18022), .B(n18021), .Y(n18023) );
  NAND2XL U19847 ( .A(n18020), .B(n18072), .Y(n18021) );
  MXI2XL U19848 ( .A(Q7[7]), .B(n18085), .S0(U1_valid[1]), .Y(n3916) );
  XOR2XL U19849 ( .A(n18267), .B(n18084), .Y(n18085) );
  NAND2XL U19850 ( .A(n18083), .B(n18168), .Y(n18084) );
  INVXL U19851 ( .A(n18166), .Y(n18083) );
  MXI2XL U19852 ( .A(Q7[8]), .B(n18125), .S0(U1_valid[1]), .Y(n3917) );
  XNOR2XL U19853 ( .A(n18124), .B(n18123), .Y(n18125) );
  NAND2XL U19854 ( .A(n18122), .B(n18167), .Y(n18123) );
  MXI2XL U19855 ( .A(Q7[9]), .B(n18175), .S0(U1_valid[1]), .Y(n3918) );
  XNOR2XL U19856 ( .A(n18224), .B(n18174), .Y(n18175) );
  NAND2XL U19857 ( .A(n18223), .B(n18262), .Y(n18174) );
  MXI2XL U19858 ( .A(Q7[10]), .B(n18230), .S0(n18351), .Y(n3919) );
  XOR2XL U19859 ( .A(n18229), .B(n18228), .Y(n18230) );
  NAND2XL U19860 ( .A(n18227), .B(n18261), .Y(n18228) );
  AOI21XL U19861 ( .A0(n18224), .A1(n18223), .B0(n18222), .Y(n18229) );
  MXI2XL U19862 ( .A(Q7[11]), .B(n18271), .S0(n18351), .Y(n3920) );
  XOR2XL U19863 ( .A(n18372), .B(n18270), .Y(n18271) );
  NAND2XL U19864 ( .A(n18311), .B(n18368), .Y(n18270) );
  MXI2XL U19865 ( .A(Q7[12]), .B(n18318), .S0(n18351), .Y(n3921) );
  XOR2XL U19866 ( .A(n18317), .B(n18316), .Y(n18318) );
  NAND2XL U19867 ( .A(n18315), .B(n18367), .Y(n18316) );
  AOI21XL U19868 ( .A0(n18312), .A1(n18311), .B0(n18310), .Y(n18317) );
  MXI2XL U19869 ( .A(Q7[13]), .B(n18376), .S0(n24128), .Y(n3922) );
  XNOR2XL U19870 ( .A(n18417), .B(n18375), .Y(n18376) );
  NAND2XL U19871 ( .A(n18416), .B(n18504), .Y(n18375) );
  MXI2XL U19872 ( .A(Q7[14]), .B(n18423), .S0(n23239), .Y(n3923) );
  XOR2XL U19873 ( .A(n18422), .B(n18421), .Y(n18423) );
  NAND2XL U19874 ( .A(n18420), .B(n18503), .Y(n18421) );
  AOI21XL U19875 ( .A0(n18417), .A1(n18416), .B0(n18415), .Y(n18422) );
  MXI2XL U19876 ( .A(Q7[15]), .B(n18519), .S0(n23239), .Y(n3924) );
  MXI2XL U19877 ( .A(Q7[16]), .B(n18560), .S0(n23239), .Y(n3925) );
  XOR2XL U19878 ( .A(n18559), .B(n18558), .Y(n18560) );
  NAND2XL U19879 ( .A(n18555), .B(n18602), .Y(n18558) );
  AOI21XL U19880 ( .A0(n18660), .A1(n18515), .B0(n18604), .Y(n18559) );
  MXI2XL U19881 ( .A(Q7[17]), .B(n18612), .S0(n18739), .Y(n3926) );
  XOR2XL U19882 ( .A(n18611), .B(n18610), .Y(n18612) );
  NAND2XL U19883 ( .A(n18609), .B(n18657), .Y(n18610) );
  AOI21XL U19884 ( .A0(n18660), .A1(n18606), .B0(n18605), .Y(n18611) );
  MXI2XL U19885 ( .A(Q7[18]), .B(n18666), .S0(n18739), .Y(n3927) );
  XOR2XL U19886 ( .A(n18665), .B(n18664), .Y(n18666) );
  NAND2XL U19887 ( .A(n18661), .B(n18717), .Y(n18664) );
  MXI2XL U19888 ( .A(Q7[19]), .B(n18727), .S0(n18739), .Y(n3928) );
  XNOR2XL U19889 ( .A(n18776), .B(n18726), .Y(n18727) );
  NAND2XL U19890 ( .A(n18723), .B(n18774), .Y(n18726) );
  MXI2XL U19891 ( .A(Q7[20]), .B(n18781), .S0(n18893), .Y(n3929) );
  XOR2XL U19892 ( .A(n18826), .B(n18780), .Y(n18781) );
  NAND2XL U19893 ( .A(n18779), .B(n18824), .Y(n18780) );
  INVXL U19894 ( .A(n18825), .Y(n18779) );
  MXI2XL U19895 ( .A(Q7[21]), .B(n18831), .S0(n18893), .Y(n3930) );
  XNOR2XL U19896 ( .A(n18872), .B(n18830), .Y(n18831) );
  NAND2XL U19897 ( .A(n18827), .B(n18870), .Y(n18830) );
  MXI2XL U19898 ( .A(Q7[22]), .B(n18877), .S0(n18893), .Y(n3931) );
  XOR2XL U19899 ( .A(n18913), .B(n18876), .Y(n18877) );
  NAND2XL U19900 ( .A(n18875), .B(n18911), .Y(n18876) );
  INVXL U19901 ( .A(n18912), .Y(n18875) );
  MXI2XL U19902 ( .A(Q7[23]), .B(n18918), .S0(U1_valid[1]), .Y(n3932) );
  XNOR2XL U19903 ( .A(n18949), .B(n18917), .Y(n18918) );
  NAND2XL U19904 ( .A(n18914), .B(n18947), .Y(n18917) );
  MXI2XL U19905 ( .A(Q7[24]), .B(n18954), .S0(U1_valid[1]), .Y(n3933) );
  XOR2XL U19906 ( .A(n18990), .B(n18953), .Y(n18954) );
  NAND2XL U19907 ( .A(n18952), .B(n18988), .Y(n18953) );
  INVXL U19908 ( .A(n18989), .Y(n18952) );
  MXI2XL U19909 ( .A(Q4[28]), .B(n19708), .S0(n23239), .Y(n3935) );
  XOR2XL U19910 ( .A(n20482), .B(n19707), .Y(n19708) );
  NAND2XL U19911 ( .A(n19706), .B(n20524), .Y(n19707) );
  INVXL U19912 ( .A(n20522), .Y(n19706) );
  MXI2XL U19913 ( .A(Q4[0]), .B(n17173), .S0(n23239), .Y(n3936) );
  XOR2XL U19914 ( .A(n17765), .B(n17172), .Y(n17173) );
  NAND2XL U19915 ( .A(n17171), .B(n17810), .Y(n17172) );
  INVXL U19916 ( .A(n17808), .Y(n17171) );
  MXI2XL U19917 ( .A(Q4[1]), .B(n17771), .S0(n23239), .Y(n3937) );
  XNOR2XL U19918 ( .A(n17770), .B(n17769), .Y(n17771) );
  NAND2XL U19919 ( .A(n17768), .B(n17809), .Y(n17769) );
  MXI2XL U19920 ( .A(Q4[2]), .B(n17818), .S0(n23239), .Y(n3938) );
  XNOR2XL U19921 ( .A(n17909), .B(n17817), .Y(n17818) );
  NAND2XL U19922 ( .A(n17859), .B(n17907), .Y(n17817) );
  MXI2XL U19923 ( .A(Q4[3]), .B(n17865), .S0(n23239), .Y(n3939) );
  AOI21XL U19924 ( .A0(n17909), .A1(n17859), .B0(n17858), .Y(n17864) );
  MXI2XL U19925 ( .A(Q4[4]), .B(n17914), .S0(n24128), .Y(n3940) );
  XOR2XL U19926 ( .A(n17952), .B(n17913), .Y(n17914) );
  NAND2XL U19927 ( .A(n17912), .B(n18004), .Y(n17913) );
  INVXL U19928 ( .A(n18001), .Y(n17912) );
  MXI2XL U19929 ( .A(Q4[5]), .B(n17958), .S0(n24128), .Y(n3941) );
  XNOR2XL U19930 ( .A(n17957), .B(n17956), .Y(n17958) );
  NAND2XL U19931 ( .A(n17955), .B(n18003), .Y(n17956) );
  MXI2XL U19932 ( .A(Q4[6]), .B(n18016), .S0(n24128), .Y(n3942) );
  XOR2XL U19933 ( .A(n18217), .B(n18015), .Y(n18016) );
  NAND2XL U19934 ( .A(n18014), .B(n18112), .Y(n18015) );
  INVXL U19935 ( .A(n18110), .Y(n18014) );
  MXI2XL U19936 ( .A(Q4[7]), .B(n18069), .S0(U1_valid[1]), .Y(n3943) );
  XNOR2XL U19937 ( .A(n18068), .B(n18067), .Y(n18069) );
  NAND2XL U19938 ( .A(n18066), .B(n18111), .Y(n18067) );
  MXI2XL U19939 ( .A(Q4[8]), .B(n18119), .S0(U1_valid[1]), .Y(n3944) );
  XNOR2XL U19940 ( .A(n18159), .B(n18118), .Y(n18119) );
  NAND2XL U19941 ( .A(n18158), .B(n18212), .Y(n18118) );
  MXI2XL U19942 ( .A(Q4[9]), .B(n18165), .S0(U1_valid[1]), .Y(n3945) );
  XOR2XL U19943 ( .A(n18164), .B(n18163), .Y(n18165) );
  NAND2XL U19944 ( .A(n18162), .B(n18211), .Y(n18163) );
  AOI21XL U19945 ( .A0(n18159), .A1(n18158), .B0(n18157), .Y(n18164) );
  MXI2XL U19946 ( .A(Q4[10]), .B(n18221), .S0(n18351), .Y(n3946) );
  XOR2XL U19947 ( .A(n18336), .B(n18220), .Y(n18221) );
  NAND2XL U19948 ( .A(n18282), .B(n18332), .Y(n18220) );
  MXI2XL U19949 ( .A(Q4[11]), .B(n18289), .S0(n18351), .Y(n3947) );
  XOR2XL U19950 ( .A(n18288), .B(n18287), .Y(n18289) );
  NAND2XL U19951 ( .A(n18286), .B(n18331), .Y(n18287) );
  AOI21XL U19952 ( .A0(n18283), .A1(n18282), .B0(n18281), .Y(n18288) );
  MXI2XL U19953 ( .A(Q4[12]), .B(n18340), .S0(n18351), .Y(n3948) );
  XNOR2XL U19954 ( .A(n18388), .B(n18339), .Y(n18340) );
  NAND2XL U19955 ( .A(n18387), .B(n18447), .Y(n18339) );
  MXI2XL U19956 ( .A(Q4[13]), .B(n18394), .S0(n23239), .Y(n3949) );
  XOR2XL U19957 ( .A(n18393), .B(n18392), .Y(n18394) );
  NAND2XL U19958 ( .A(n18391), .B(n18446), .Y(n18392) );
  MXI2XL U19959 ( .A(Q4[14]), .B(n18461), .S0(n23239), .Y(n3950) );
  XNOR2XL U19960 ( .A(n18682), .B(n18460), .Y(n18461) );
  NAND2XL U19961 ( .A(n18529), .B(n18573), .Y(n18460) );
  MXI2XL U19962 ( .A(Q4[15]), .B(n18535), .S0(n23239), .Y(n3951) );
  XOR2XL U19963 ( .A(n18534), .B(n18533), .Y(n18535) );
  NAND2XL U19964 ( .A(n18532), .B(n18572), .Y(n18533) );
  AOI21XL U19965 ( .A0(n18682), .A1(n18529), .B0(n18528), .Y(n18534) );
  MXI2XL U19966 ( .A(Q4[16]), .B(n18580), .S0(n18739), .Y(n3952) );
  XOR2XL U19967 ( .A(n18579), .B(n18578), .Y(n18580) );
  NAND2XL U19968 ( .A(n18575), .B(n18626), .Y(n18578) );
  AOI21XL U19969 ( .A0(n18682), .A1(n18625), .B0(n18628), .Y(n18579) );
  MXI2XL U19970 ( .A(Q4[17]), .B(n18636), .S0(n18739), .Y(n3953) );
  XOR2XL U19971 ( .A(n18635), .B(n18634), .Y(n18636) );
  NAND2XL U19972 ( .A(n18633), .B(n18679), .Y(n18634) );
  AOI21XL U19973 ( .A0(n18682), .A1(n18630), .B0(n18629), .Y(n18635) );
  MXI2XL U19974 ( .A(Q4[18]), .B(n18688), .S0(n18739), .Y(n3954) );
  NAND2XL U19975 ( .A(n18683), .B(n18742), .Y(n18686) );
  AOI21XL U19976 ( .A0(n18682), .A1(n18741), .B0(n18744), .Y(n18687) );
  MXI2XL U19977 ( .A(Q4[19]), .B(n18752), .S0(n18893), .Y(n3955) );
  XNOR2XL U19978 ( .A(n18792), .B(n18751), .Y(n18752) );
  NAND2XL U19979 ( .A(n18748), .B(n18790), .Y(n18751) );
  MXI2XL U19980 ( .A(Q4[20]), .B(n18797), .S0(n18893), .Y(n3956) );
  XOR2XL U19981 ( .A(n18842), .B(n18796), .Y(n18797) );
  NAND2XL U19982 ( .A(n18795), .B(n18840), .Y(n18796) );
  INVXL U19983 ( .A(n18841), .Y(n18795) );
  MXI2XL U19984 ( .A(Q4[21]), .B(n18847), .S0(n18893), .Y(n3957) );
  XNOR2XL U19985 ( .A(n18888), .B(n18846), .Y(n18847) );
  NAND2XL U19986 ( .A(n18843), .B(n18886), .Y(n18846) );
  MXI2XL U19987 ( .A(Q4[22]), .B(n18894), .S0(n18893), .Y(n3958) );
  XOR2XL U19988 ( .A(n18929), .B(n18892), .Y(n18894) );
  NAND2XL U19989 ( .A(n18891), .B(n18927), .Y(n18892) );
  INVXL U19990 ( .A(n18928), .Y(n18891) );
  MXI2XL U19991 ( .A(Q4[23]), .B(n18934), .S0(U1_valid[1]), .Y(n3959) );
  XNOR2XL U19992 ( .A(n18965), .B(n18933), .Y(n18934) );
  NAND2XL U19993 ( .A(n18930), .B(n18963), .Y(n18933) );
  MXI2XL U19994 ( .A(Q4[24]), .B(n18970), .S0(U1_valid[1]), .Y(n3960) );
  XOR2XL U19995 ( .A(n19004), .B(n18969), .Y(n18970) );
  NAND2XL U19996 ( .A(n18968), .B(n19002), .Y(n18969) );
  INVXL U19997 ( .A(n19003), .Y(n18968) );
  XOR2XL U19998 ( .A(n28694), .B(n28990), .Y(n19007) );
  MXI2XL U19999 ( .A(Q5[28]), .B(n20465), .S0(n23239), .Y(n3962) );
  XOR2XL U20000 ( .A(n20464), .B(n20499), .Y(n20465) );
  NAND2XL U20001 ( .A(n20460), .B(n20497), .Y(n20464) );
  INVXL U20002 ( .A(n20498), .Y(n20460) );
  MXI2XL U20003 ( .A(Q5[29]), .B(n20504), .S0(n23239), .Y(n3963) );
  XOR2XL U20004 ( .A(n20540), .B(n20503), .Y(n20504) );
  NAND2XL U20005 ( .A(n20502), .B(n20562), .Y(n20503) );
  INVXL U20006 ( .A(n20560), .Y(n20502) );
  MXI2XL U20007 ( .A(Q5[30]), .B(n20546), .S0(n23239), .Y(n3964) );
  XNOR2XL U20008 ( .A(n20545), .B(n20544), .Y(n20546) );
  NAND2XL U20009 ( .A(n20543), .B(n20561), .Y(n20544) );
  MXI2XL U20010 ( .A(Q5[31]), .B(n20570), .S0(n24128), .Y(n3965) );
  XNOR2XL U20011 ( .A(n20688), .B(n20569), .Y(n20570) );
  NAND2XL U20012 ( .A(n20638), .B(n20686), .Y(n20569) );
  MXI2XL U20013 ( .A(Q5[32]), .B(n20644), .S0(n23239), .Y(n3966) );
  XOR2XL U20014 ( .A(n20643), .B(n20642), .Y(n20644) );
  NAND2XL U20015 ( .A(n20641), .B(n20685), .Y(n20642) );
  AOI21XL U20016 ( .A0(n20688), .A1(n20638), .B0(n20637), .Y(n20643) );
  MXI2XL U20017 ( .A(Q5[33]), .B(n20693), .S0(n24128), .Y(n3967) );
  XOR2XL U20018 ( .A(n20703), .B(n20692), .Y(n20693) );
  NAND2XL U20019 ( .A(n20691), .B(n20761), .Y(n20692) );
  INVXL U20020 ( .A(n20758), .Y(n20691) );
  MXI2XL U20021 ( .A(Q5[34]), .B(n20709), .S0(n24128), .Y(n3968) );
  XNOR2XL U20022 ( .A(n20708), .B(n20707), .Y(n20709) );
  NAND2XL U20023 ( .A(n20706), .B(n20760), .Y(n20707) );
  MXI2XL U20024 ( .A(Q5[35]), .B(n20773), .S0(n24128), .Y(n3969) );
  INVXL U20025 ( .A(n20889), .Y(n20771) );
  MXI2XL U20026 ( .A(Q5[36]), .B(n20847), .S0(n23239), .Y(n3970) );
  XNOR2XL U20027 ( .A(n20846), .B(n20845), .Y(n20847) );
  NAND2XL U20028 ( .A(n20844), .B(n20890), .Y(n20845) );
  MXI2XL U20029 ( .A(Q5[37]), .B(n20898), .S0(n23239), .Y(n3971) );
  XNOR2XL U20030 ( .A(n20943), .B(n20897), .Y(n20898) );
  NAND2XL U20031 ( .A(n20942), .B(n20981), .Y(n20897) );
  MXI2XL U20032 ( .A(Q5[38]), .B(n20949), .S0(n23239), .Y(n3972) );
  XOR2XL U20033 ( .A(n20948), .B(n20947), .Y(n20949) );
  NAND2XL U20034 ( .A(n20946), .B(n20980), .Y(n20947) );
  AOI21XL U20035 ( .A0(n20943), .A1(n20942), .B0(n20941), .Y(n20948) );
  MXI2XL U20036 ( .A(Q5[39]), .B(n20990), .S0(n24128), .Y(n3973) );
  XOR2XL U20037 ( .A(n21093), .B(n20989), .Y(n20990) );
  NAND2XL U20038 ( .A(n21035), .B(n21089), .Y(n20989) );
  MXI2XL U20039 ( .A(Q5[40]), .B(n21042), .S0(n24128), .Y(n3974) );
  XOR2XL U20040 ( .A(n21041), .B(n21040), .Y(n21042) );
  NAND2XL U20041 ( .A(n21039), .B(n21088), .Y(n21040) );
  AOI21XL U20042 ( .A0(n21036), .A1(n21035), .B0(n21034), .Y(n21041) );
  MXI2XL U20043 ( .A(Q5[41]), .B(n21097), .S0(n23239), .Y(n3975) );
  XNOR2XL U20044 ( .A(n21140), .B(n21096), .Y(n21097) );
  NAND2XL U20045 ( .A(n21139), .B(n21248), .Y(n21096) );
  MXI2XL U20046 ( .A(Q5[42]), .B(n21146), .S0(n23239), .Y(n3976) );
  XOR2XL U20047 ( .A(n21145), .B(n21144), .Y(n21146) );
  NAND2XL U20048 ( .A(n21143), .B(n21247), .Y(n21144) );
  AOI21XL U20049 ( .A0(n21140), .A1(n21139), .B0(n21138), .Y(n21145) );
  MXI2XL U20050 ( .A(Q5[43]), .B(n21263), .S0(n24128), .Y(n3977) );
  XNOR2XL U20051 ( .A(n21406), .B(n21262), .Y(n21263) );
  NAND2XL U20052 ( .A(n21259), .B(n21280), .Y(n21262) );
  MXI2XL U20053 ( .A(Q5[44]), .B(n21286), .S0(n23239), .Y(n3978) );
  XOR2XL U20054 ( .A(n21285), .B(n21284), .Y(n21286) );
  NAND2XL U20055 ( .A(n21281), .B(n21349), .Y(n21284) );
  AOI21XL U20056 ( .A0(n21406), .A1(n21259), .B0(n21351), .Y(n21285) );
  MXI2XL U20057 ( .A(Q5[45]), .B(n21359), .S0(n24128), .Y(n3979) );
  XOR2XL U20058 ( .A(n21358), .B(n21357), .Y(n21359) );
  NAND2XL U20059 ( .A(n21356), .B(n21403), .Y(n21357) );
  AOI21XL U20060 ( .A0(n21406), .A1(n21353), .B0(n21352), .Y(n21358) );
  MXI2XL U20061 ( .A(Q5[46]), .B(n21412), .S0(n23239), .Y(n3980) );
  XOR2XL U20062 ( .A(n21411), .B(n21410), .Y(n21412) );
  NAND2XL U20063 ( .A(n21407), .B(n21466), .Y(n21410) );
  AOI21XL U20064 ( .A0(n21406), .A1(n21465), .B0(n21468), .Y(n21411) );
  MXI2XL U20065 ( .A(Q5[47]), .B(n21476), .S0(n24128), .Y(n3981) );
  XNOR2XL U20066 ( .A(n21496), .B(n21475), .Y(n21476) );
  NAND2XL U20067 ( .A(n21472), .B(n21494), .Y(n21475) );
  MXI2XL U20068 ( .A(Q5[48]), .B(n21501), .S0(n24128), .Y(n3982) );
  XOR2XL U20069 ( .A(n21546), .B(n21500), .Y(n21501) );
  NAND2XL U20070 ( .A(n21499), .B(n21544), .Y(n21500) );
  INVXL U20071 ( .A(n21545), .Y(n21499) );
  MXI2XL U20072 ( .A(Q5[49]), .B(n21551), .S0(n24128), .Y(n3983) );
  XNOR2XL U20073 ( .A(n21590), .B(n21550), .Y(n21551) );
  NAND2XL U20074 ( .A(n21547), .B(n21588), .Y(n21550) );
  MXI2XL U20075 ( .A(Q5[50]), .B(n21595), .S0(n23239), .Y(n3984) );
  NAND2XL U20076 ( .A(n21593), .B(n21646), .Y(n21594) );
  INVXL U20077 ( .A(n21647), .Y(n21593) );
  MXI2XL U20078 ( .A(Q5[51]), .B(n21653), .S0(n24128), .Y(n3985) );
  XNOR2XL U20079 ( .A(n21686), .B(n21652), .Y(n21653) );
  NAND2XL U20080 ( .A(n21649), .B(n21684), .Y(n21652) );
  XOR2XL U20081 ( .A(n21725), .B(n21690), .Y(n21691) );
  NAND2XL U20082 ( .A(n21689), .B(n21723), .Y(n21690) );
  INVXL U20083 ( .A(n21724), .Y(n21689) );
  XOR2XL U20084 ( .A(n28987), .B(U1_pipe9[27]), .Y(n21728) );
  MXI2XL U20085 ( .A(Q5[0]), .B(n17749), .S0(n23239), .Y(n3988) );
  XOR2XL U20086 ( .A(n17780), .B(n17748), .Y(n17749) );
  NAND2XL U20087 ( .A(n17747), .B(n17828), .Y(n17748) );
  INVXL U20088 ( .A(n17826), .Y(n17747) );
  MXI2XL U20089 ( .A(Q5[1]), .B(n17786), .S0(n24128), .Y(n3989) );
  XNOR2XL U20090 ( .A(n17785), .B(n17784), .Y(n17786) );
  NAND2XL U20091 ( .A(n17783), .B(n17827), .Y(n17784) );
  MXI2XL U20092 ( .A(Q5[2]), .B(n17836), .S0(n24128), .Y(n3990) );
  XNOR2XL U20093 ( .A(n17899), .B(n17835), .Y(n17836) );
  NAND2XL U20094 ( .A(n17878), .B(n17897), .Y(n17835) );
  MXI2XL U20095 ( .A(Q5[3]), .B(n17884), .S0(n24128), .Y(n3991) );
  XOR2XL U20096 ( .A(n17883), .B(n17882), .Y(n17884) );
  NAND2XL U20097 ( .A(n17881), .B(n17896), .Y(n17882) );
  AOI21XL U20098 ( .A0(n17899), .A1(n17878), .B0(n17877), .Y(n17883) );
  MXI2XL U20099 ( .A(Q5[4]), .B(n17904), .S0(n24128), .Y(n3992) );
  XOR2XL U20100 ( .A(n17969), .B(n17903), .Y(n17904) );
  NAND2XL U20101 ( .A(n17902), .B(n18027), .Y(n17903) );
  INVXL U20102 ( .A(n18024), .Y(n17902) );
  MXI2XL U20103 ( .A(Q5[5]), .B(n17975), .S0(n24128), .Y(n3993) );
  XNOR2XL U20104 ( .A(n17974), .B(n17973), .Y(n17975) );
  NAND2XL U20105 ( .A(n17972), .B(n18026), .Y(n17973) );
  MXI2XL U20106 ( .A(Q5[6]), .B(n18039), .S0(U1_valid[1]), .Y(n3994) );
  XOR2XL U20107 ( .A(n18204), .B(n18038), .Y(n18039) );
  NAND2XL U20108 ( .A(n18037), .B(n18128), .Y(n18038) );
  INVXL U20109 ( .A(n18126), .Y(n18037) );
  MXI2XL U20110 ( .A(Q5[7]), .B(n18063), .S0(U1_valid[1]), .Y(n3995) );
  XNOR2XL U20111 ( .A(n18062), .B(n18061), .Y(n18063) );
  NAND2XL U20112 ( .A(n18060), .B(n18127), .Y(n18061) );
  MXI2XL U20113 ( .A(Q5[8]), .B(n18135), .S0(U1_valid[1]), .Y(n3996) );
  MXI2XL U20114 ( .A(Q5[9]), .B(n18184), .S0(n18351), .Y(n3997) );
  XOR2XL U20115 ( .A(n18183), .B(n18182), .Y(n18184) );
  NAND2XL U20116 ( .A(n18181), .B(n18198), .Y(n18182) );
  AOI21XL U20117 ( .A0(n18178), .A1(n18177), .B0(n18176), .Y(n18183) );
  MXI2XL U20118 ( .A(Q5[10]), .B(n18208), .S0(n18351), .Y(n3998) );
  XOR2XL U20119 ( .A(n18347), .B(n18207), .Y(n18208) );
  NAND2XL U20120 ( .A(n18291), .B(n18343), .Y(n18207) );
  MXI2XL U20121 ( .A(Q5[11]), .B(n18298), .S0(n18351), .Y(n3999) );
  XOR2XL U20122 ( .A(n18297), .B(n18296), .Y(n18298) );
  NAND2XL U20123 ( .A(n18295), .B(n18342), .Y(n18296) );
  AOI21XL U20124 ( .A0(n18292), .A1(n18291), .B0(n18290), .Y(n18297) );
  MXI2XL U20125 ( .A(Q5[12]), .B(n18352), .S0(n18351), .Y(n4000) );
  XNOR2XL U20126 ( .A(n18379), .B(n18350), .Y(n18352) );
  NAND2XL U20127 ( .A(n18378), .B(n18466), .Y(n18350) );
  MXI2XL U20128 ( .A(Q5[13]), .B(n18385), .S0(n24128), .Y(n4001) );
  XOR2XL U20129 ( .A(n18384), .B(n18383), .Y(n18385) );
  NAND2XL U20130 ( .A(n18382), .B(n18465), .Y(n18383) );
  AOI21XL U20131 ( .A0(n18379), .A1(n18378), .B0(n18377), .Y(n18384) );
  MXI2XL U20132 ( .A(Q5[14]), .B(n18480), .S0(n24128), .Y(n4002) );
  XNOR2XL U20133 ( .A(n18671), .B(n18479), .Y(n18480) );
  NAND2XL U20134 ( .A(n18537), .B(n18563), .Y(n18479) );
  MXI2XL U20135 ( .A(Q5[15]), .B(n18543), .S0(n24128), .Y(n4003) );
  XOR2XL U20136 ( .A(n18542), .B(n18541), .Y(n18543) );
  NAND2XL U20137 ( .A(n18540), .B(n18562), .Y(n18541) );
  AOI21XL U20138 ( .A0(n18671), .A1(n18537), .B0(n18536), .Y(n18542) );
  MXI2XL U20139 ( .A(Q5[16]), .B(n18570), .S0(n18739), .Y(n4004) );
  XOR2XL U20140 ( .A(n18569), .B(n18568), .Y(n18570) );
  NAND2XL U20141 ( .A(n18565), .B(n18638), .Y(n18568) );
  AOI21XL U20142 ( .A0(n18671), .A1(n18637), .B0(n18640), .Y(n18569) );
  MXI2XL U20143 ( .A(Q5[17]), .B(n18648), .S0(n18739), .Y(n4005) );
  XOR2XL U20144 ( .A(n18647), .B(n18646), .Y(n18648) );
  NAND2XL U20145 ( .A(n18645), .B(n18668), .Y(n18646) );
  AOI21XL U20146 ( .A0(n18671), .A1(n18642), .B0(n18641), .Y(n18647) );
  MXI2XL U20147 ( .A(Q5[18]), .B(n18677), .S0(n18739), .Y(n4006) );
  XOR2XL U20148 ( .A(n18676), .B(n18675), .Y(n18677) );
  NAND2XL U20149 ( .A(n18672), .B(n18729), .Y(n18675) );
  AOI21XL U20150 ( .A0(n18671), .A1(n18728), .B0(n18731), .Y(n18676) );
  MXI2XL U20151 ( .A(Q5[19]), .B(n18740), .S0(n18739), .Y(n4007) );
  XNOR2XL U20152 ( .A(n18800), .B(n18738), .Y(n18740) );
  NAND2XL U20153 ( .A(n18735), .B(n18798), .Y(n18738) );
  MXI2XL U20154 ( .A(Q5[20]), .B(n18805), .S0(n18893), .Y(n4008) );
  NAND2XL U20155 ( .A(n18803), .B(n18832), .Y(n18804) );
  INVXL U20156 ( .A(n18833), .Y(n18803) );
  MXI2XL U20157 ( .A(Q5[21]), .B(n18839), .S0(n18893), .Y(n4009) );
  XNOR2XL U20158 ( .A(n18880), .B(n18838), .Y(n18839) );
  NAND2XL U20159 ( .A(n18835), .B(n18878), .Y(n18838) );
  MXI2XL U20160 ( .A(Q5[22]), .B(n18885), .S0(n18893), .Y(n4010) );
  XOR2XL U20161 ( .A(n18921), .B(n18884), .Y(n18885) );
  NAND2XL U20162 ( .A(n18883), .B(n18919), .Y(n18884) );
  INVXL U20163 ( .A(n18920), .Y(n18883) );
  MXI2XL U20164 ( .A(Q5[23]), .B(n18926), .S0(U1_valid[1]), .Y(n4011) );
  XNOR2XL U20165 ( .A(n18957), .B(n18925), .Y(n18926) );
  NAND2XL U20166 ( .A(n18922), .B(n18955), .Y(n18925) );
  MXI2XL U20167 ( .A(Q5[24]), .B(n18962), .S0(U1_valid[1]), .Y(n4012) );
  XOR2XL U20168 ( .A(n19011), .B(n18961), .Y(n18962) );
  NAND2XL U20169 ( .A(n18960), .B(n19009), .Y(n18961) );
  INVXL U20170 ( .A(n19010), .Y(n18960) );
  XOR2XL U20171 ( .A(n28695), .B(n28991), .Y(n19014) );
  MXI2XL U20172 ( .A(Q6[28]), .B(n19384), .S0(n23239), .Y(n4014) );
  XOR2XL U20173 ( .A(n19383), .B(n20476), .Y(n19384) );
  NAND2XL U20174 ( .A(n19379), .B(n20474), .Y(n19383) );
  INVXL U20175 ( .A(n20475), .Y(n19379) );
  MXI2XL U20176 ( .A(Q6[29]), .B(n20481), .S0(n24128), .Y(n4015) );
  XOR2XL U20177 ( .A(n20515), .B(n20480), .Y(n20481) );
  NAND2XL U20178 ( .A(n20479), .B(n20592), .Y(n20480) );
  INVXL U20179 ( .A(n20590), .Y(n20479) );
  MXI2XL U20180 ( .A(Q6[30]), .B(n20521), .S0(n24128), .Y(n4016) );
  XNOR2XL U20181 ( .A(n20520), .B(n20519), .Y(n20521) );
  NAND2XL U20182 ( .A(n20518), .B(n20591), .Y(n20519) );
  MXI2XL U20183 ( .A(Q6[31]), .B(n20600), .S0(n23239), .Y(n4017) );
  XNOR2XL U20184 ( .A(n20661), .B(n20599), .Y(n20600) );
  NAND2XL U20185 ( .A(n20612), .B(n20659), .Y(n20599) );
  MXI2XL U20186 ( .A(Q6[32]), .B(n20618), .S0(n23239), .Y(n4018) );
  XOR2XL U20187 ( .A(n20617), .B(n20616), .Y(n20618) );
  NAND2XL U20188 ( .A(n20615), .B(n20658), .Y(n20616) );
  AOI21XL U20189 ( .A0(n20661), .A1(n20612), .B0(n20611), .Y(n20617) );
  MXI2XL U20190 ( .A(Q6[33]), .B(n20666), .S0(n23239), .Y(n4019) );
  XOR2XL U20191 ( .A(n20733), .B(n20665), .Y(n20666) );
  NAND2XL U20192 ( .A(n20664), .B(n20799), .Y(n20665) );
  INVXL U20193 ( .A(n20796), .Y(n20664) );
  MXI2XL U20194 ( .A(Q6[34]), .B(n20739), .S0(n24128), .Y(n4020) );
  XNOR2XL U20195 ( .A(n20738), .B(n20737), .Y(n20739) );
  NAND2XL U20196 ( .A(n20736), .B(n20798), .Y(n20737) );
  MXI2XL U20197 ( .A(Q6[35]), .B(n20811), .S0(n23239), .Y(n4021) );
  XOR2XL U20198 ( .A(n21008), .B(n20810), .Y(n20811) );
  NAND2XL U20199 ( .A(n20809), .B(n20862), .Y(n20810) );
  INVXL U20200 ( .A(n20860), .Y(n20809) );
  MXI2XL U20201 ( .A(Q6[36]), .B(n20825), .S0(n23239), .Y(n4022) );
  MXI2XL U20202 ( .A(Q6[37]), .B(n20869), .S0(n24128), .Y(n4023) );
  XNOR2XL U20203 ( .A(n20912), .B(n20868), .Y(n20869) );
  NAND2XL U20204 ( .A(n20911), .B(n21003), .Y(n20868) );
  MXI2XL U20205 ( .A(Q6[38]), .B(n20918), .S0(n24128), .Y(n4024) );
  XOR2XL U20206 ( .A(n20917), .B(n20916), .Y(n20918) );
  NAND2XL U20207 ( .A(n20915), .B(n21002), .Y(n20916) );
  AOI21XL U20208 ( .A0(n20912), .A1(n20911), .B0(n20910), .Y(n20917) );
  MXI2XL U20209 ( .A(Q6[39]), .B(n21012), .S0(n23239), .Y(n4025) );
  XOR2XL U20210 ( .A(n21113), .B(n21011), .Y(n21012) );
  NAND2XL U20211 ( .A(n21055), .B(n21109), .Y(n21011) );
  MXI2XL U20212 ( .A(Q6[40]), .B(n21062), .S0(n24128), .Y(n4026) );
  XOR2XL U20213 ( .A(n21061), .B(n21060), .Y(n21062) );
  NAND2XL U20214 ( .A(n21059), .B(n21108), .Y(n21060) );
  AOI21XL U20215 ( .A0(n21056), .A1(n21055), .B0(n21054), .Y(n21061) );
  MXI2XL U20216 ( .A(Q4[29]), .B(n20488), .S0(n23239), .Y(n4027) );
  XNOR2XL U20217 ( .A(n20487), .B(n20486), .Y(n20488) );
  NAND2XL U20218 ( .A(n20485), .B(n20523), .Y(n20486) );
  MXI2XL U20219 ( .A(Q4[31]), .B(n20578), .S0(n24128), .Y(n4028) );
  XOR2XL U20220 ( .A(n20577), .B(n20576), .Y(n20578) );
  NAND2XL U20221 ( .A(n20575), .B(n20620), .Y(n20576) );
  AOI21XL U20222 ( .A0(n20623), .A1(n20572), .B0(n20571), .Y(n20577) );
  MXI2XL U20223 ( .A(Q4[32]), .B(n20628), .S0(n24128), .Y(n4029) );
  XOR2XL U20224 ( .A(n20667), .B(n20627), .Y(n20628) );
  NAND2XL U20225 ( .A(n20626), .B(n20713), .Y(n20627) );
  INVXL U20226 ( .A(n20710), .Y(n20626) );
  MXI2XL U20227 ( .A(Q4[33]), .B(n20673), .S0(n23239), .Y(n4030) );
  XNOR2XL U20228 ( .A(n20672), .B(n20671), .Y(n20673) );
  NAND2XL U20229 ( .A(n20670), .B(n20712), .Y(n20671) );
  MXI2XL U20230 ( .A(Q4[34]), .B(n20725), .S0(n23239), .Y(n4031) );
  XOR2XL U20231 ( .A(n20927), .B(n20724), .Y(n20725) );
  NAND2XL U20232 ( .A(n20723), .B(n20828), .Y(n20724) );
  INVXL U20233 ( .A(n20826), .Y(n20723) );
  MXI2XL U20234 ( .A(Q4[35]), .B(n20779), .S0(n24128), .Y(n4032) );
  XNOR2XL U20235 ( .A(n20778), .B(n20777), .Y(n20779) );
  NAND2XL U20236 ( .A(n20776), .B(n20827), .Y(n20777) );
  MXI2XL U20237 ( .A(Q4[36]), .B(n20835), .S0(n23239), .Y(n4033) );
  XNOR2XL U20238 ( .A(n20872), .B(n20834), .Y(n20835) );
  NAND2XL U20239 ( .A(n20871), .B(n20922), .Y(n20834) );
  MXI2XL U20240 ( .A(Q4[37]), .B(n20878), .S0(n23239), .Y(n4034) );
  XOR2XL U20241 ( .A(n20877), .B(n20876), .Y(n20878) );
  NAND2XL U20242 ( .A(n20875), .B(n20921), .Y(n20876) );
  AOI21XL U20243 ( .A0(n20872), .A1(n20871), .B0(n20870), .Y(n20877) );
  MXI2XL U20244 ( .A(Q4[38]), .B(n20931), .S0(n23239), .Y(n4035) );
  MXI2XL U20245 ( .A(Q4[39]), .B(n20999), .S0(n24128), .Y(n4036) );
  XOR2XL U20246 ( .A(n20998), .B(n20997), .Y(n20999) );
  NAND2XL U20247 ( .A(n20996), .B(n21044), .Y(n20997) );
  AOI21XL U20248 ( .A0(n20993), .A1(n20992), .B0(n20991), .Y(n20998) );
  MXI2XL U20249 ( .A(Q4[40]), .B(n21053), .S0(n24128), .Y(n4037) );
  XNOR2XL U20250 ( .A(n21100), .B(n21052), .Y(n21053) );
  NAND2XL U20251 ( .A(n21099), .B(n21151), .Y(n21052) );
  MXI2XL U20252 ( .A(Q4[41]), .B(n21106), .S0(n23239), .Y(n4038) );
  XOR2XL U20253 ( .A(n21105), .B(n21104), .Y(n21106) );
  NAND2XL U20254 ( .A(n21103), .B(n21150), .Y(n21104) );
  AOI21XL U20255 ( .A0(n21100), .A1(n21099), .B0(n21098), .Y(n21105) );
  MXI2XL U20256 ( .A(Q4[42]), .B(n21165), .S0(n23239), .Y(n4039) );
  XNOR2XL U20257 ( .A(n21395), .B(n21164), .Y(n21165) );
  NAND2XL U20258 ( .A(n21237), .B(n21289), .Y(n21164) );
  MXI2XL U20259 ( .A(Q4[43]), .B(n21243), .S0(n24128), .Y(n4040) );
  XOR2XL U20260 ( .A(n21242), .B(n21241), .Y(n21243) );
  NAND2XL U20261 ( .A(n21240), .B(n21288), .Y(n21241) );
  AOI21XL U20262 ( .A0(n21395), .A1(n21237), .B0(n21236), .Y(n21242) );
  MXI2XL U20263 ( .A(Q4[44]), .B(n21296), .S0(n24128), .Y(n4041) );
  XOR2XL U20264 ( .A(n21295), .B(n21294), .Y(n21296) );
  NAND2XL U20265 ( .A(n21291), .B(n21338), .Y(n21294) );
  AOI21XL U20266 ( .A0(n21395), .A1(n21337), .B0(n21340), .Y(n21295) );
  MXI2XL U20267 ( .A(Q4[45]), .B(n21348), .S0(n24128), .Y(n4042) );
  XOR2XL U20268 ( .A(n21347), .B(n21346), .Y(n21348) );
  NAND2XL U20269 ( .A(n21345), .B(n21392), .Y(n21346) );
  AOI21XL U20270 ( .A0(n21395), .A1(n21342), .B0(n21341), .Y(n21347) );
  MXI2XL U20271 ( .A(Q4[46]), .B(n21401), .S0(n23239), .Y(n4043) );
  XOR2XL U20272 ( .A(n21400), .B(n21399), .Y(n21401) );
  NAND2XL U20273 ( .A(n21396), .B(n21454), .Y(n21399) );
  AOI21XL U20274 ( .A0(n21395), .A1(n21453), .B0(n21456), .Y(n21400) );
  MXI2XL U20275 ( .A(Q4[47]), .B(n21464), .S0(n24128), .Y(n4044) );
  XNOR2XL U20276 ( .A(n21504), .B(n21463), .Y(n21464) );
  NAND2XL U20277 ( .A(n21460), .B(n21502), .Y(n21463) );
  MXI2XL U20278 ( .A(Q4[48]), .B(n21509), .S0(n24128), .Y(n4045) );
  XOR2XL U20279 ( .A(n21554), .B(n21508), .Y(n21509) );
  NAND2XL U20280 ( .A(n21507), .B(n21552), .Y(n21508) );
  INVXL U20281 ( .A(n21553), .Y(n21507) );
  MXI2XL U20282 ( .A(Q4[49]), .B(n21559), .S0(n23239), .Y(n4046) );
  XNOR2XL U20283 ( .A(n21598), .B(n21558), .Y(n21559) );
  NAND2XL U20284 ( .A(n21555), .B(n21596), .Y(n21558) );
  MXI2XL U20285 ( .A(Q4[50]), .B(n21603), .S0(n23239), .Y(n4047) );
  XOR2XL U20286 ( .A(n21640), .B(n21602), .Y(n21603) );
  NAND2XL U20287 ( .A(n21601), .B(n21638), .Y(n21602) );
  INVXL U20288 ( .A(n21639), .Y(n21601) );
  MXI2XL U20289 ( .A(Q4[51]), .B(n21645), .S0(n23239), .Y(n4048) );
  XNOR2XL U20290 ( .A(n21678), .B(n21644), .Y(n21645) );
  NAND2XL U20291 ( .A(n21641), .B(n21676), .Y(n21644) );
  MXI2XL U20292 ( .A(Q4[52]), .B(n21683), .S0(n23239), .Y(n4049) );
  XOR2XL U20293 ( .A(n21718), .B(n21682), .Y(n21683) );
  NAND2XL U20294 ( .A(n21681), .B(n21716), .Y(n21682) );
  INVXL U20295 ( .A(n21717), .Y(n21681) );
  XOR2XL U20296 ( .A(n28693), .B(n28989), .Y(n21721) );
  MXI2XL U20297 ( .A(Q4[30]), .B(n20532), .S0(n23239), .Y(n4051) );
  XNOR2XL U20298 ( .A(n20623), .B(n20531), .Y(n20532) );
  NAND2XL U20299 ( .A(n20572), .B(n20621), .Y(n20531) );
  MXI2XL U20300 ( .A(CQ0[31]), .B(U2_pipe0[5]), .S0(U2_valid_1_), .Y(n4052) );
  XOR2XL U20301 ( .A(n25991), .B(n25990), .Y(n25992) );
  NAND2XL U20302 ( .A(n25989), .B(n26031), .Y(n25990) );
  AOI21XL U20303 ( .A0(n26034), .A1(n25984), .B0(n25983), .Y(n25991) );
  MXI2XL U20304 ( .A(CQ0[32]), .B(U2_pipe0[6]), .S0(U2_valid_1_), .Y(n4054) );
  XOR2XL U20305 ( .A(n26079), .B(n26040), .Y(n26041) );
  NAND2XL U20306 ( .A(n26039), .B(n26145), .Y(n26040) );
  INVXL U20307 ( .A(n26142), .Y(n26039) );
  MXI2XL U20308 ( .A(CQ0[33]), .B(U2_pipe0[7]), .S0(U2_valid_1_), .Y(n4056) );
  XNOR2XL U20309 ( .A(n26086), .B(n26085), .Y(n26087) );
  NAND2XL U20310 ( .A(n26084), .B(n26144), .Y(n26085) );
  MXI2XL U20311 ( .A(CQ0[34]), .B(U2_pipe0[8]), .S0(U2_valid_1_), .Y(n4058) );
  XOR2XL U20312 ( .A(n26354), .B(n26158), .Y(n26159) );
  INVXL U20313 ( .A(n26235), .Y(n26157) );
  MXI2XL U20314 ( .A(CQ0[35]), .B(U2_pipe0[9]), .S0(U2_valid_1_), .Y(n4060) );
  MXI2XL U20315 ( .A(CQ0[36]), .B(U2_pipe0[10]), .S0(U2_valid_1_), .Y(n4062)
         );
  MXI2XL U20316 ( .A(CQ0[37]), .B(U2_pipe0[11]), .S0(U2_valid_1_), .Y(n4064)
         );
  NAND2XL U20317 ( .A(n26294), .B(n26348), .Y(n26295) );
  AOI21XL U20318 ( .A0(n26289), .A1(n26288), .B0(n26287), .Y(n26296) );
  MXI2XL U20319 ( .A(CQ0[38]), .B(U2_pipe0[12]), .S0(U2_valid_1_), .Y(n4066)
         );
  MXI2XL U20320 ( .A(CQ0[39]), .B(U2_pipe0[13]), .S0(n27042), .Y(n4068) );
  AOI21XL U20321 ( .A0(n26402), .A1(n26401), .B0(n26400), .Y(n26409) );
  MXI2XL U20322 ( .A(CQ0[40]), .B(U2_pipe0[14]), .S0(n27042), .Y(n4070) );
  MXI2XL U20323 ( .A(CQ0[41]), .B(U2_pipe0[15]), .S0(n27042), .Y(n4072) );
  NAND2XL U20324 ( .A(n26519), .B(n26594), .Y(n26520) );
  MXI2XL U20325 ( .A(CQ0[42]), .B(U2_pipe0[16]), .S0(n27042), .Y(n4074) );
  MXI2XL U20326 ( .A(CQ0[43]), .B(U2_pipe0[17]), .S0(n27042), .Y(n4076) );
  MXI2XL U20327 ( .A(CQ0[44]), .B(U2_pipe0[18]), .S0(n27042), .Y(n4078) );
  MXI2XL U20328 ( .A(CQ0[45]), .B(U2_pipe0[19]), .S0(n27042), .Y(n4080) );
  NAND2XL U20329 ( .A(n26763), .B(n26816), .Y(n26764) );
  MXI2XL U20330 ( .A(CQ0[46]), .B(U2_pipe0[20]), .S0(n27042), .Y(n4082) );
  NAND2XL U20331 ( .A(n26821), .B(n26860), .Y(n26824) );
  MXI2XL U20332 ( .A(CQ0[47]), .B(U2_pipe0[21]), .S0(n27042), .Y(n4084) );
  NAND2XL U20333 ( .A(n26906), .B(n26904), .Y(n26870) );
  MXI2XL U20334 ( .A(CQ0[48]), .B(U2_pipe0[22]), .S0(n27042), .Y(n4086) );
  AND2XL U20335 ( .A(n26912), .B(n26946), .Y(n7026) );
  OAI2BB1X1 U20336 ( .A0N(n26906), .A1N(n26907), .B0(n26904), .Y(n7541) );
  MXI2XL U20337 ( .A(CQ0[49]), .B(U2_pipe0[23]), .S0(n27042), .Y(n4088) );
  XNOR2X1 U20338 ( .A(n26989), .B(n26952), .Y(n26953) );
  NAND2XL U20339 ( .A(n26988), .B(n26986), .Y(n26952) );
  MXI2XL U20340 ( .A(CQ0[50]), .B(U2_pipe0[24]), .S0(n27042), .Y(n4090) );
  XOR2X1 U20341 ( .A(n27031), .B(n26995), .Y(n26996) );
  NAND2XL U20342 ( .A(n26994), .B(n27029), .Y(n26995) );
  INVXL U20343 ( .A(n27030), .Y(n26994) );
  MXI2XL U20344 ( .A(CQ0[51]), .B(U2_pipe0[25]), .S0(n27042), .Y(n4092) );
  NAND2XL U20345 ( .A(n27037), .B(n27036), .Y(n27038) );
  MXI2XL U20346 ( .A(CQ0[0]), .B(U2_pipe1[0]), .S0(U2_valid_1_), .Y(n4094) );
  MXI2XL U20347 ( .A(U2_pipe1[0]), .B(n21733), .S0(n23695), .Y(n4095) );
  XNOR2XL U20348 ( .A(n21732), .B(n21731), .Y(n21733) );
  NAND2XL U20349 ( .A(n23166), .B(n23167), .Y(n21731) );
  MXI2XL U20350 ( .A(CQ0[1]), .B(U2_pipe1[1]), .S0(U2_valid_1_), .Y(n4096) );
  MXI2XL U20351 ( .A(U2_pipe1[1]), .B(n23136), .S0(n23695), .Y(n4097) );
  XNOR2XL U20352 ( .A(n23135), .B(n23134), .Y(n23136) );
  NAND2XL U20353 ( .A(n23171), .B(n23168), .Y(n23134) );
  MXI2XL U20354 ( .A(CQ0[2]), .B(U2_pipe1[2]), .S0(U2_valid_1_), .Y(n4098) );
  MXI2XL U20355 ( .A(U2_pipe1[2]), .B(n23182), .S0(n23695), .Y(n4099) );
  XOR2XL U20356 ( .A(n23223), .B(n23181), .Y(n23182) );
  NAND2XL U20357 ( .A(n23180), .B(n23270), .Y(n23181) );
  INVXL U20358 ( .A(n23268), .Y(n23180) );
  MXI2XL U20359 ( .A(CQ0[3]), .B(U2_pipe1[3]), .S0(U2_valid_1_), .Y(n4100) );
  XNOR2XL U20360 ( .A(n23230), .B(n23229), .Y(n23231) );
  NAND2XL U20361 ( .A(n23228), .B(n23269), .Y(n23229) );
  MXI2XL U20362 ( .A(CQ0[4]), .B(U2_pipe1[4]), .S0(U2_valid_1_), .Y(n4102) );
  XNOR2XL U20363 ( .A(n23364), .B(n23279), .Y(n23280) );
  NAND2XL U20364 ( .A(n23320), .B(n23362), .Y(n23279) );
  MXI2XL U20365 ( .A(CQ0[5]), .B(U2_pipe1[5]), .S0(U2_valid_1_), .Y(n4104) );
  XOR2XL U20366 ( .A(n23327), .B(n23326), .Y(n23328) );
  NAND2XL U20367 ( .A(n23325), .B(n23361), .Y(n23326) );
  AOI21XL U20368 ( .A0(n23364), .A1(n23320), .B0(n23319), .Y(n23327) );
  MXI2XL U20369 ( .A(CQ0[6]), .B(U2_pipe1[6]), .S0(U2_valid_1_), .Y(n4106) );
  XOR2XL U20370 ( .A(n23427), .B(n23370), .Y(n23371) );
  NAND2XL U20371 ( .A(n23369), .B(n23473), .Y(n23370) );
  INVXL U20372 ( .A(n23470), .Y(n23369) );
  MXI2XL U20373 ( .A(CQ0[7]), .B(U2_pipe1[7]), .S0(n27042), .Y(n4108) );
  XNOR2XL U20374 ( .A(n23434), .B(n23433), .Y(n23435) );
  NAND2XL U20375 ( .A(n23432), .B(n23472), .Y(n23433) );
  MXI2XL U20376 ( .A(CQ0[8]), .B(U2_pipe1[8]), .S0(n27042), .Y(n4110) );
  INVXL U20377 ( .A(n23570), .Y(n23485) );
  MXI2XL U20378 ( .A(CQ0[9]), .B(U2_pipe1[9]), .S0(n27042), .Y(n4112) );
  XNOR2XL U20379 ( .A(n23530), .B(n23529), .Y(n23531) );
  NAND2XL U20380 ( .A(n23528), .B(n23571), .Y(n23529) );
  MXI2XL U20381 ( .A(CQ0[10]), .B(U2_pipe1[10]), .S0(n27042), .Y(n4114) );
  MXI2XL U20382 ( .A(CQ0[11]), .B(U2_pipe1[11]), .S0(n27042), .Y(n4116) );
  NAND2XL U20383 ( .A(n23637), .B(n23683), .Y(n23638) );
  MXI2XL U20384 ( .A(CQ0[12]), .B(U2_pipe1[12]), .S0(n27042), .Y(n4118) );
  MXI2XL U20385 ( .A(CQ0[13]), .B(U2_pipe1[13]), .S0(n24380), .Y(n4120) );
  XOR2XL U20386 ( .A(n23748), .B(n23747), .Y(n23749) );
  MXI2XL U20387 ( .A(CQ0[14]), .B(U2_pipe1[14]), .S0(n24380), .Y(n4122) );
  XNOR2X1 U20388 ( .A(n23869), .B(n23799), .Y(n23800) );
  MXI2XL U20389 ( .A(CQ0[15]), .B(U2_pipe1[15]), .S0(n24380), .Y(n4124) );
  NAND2XL U20390 ( .A(n23874), .B(n23925), .Y(n23875) );
  MXI2XL U20391 ( .A(CQ0[16]), .B(U2_pipe1[16]), .S0(n24380), .Y(n4126) );
  MXI2XL U20392 ( .A(CQ0[17]), .B(U2_pipe1[17]), .S0(n24380), .Y(n4128) );
  MXI2XL U20393 ( .A(CQ0[18]), .B(U2_pipe1[18]), .S0(n24380), .Y(n4130) );
  NAND2XL U20394 ( .A(n6986), .B(n24092), .Y(n24044) );
  MXI2XL U20395 ( .A(CQ0[19]), .B(U2_pipe1[19]), .S0(n24380), .Y(n4132) );
  NAND2XL U20396 ( .A(n24101), .B(n24155), .Y(n24102) );
  MXI2XL U20397 ( .A(CQ0[20]), .B(U2_pipe1[20]), .S0(n24380), .Y(n4134) );
  NAND2XL U20398 ( .A(n24161), .B(n24200), .Y(n24164) );
  MXI2XL U20399 ( .A(CQ0[21]), .B(U2_pipe1[21]), .S0(n24380), .Y(n4136) );
  XNOR2X1 U20400 ( .A(n24247), .B(n24210), .Y(n24211) );
  NAND2XL U20401 ( .A(n24246), .B(n24244), .Y(n24210) );
  MXI2XL U20402 ( .A(CQ0[22]), .B(U2_pipe1[22]), .S0(n24380), .Y(n4138) );
  NAND2XL U20403 ( .A(n7383), .B(n24286), .Y(n24252) );
  MXI2XL U20404 ( .A(CQ0[23]), .B(U2_pipe1[23]), .S0(n24380), .Y(n4140) );
  XNOR2X1 U20405 ( .A(n24330), .B(n24293), .Y(n24294) );
  NAND2XL U20406 ( .A(n24329), .B(n24327), .Y(n24293) );
  MXI2XL U20407 ( .A(CQ0[24]), .B(U2_pipe1[24]), .S0(n24380), .Y(n4142) );
  NAND2XL U20408 ( .A(n24335), .B(n24370), .Y(n24336) );
  INVXL U20409 ( .A(n24371), .Y(n24335) );
  MXI2XL U20410 ( .A(CQ0[25]), .B(U2_pipe1[25]), .S0(n24380), .Y(n4144) );
  MXI2XL U20411 ( .A(CQ1[26]), .B(U2_pipe2[0]), .S0(n24380), .Y(n4146) );
  MXI2XL U20412 ( .A(U2_pipe2[0]), .B(n19068), .S0(n21023), .Y(n4147) );
  XNOR2XL U20413 ( .A(n25845), .B(n19067), .Y(n19068) );
  NAND2XL U20414 ( .A(n19066), .B(n20466), .Y(n19067) );
  INVXL U20415 ( .A(n20467), .Y(n19066) );
  MXI2XL U20416 ( .A(CQ1[27]), .B(U2_pipe2[1]), .S0(n24380), .Y(n4148) );
  MXI2XL U20417 ( .A(U2_pipe2[1]), .B(n20473), .S0(n21023), .Y(n4149) );
  XOR2XL U20418 ( .A(n20505), .B(n20472), .Y(n20473) );
  NAND2XL U20419 ( .A(n20471), .B(n20549), .Y(n20472) );
  INVXL U20420 ( .A(n20547), .Y(n20471) );
  MXI2XL U20421 ( .A(CQ1[28]), .B(U2_pipe2[2]), .S0(n27042), .Y(n4150) );
  MXI2XL U20422 ( .A(U2_pipe2[2]), .B(n20514), .S0(n21023), .Y(n4151) );
  XNOR2XL U20423 ( .A(n20513), .B(n20512), .Y(n20514) );
  NAND2XL U20424 ( .A(n20511), .B(n20548), .Y(n20512) );
  MXI2XL U20425 ( .A(CQ1[29]), .B(U2_pipe2[3]), .S0(n27042), .Y(n4152) );
  XNOR2XL U20426 ( .A(n20649), .B(n20558), .Y(n20559) );
  NAND2XL U20427 ( .A(n20602), .B(n20647), .Y(n20558) );
  MXI2XL U20428 ( .A(CQ1[30]), .B(U2_pipe2[4]), .S0(U2_valid_1_), .Y(n4154) );
  XOR2XL U20429 ( .A(n20609), .B(n20608), .Y(n20610) );
  NAND2XL U20430 ( .A(n20607), .B(n20646), .Y(n20608) );
  AOI21XL U20431 ( .A0(n20649), .A1(n20602), .B0(n20601), .Y(n20609) );
  MXI2XL U20432 ( .A(CQ1[31]), .B(U2_pipe2[5]), .S0(n27042), .Y(n4156) );
  XOR2XL U20433 ( .A(n20694), .B(n20655), .Y(n20656) );
  NAND2XL U20434 ( .A(n20654), .B(n20743), .Y(n20655) );
  MXI2XL U20435 ( .A(CQ1[32]), .B(U2_pipe2[6]), .S0(n24380), .Y(n4158) );
  XNOR2XL U20436 ( .A(n20701), .B(n20700), .Y(n20702) );
  NAND2XL U20437 ( .A(n20699), .B(n20742), .Y(n20700) );
  MXI2XL U20438 ( .A(CQ1[33]), .B(U2_pipe2[7]), .S0(U2_valid_1_), .Y(n4160) );
  XOR2XL U20439 ( .A(n20958), .B(n20756), .Y(n20757) );
  INVXL U20440 ( .A(n20848), .Y(n20755) );
  MXI2XL U20441 ( .A(CQ1[34]), .B(U2_pipe2[8]), .S0(n27042), .Y(n4162) );
  NAND2XL U20442 ( .A(n20816), .B(n20849), .Y(n20817) );
  MXI2XL U20443 ( .A(CQ1[35]), .B(U2_pipe2[9]), .S0(n27042), .Y(n4164) );
  MXI2XL U20444 ( .A(CQ1[36]), .B(U2_pipe2[10]), .S0(U2_valid_1_), .Y(n4166)
         );
  NAND2XL U20445 ( .A(n20906), .B(n20952), .Y(n20907) );
  AOI21XL U20446 ( .A0(n20901), .A1(n20900), .B0(n20899), .Y(n20908) );
  MXI2XL U20447 ( .A(CQ1[37]), .B(U2_pipe2[11]), .S0(n27042), .Y(n4168) );
  MXI2XL U20448 ( .A(CQ1[38]), .B(U2_pipe2[12]), .S0(n24380), .Y(n4170) );
  NAND2XL U20449 ( .A(n21020), .B(n21064), .Y(n21021) );
  MXI2XL U20450 ( .A(CQ1[39]), .B(U2_pipe2[13]), .S0(U2_valid_1_), .Y(n4172)
         );
  NAND2XL U20451 ( .A(n21119), .B(n21179), .Y(n21074) );
  MXI2XL U20452 ( .A(CQ1[40]), .B(U2_pipe2[14]), .S0(n24380), .Y(n4174) );
  NAND2XL U20453 ( .A(n21125), .B(n21178), .Y(n21126) );
  MXI2XL U20454 ( .A(CQ1[41]), .B(U2_pipe2[15]), .S0(n27042), .Y(n4176) );
  XNOR2X1 U20455 ( .A(n21528), .B(n21194), .Y(n21195) );
  MXI2XL U20456 ( .A(CQ1[42]), .B(U2_pipe2[16]), .S0(n27042), .Y(n4178) );
  MXI2XL U20457 ( .A(CQ1[43]), .B(U2_pipe2[17]), .S0(n27042), .Y(n4180) );
  NAND2XL U20458 ( .A(n21312), .B(n21416), .Y(n21313) );
  INVXL U20459 ( .A(n21413), .Y(n21312) );
  MXI2XL U20460 ( .A(CQ1[44]), .B(U2_pipe2[18]), .S0(U2_valid_1_), .Y(n4182)
         );
  NAND2XL U20461 ( .A(n21365), .B(n21415), .Y(n21366) );
  MXI2XL U20462 ( .A(CQ1[45]), .B(U2_pipe2[19]), .S0(U2_valid_1_), .Y(n4184)
         );
  NAND2XL U20463 ( .A(n21518), .B(n21520), .Y(n21427) );
  MXI2XL U20464 ( .A(CQ1[46]), .B(U2_pipe2[20]), .S0(n24380), .Y(n4186) );
  NAND2XL U20465 ( .A(n21524), .B(n21521), .Y(n21483) );
  MXI2XL U20466 ( .A(CQ1[47]), .B(U2_pipe2[21]), .S0(n27042), .Y(n4188) );
  NAND2XL U20467 ( .A(n5765), .B(n21569), .Y(n21533) );
  MXI2XL U20468 ( .A(CQ1[48]), .B(U2_pipe2[22]), .S0(n27042), .Y(n4190) );
  NAND2XL U20469 ( .A(n21575), .B(n21612), .Y(n21578) );
  MXI2XL U20470 ( .A(CQ1[49]), .B(U2_pipe2[23]), .S0(n24380), .Y(n4192) );
  XOR2X1 U20471 ( .A(n21658), .B(n21620), .Y(n21621) );
  NAND2XL U20472 ( .A(n21619), .B(n21656), .Y(n21620) );
  INVXL U20473 ( .A(n21657), .Y(n21619) );
  MXI2XL U20474 ( .A(CQ1[50]), .B(U2_pipe2[24]), .S0(n24380), .Y(n4194) );
  XOR2X1 U20475 ( .A(n7417), .B(n7416), .Y(n21659) );
  MXI2XL U20476 ( .A(CQ1[51]), .B(U2_pipe2[25]), .S0(U2_valid_1_), .Y(n4196)
         );
  MXI2XL U20477 ( .A(CQ1[0]), .B(U2_pipe3[0]), .S0(n24380), .Y(n4198) );
  MXI2XL U20478 ( .A(U2_pipe3[0]), .B(n16627), .S0(n8054), .Y(n4199) );
  NAND2XL U20479 ( .A(n16625), .B(n17750), .Y(n16626) );
  INVXL U20480 ( .A(n17751), .Y(n16625) );
  MXI2XL U20481 ( .A(CQ1[1]), .B(U2_pipe3[1]), .S0(n24380), .Y(n4200) );
  MXI2XL U20482 ( .A(U2_pipe3[1]), .B(n17757), .S0(n8054), .Y(n4201) );
  XOR2XL U20483 ( .A(n17787), .B(n17756), .Y(n17757) );
  NAND2XL U20484 ( .A(n17755), .B(n17839), .Y(n17756) );
  INVXL U20485 ( .A(n17837), .Y(n17755) );
  MXI2XL U20486 ( .A(CQ1[2]), .B(U2_pipe3[2]), .S0(n24380), .Y(n4202) );
  NAND2XL U20487 ( .A(n17793), .B(n17838), .Y(n17794) );
  MXI2XL U20488 ( .A(CQ1[3]), .B(U2_pipe3[3]), .S0(n24380), .Y(n4204) );
  XNOR2XL U20489 ( .A(n17937), .B(n17848), .Y(n17849) );
  NAND2XL U20490 ( .A(n17886), .B(n17935), .Y(n17848) );
  MXI2XL U20491 ( .A(CQ1[4]), .B(U2_pipe3[4]), .S0(n24380), .Y(n4206) );
  XOR2XL U20492 ( .A(n17893), .B(n17892), .Y(n17894) );
  NAND2XL U20493 ( .A(n17891), .B(n17934), .Y(n17892) );
  AOI21XL U20494 ( .A0(n17937), .A1(n17886), .B0(n17885), .Y(n17893) );
  MXI2XL U20495 ( .A(CQ1[5]), .B(U2_pipe3[5]), .S0(n24380), .Y(n4208) );
  XOR2XL U20496 ( .A(n17976), .B(n17943), .Y(n17944) );
  NAND2XL U20497 ( .A(n17942), .B(n18043), .Y(n17943) );
  MXI2XL U20498 ( .A(CQ1[6]), .B(U2_pipe3[6]), .S0(n24380), .Y(n4210) );
  NAND2XL U20499 ( .A(n17981), .B(n18042), .Y(n17982) );
  MXI2XL U20500 ( .A(CQ1[7]), .B(U2_pipe3[7]), .S0(n24380), .Y(n4212) );
  XOR2XL U20501 ( .A(n18252), .B(n18056), .Y(n18057) );
  NAND2XL U20502 ( .A(n18055), .B(n18138), .Y(n18056) );
  MXI2XL U20503 ( .A(CQ1[8]), .B(U2_pipe3[8]), .S0(n24380), .Y(n4214) );
  NAND2XL U20504 ( .A(n18096), .B(n18137), .Y(n18097) );
  MXI2XL U20505 ( .A(CQ1[9]), .B(U2_pipe3[9]), .S0(n24380), .Y(n4216) );
  MXI2XL U20506 ( .A(CQ1[10]), .B(U2_pipe3[10]), .S0(n24380), .Y(n4218) );
  NAND2XL U20507 ( .A(n18192), .B(n18246), .Y(n18193) );
  MXI2XL U20508 ( .A(CQ1[11]), .B(U2_pipe3[11]), .S0(n24380), .Y(n4220) );
  MXI2XL U20509 ( .A(CQ1[12]), .B(U2_pipe3[12]), .S0(n24380), .Y(n4222) );
  MXI2XL U20510 ( .A(CQ1[13]), .B(U2_pipe3[13]), .S0(n27042), .Y(n4224) );
  NAND2XL U20511 ( .A(n18405), .B(n18485), .Y(n18364) );
  MXI2XL U20512 ( .A(CQ1[14]), .B(U2_pipe3[14]), .S0(n24380), .Y(n4226) );
  NAND2XL U20513 ( .A(n18411), .B(n18484), .Y(n18412) );
  AOI21XL U20514 ( .A0(n18406), .A1(n18405), .B0(n18404), .Y(n18413) );
  MXI2XL U20515 ( .A(CQ1[15]), .B(U2_pipe3[15]), .S0(n27042), .Y(n4228) );
  MXI2XL U20516 ( .A(CQ1[16]), .B(U2_pipe3[16]), .S0(n24380), .Y(n4230) );
  MXI2XL U20517 ( .A(CQ1[17]), .B(U2_pipe3[17]), .S0(n27042), .Y(n4232) );
  NAND2XL U20518 ( .A(n18599), .B(n18703), .Y(n18600) );
  INVXL U20519 ( .A(n18700), .Y(n18599) );
  MXI2XL U20520 ( .A(CQ1[18]), .B(U2_pipe3[18]), .S0(n24380), .Y(n4234) );
  MXI2XL U20521 ( .A(CQ1[19]), .B(U2_pipe3[19]), .S0(n27042), .Y(n4236) );
  NAND2XL U20522 ( .A(n18806), .B(n18808), .Y(n18714) );
  MXI2XL U20523 ( .A(CQ1[20]), .B(U2_pipe3[20]), .S0(n24380), .Y(n4238) );
  NAND2XL U20524 ( .A(n18812), .B(n18809), .Y(n18771) );
  MXI2XL U20525 ( .A(CQ1[21]), .B(U2_pipe3[21]), .S0(n27042), .Y(n4240) );
  NAND2XL U20526 ( .A(n6935), .B(n18857), .Y(n18821) );
  MXI2XL U20527 ( .A(CQ1[22]), .B(U2_pipe3[22]), .S0(n24380), .Y(n4242) );
  XNOR2X1 U20528 ( .A(n18905), .B(n18868), .Y(n18869) );
  NAND2XL U20529 ( .A(n18865), .B(n18903), .Y(n18868) );
  MXI2XL U20530 ( .A(CQ1[23]), .B(U2_pipe3[23]), .S0(n27042), .Y(n4244) );
  AND2XL U20531 ( .A(n7050), .B(n18945), .Y(n7027) );
  MXI2XL U20532 ( .A(CQ1[24]), .B(U2_pipe3[24]), .S0(n24380), .Y(n4246) );
  MXI2XL U20533 ( .A(CQ1[25]), .B(U2_pipe3[25]), .S0(n27042), .Y(n4248) );
  MXI2XL U20534 ( .A(CQ0[26]), .B(U2_pipe0[0]), .S0(U2_valid_1_), .Y(n4250) );
  MXI2XL U20535 ( .A(U2_pipe0[0]), .B(n24412), .S0(n8054), .Y(n4251) );
  XNOR2XL U20536 ( .A(n24411), .B(n24410), .Y(n24412) );
  NAND2XL U20537 ( .A(n25837), .B(n25838), .Y(n24410) );
  MXI2XL U20538 ( .A(CQ0[28]), .B(U2_pipe0[2]), .S0(U2_valid_1_), .Y(n4252) );
  MXI2XL U20539 ( .A(U2_pipe0[2]), .B(n25853), .S0(n8054), .Y(n4253) );
  XOR2XL U20540 ( .A(n25886), .B(n25852), .Y(n25853) );
  NAND2XL U20541 ( .A(n25851), .B(n25938), .Y(n25852) );
  INVXL U20542 ( .A(n25936), .Y(n25851) );
  MXI2XL U20543 ( .A(CQ0[29]), .B(U2_pipe0[3]), .S0(U2_valid_1_), .Y(n4254) );
  MXI2XL U20544 ( .A(U2_pipe0[3]), .B(n25894), .S0(n8054), .Y(n4255) );
  XNOR2XL U20545 ( .A(n25893), .B(n25892), .Y(n25894) );
  NAND2XL U20546 ( .A(n25891), .B(n25937), .Y(n25892) );
  MXI2XL U20547 ( .A(CQ0[30]), .B(U2_pipe0[4]), .S0(U2_valid_1_), .Y(n4256) );
  XNOR2XL U20548 ( .A(n26034), .B(n25947), .Y(n25948) );
  NAND2XL U20549 ( .A(n25984), .B(n26032), .Y(n25947) );
  MXI2XL U20550 ( .A(CQ0[27]), .B(U2_pipe0[1]), .S0(U2_valid_1_), .Y(n4258) );
  MXI2XL U20551 ( .A(U2_pipe0[1]), .B(n25805), .S0(n8054), .Y(n4259) );
  XNOR2XL U20552 ( .A(n25804), .B(n25803), .Y(n25805) );
  NAND2XL U20553 ( .A(n25842), .B(n25839), .Y(n25803) );
  MXI2XL U20554 ( .A(U0_pipe0[4]), .B(n24970), .S0(n5920), .Y(n4260) );
  XNOR2XL U20555 ( .A(n24969), .B(n24968), .Y(n24970) );
  NAND2XL U20556 ( .A(n24967), .B(n24966), .Y(n24968) );
  XNOR2X1 U20557 ( .A(n24995), .B(n24994), .Y(n24996) );
  XNOR2X1 U20558 ( .A(n24999), .B(n24998), .Y(n25000) );
  XOR2X1 U20559 ( .A(n25004), .B(n25003), .Y(n25005) );
  INVXL U20560 ( .A(n25014), .Y(n25015) );
  INVXL U20561 ( .A(n25020), .Y(n25021) );
  XOR2X1 U20562 ( .A(n25019), .B(n25025), .Y(n25026) );
  NAND2XL U20563 ( .A(n25018), .B(n25024), .Y(n25025) );
  XOR2XL U20564 ( .A(n25036), .B(n25035), .Y(n25037) );
  XOR2XL U20565 ( .A(n25042), .B(n25041), .Y(n25043) );
  NAND2XL U20566 ( .A(n25040), .B(n25039), .Y(n25041) );
  XOR2XL U20567 ( .A(n25053), .B(n25052), .Y(n25054) );
  XNOR2XL U20568 ( .A(n25056), .B(n25055), .Y(n25057) );
  XOR2XL U20569 ( .A(n25064), .B(n25063), .Y(n25065) );
  AOI21XL U20570 ( .A0(n25067), .A1(n25062), .B0(n25061), .Y(n25064) );
  XNOR2XL U20571 ( .A(n25067), .B(n25066), .Y(n25068) );
  XOR2XL U20572 ( .A(n25070), .B(n25069), .Y(n25071) );
  XOR2XL U20573 ( .A(n25077), .B(n25076), .Y(n25078) );
  NAND2XL U20574 ( .A(n8839), .B(n25075), .Y(n25076) );
  XOR2XL U20575 ( .A(n25085), .B(n25084), .Y(n25086) );
  NAND2XL U20576 ( .A(n25083), .B(n25082), .Y(n25084) );
  AOI21XL U20577 ( .A0(n25090), .A1(n25088), .B0(n25080), .Y(n25085) );
  MXI2XL U20578 ( .A(U0_pipe1[5]), .B(n25092), .S0(n25091), .Y(n4279) );
  XNOR2XL U20579 ( .A(n25090), .B(n25089), .Y(n25092) );
  NAND2XL U20580 ( .A(n25088), .B(n25087), .Y(n25089) );
  MXI2XL U20581 ( .A(U0_pipe1[4]), .B(n25102), .S0(n25101), .Y(n4280) );
  XNOR2XL U20582 ( .A(n25100), .B(n25099), .Y(n25102) );
  NAND2XL U20583 ( .A(n25098), .B(n25097), .Y(n25099) );
  MXI2XL U20584 ( .A(U0_pipe1[3]), .B(n25105), .S0(n5810), .Y(n4281) );
  XOR2XL U20585 ( .A(n25104), .B(n25103), .Y(n25105) );
  MXI2XL U20586 ( .A(U0_pipe1[2]), .B(n25110), .S0(n5810), .Y(n4282) );
  XNOR2XL U20587 ( .A(n25109), .B(n25108), .Y(n25110) );
  MXI2XL U20588 ( .A(U0_pipe1[1]), .B(n25113), .S0(n5810), .Y(n4283) );
  MXI2XL U20589 ( .A(U0_pipe1[0]), .B(n25114), .S0(n5810), .Y(n4284) );
  NAND2XL U20590 ( .A(n24866), .B(n24865), .Y(n24867) );
  XOR2XL U20591 ( .A(n24909), .B(n24908), .Y(n24910) );
  XOR2XL U20592 ( .A(n24914), .B(n24913), .Y(n24915) );
  XNOR2XL U20593 ( .A(n24927), .B(n24926), .Y(n24928) );
  XOR2XL U20594 ( .A(n24935), .B(n24934), .Y(n24936) );
  AOI21XL U20595 ( .A0(n24938), .A1(n24933), .B0(n24932), .Y(n24935) );
  XNOR2XL U20596 ( .A(n24938), .B(n24937), .Y(n24939) );
  XOR2XL U20597 ( .A(n24941), .B(n24940), .Y(n24942) );
  XOR2XL U20598 ( .A(n24949), .B(n24948), .Y(n24950) );
  NAND2XL U20599 ( .A(n24947), .B(n24946), .Y(n24948) );
  XOR2XL U20600 ( .A(n24957), .B(n24956), .Y(n24958) );
  NAND2XL U20601 ( .A(n24955), .B(n24954), .Y(n24956) );
  AOI21XL U20602 ( .A0(n24962), .A1(n24960), .B0(n24952), .Y(n24957) );
  MXI2XL U20603 ( .A(U0_pipe0[5]), .B(n24963), .S0(n5920), .Y(n4307) );
  XNOR2XL U20604 ( .A(n24962), .B(n24961), .Y(n24963) );
  NAND2XL U20605 ( .A(n24960), .B(n24959), .Y(n24961) );
  MXI2XL U20606 ( .A(U0_pipe0[3]), .B(n24976), .S0(n5920), .Y(n4308) );
  XOR2XL U20607 ( .A(n24975), .B(n24974), .Y(n24976) );
  NAND2XL U20608 ( .A(n24973), .B(n24972), .Y(n24974) );
  INVXL U20609 ( .A(n24971), .Y(n24973) );
  XOR2XL U20610 ( .A(n22378), .B(n22377), .Y(n22379) );
  XNOR2XL U20611 ( .A(n22381), .B(n22380), .Y(n22382) );
  XOR2XL U20612 ( .A(n22384), .B(n22383), .Y(n22385) );
  MXI2XL U20613 ( .A(U0_pipe5[7]), .B(n22392), .S0(n25330), .Y(n4312) );
  XOR2XL U20614 ( .A(n22391), .B(n22390), .Y(n22392) );
  NAND2XL U20615 ( .A(n13097), .B(n22389), .Y(n22390) );
  XOR2XL U20616 ( .A(n22399), .B(n22398), .Y(n22400) );
  NAND2XL U20617 ( .A(n22397), .B(n22396), .Y(n22398) );
  AOI21XL U20618 ( .A0(n22404), .A1(n22402), .B0(n22394), .Y(n22399) );
  MXI2XL U20619 ( .A(U0_pipe5[5]), .B(n22405), .S0(n6888), .Y(n4314) );
  XNOR2XL U20620 ( .A(n22404), .B(n22403), .Y(n22405) );
  NAND2XL U20621 ( .A(n22402), .B(n22401), .Y(n22403) );
  MXI2XL U20622 ( .A(U0_pipe5[4]), .B(n22414), .S0(n6888), .Y(n4315) );
  NAND2XL U20623 ( .A(n22411), .B(n22410), .Y(n22412) );
  MXI2XL U20624 ( .A(U0_pipe5[3]), .B(n22417), .S0(n22620), .Y(n4316) );
  XOR2XL U20625 ( .A(n22416), .B(n22415), .Y(n22417) );
  MXI2XL U20626 ( .A(U0_pipe5[2]), .B(n22420), .S0(n6888), .Y(n4317) );
  MXI2XL U20627 ( .A(U0_pipe5[1]), .B(n22423), .S0(n5920), .Y(n4318) );
  MXI2XL U20628 ( .A(U0_pipe5[0]), .B(n22424), .S0(n5805), .Y(n4319) );
  XOR2X1 U20629 ( .A(n7710), .B(n7708), .Y(n22179) );
  XOR2XL U20630 ( .A(n22197), .B(n22196), .Y(n22198) );
  XOR2XL U20631 ( .A(n22208), .B(n22207), .Y(n22209) );
  XOR2XL U20632 ( .A(n22233), .B(n22232), .Y(n22234) );
  AOI21XL U20633 ( .A0(n22236), .A1(n22231), .B0(n22230), .Y(n22233) );
  XNOR2XL U20634 ( .A(n22236), .B(n22235), .Y(n22237) );
  XOR2XL U20635 ( .A(n22244), .B(n22243), .Y(n22245) );
  XNOR2XL U20636 ( .A(n22247), .B(n22246), .Y(n22249) );
  XOR2XL U20637 ( .A(n22256), .B(n22255), .Y(n22257) );
  AOI21XL U20638 ( .A0(n22259), .A1(n22254), .B0(n22253), .Y(n22256) );
  INVXL U20639 ( .A(n22252), .Y(n22253) );
  XNOR2XL U20640 ( .A(n22259), .B(n22258), .Y(n22260) );
  XOR2XL U20641 ( .A(n22262), .B(n22261), .Y(n22263) );
  XOR2XL U20642 ( .A(n22268), .B(n22267), .Y(n22269) );
  XOR2XL U20643 ( .A(n22274), .B(n22273), .Y(n22275) );
  AOI21XL U20644 ( .A0(n22277), .A1(n22272), .B0(n22271), .Y(n22274) );
  INVXL U20645 ( .A(n22270), .Y(n22271) );
  MXI2XL U20646 ( .A(U0_pipe4[5]), .B(n22278), .S0(n22248), .Y(n4342) );
  XNOR2XL U20647 ( .A(n22277), .B(n22276), .Y(n22278) );
  MXI2XL U20648 ( .A(U0_pipe4[4]), .B(n22284), .S0(n22248), .Y(n4343) );
  XNOR2XL U20649 ( .A(n22283), .B(n22282), .Y(n22284) );
  MXI2XL U20650 ( .A(U0_pipe4[3]), .B(n22287), .S0(n22248), .Y(n4344) );
  XOR2XL U20651 ( .A(n22286), .B(n22285), .Y(n22287) );
  MXI2XL U20652 ( .A(U0_pipe4[2]), .B(n22290), .S0(n22248), .Y(n4345) );
  MXI2XL U20653 ( .A(U0_pipe4[1]), .B(n22293), .S0(n22248), .Y(n4346) );
  MXI2XL U20654 ( .A(U0_pipe4[0]), .B(n22294), .S0(n22248), .Y(n4347) );
  XOR2X1 U20655 ( .A(n24727), .B(n24726), .Y(n24728) );
  NAND2XL U20656 ( .A(n6984), .B(n24767), .Y(n24768) );
  NAND2XL U20657 ( .A(n24648), .B(n24771), .Y(n24772) );
  INVXL U20658 ( .A(n25052), .Y(n24782) );
  AOI21XL U20659 ( .A0(n24788), .A1(n24779), .B0(n24778), .Y(n24783) );
  INVXL U20660 ( .A(n25055), .Y(n24787) );
  INVXL U20661 ( .A(n25063), .Y(n24799) );
  AOI21XL U20662 ( .A0(n24804), .A1(n24795), .B0(n24794), .Y(n24800) );
  INVXL U20663 ( .A(n25066), .Y(n24803) );
  XOR2XL U20664 ( .A(n24808), .B(n24807), .Y(n24809) );
  INVXL U20665 ( .A(n25069), .Y(n24807) );
  XOR2XL U20666 ( .A(n24815), .B(n24814), .Y(n24816) );
  NAND2XL U20667 ( .A(n24585), .B(n24813), .Y(n24814) );
  AOI21XL U20668 ( .A0(n24828), .A1(n24812), .B0(n24811), .Y(n24815) );
  NAND2XL U20669 ( .A(n24821), .B(n24820), .Y(n24822) );
  AOI21XL U20670 ( .A0(n24828), .A1(n24826), .B0(n24818), .Y(n24823) );
  XNOR2XL U20671 ( .A(n24828), .B(n24827), .Y(n24829) );
  NAND2XL U20672 ( .A(n24826), .B(n24825), .Y(n24827) );
  MXI2XL U20673 ( .A(U0_pipe3[4]), .B(n24838), .S0(n24784), .Y(n4371) );
  XNOR2XL U20674 ( .A(n24837), .B(n24836), .Y(n24838) );
  NAND2XL U20675 ( .A(n24835), .B(n24834), .Y(n24836) );
  MXI2XL U20676 ( .A(U0_pipe3[3]), .B(n24842), .S0(n24784), .Y(n4372) );
  XOR2XL U20677 ( .A(n24841), .B(n24840), .Y(n24842) );
  INVXL U20678 ( .A(n25103), .Y(n24840) );
  MXI2XL U20679 ( .A(U0_pipe3[2]), .B(n24846), .S0(n24784), .Y(n4373) );
  INVXL U20680 ( .A(n25108), .Y(n24845) );
  MXI2XL U20681 ( .A(U0_pipe3[1]), .B(n24850), .S0(n24784), .Y(n4374) );
  INVXL U20682 ( .A(n25112), .Y(n24849) );
  MXI2XL U20683 ( .A(U0_pipe3[0]), .B(n25114), .S0(n24784), .Y(n4375) );
  NAND2XL U20684 ( .A(n24418), .B(n24417), .Y(n24419) );
  INVXL U20685 ( .A(n24870), .Y(n24427) );
  INVXL U20686 ( .A(n24876), .Y(n24436) );
  OAI21XL U20687 ( .A0(n24447), .A1(n24433), .B0(n24432), .Y(n24437) );
  INVXL U20688 ( .A(n24881), .Y(n24442) );
  INVXL U20689 ( .A(n24884), .Y(n24446) );
  INVXL U20690 ( .A(n24456), .Y(n24457) );
  AOI21XL U20691 ( .A0(n24463), .A1(n24455), .B0(n24454), .Y(n24458) );
  INVXL U20692 ( .A(n24887), .Y(n24462) );
  INVXL U20693 ( .A(n24893), .Y(n24470) );
  INVXL U20694 ( .A(n24896), .Y(n24474) );
  INVXL U20695 ( .A(n24905), .Y(n24485) );
  XOR2XL U20696 ( .A(n24490), .B(n24489), .Y(n24491) );
  INVXL U20697 ( .A(n24908), .Y(n24489) );
  XOR2XL U20698 ( .A(n24497), .B(n24496), .Y(n24498) );
  INVXL U20699 ( .A(n24913), .Y(n24496) );
  XNOR2XL U20700 ( .A(n24501), .B(n24500), .Y(n24502) );
  INVXL U20701 ( .A(n24916), .Y(n24500) );
  INVXL U20702 ( .A(n24923), .Y(n24510) );
  INVXL U20703 ( .A(n24926), .Y(n24514) );
  INVXL U20704 ( .A(n24934), .Y(n24526) );
  AOI21XL U20705 ( .A0(n24531), .A1(n24522), .B0(n24521), .Y(n24527) );
  XNOR2XL U20706 ( .A(n24531), .B(n24530), .Y(n24532) );
  INVXL U20707 ( .A(n24937), .Y(n24530) );
  XOR2XL U20708 ( .A(n24535), .B(n24534), .Y(n24536) );
  INVXL U20709 ( .A(n24940), .Y(n24534) );
  XOR2XL U20710 ( .A(n24543), .B(n24542), .Y(n24544) );
  NAND2XL U20711 ( .A(n24541), .B(n24540), .Y(n24542) );
  XOR2XL U20712 ( .A(n24551), .B(n24550), .Y(n24552) );
  NAND2XL U20713 ( .A(n24549), .B(n24548), .Y(n24550) );
  AOI21XL U20714 ( .A0(n24556), .A1(n24554), .B0(n24546), .Y(n24551) );
  MXI2XL U20715 ( .A(U0_pipe2[5]), .B(n24557), .S0(n22853), .Y(n4398) );
  NAND2XL U20716 ( .A(n24554), .B(n24553), .Y(n24555) );
  MXI2XL U20717 ( .A(U0_pipe2[4]), .B(n24564), .S0(n22620), .Y(n4399) );
  XNOR2XL U20718 ( .A(n24563), .B(n24562), .Y(n24564) );
  NAND2XL U20719 ( .A(n24561), .B(n24560), .Y(n24562) );
  MXI2XL U20720 ( .A(U0_pipe2[3]), .B(n24570), .S0(n6888), .Y(n4400) );
  XOR2XL U20721 ( .A(n24569), .B(n24568), .Y(n24570) );
  NAND2XL U20722 ( .A(n24567), .B(n24566), .Y(n24568) );
  INVXL U20723 ( .A(n24565), .Y(n24567) );
  MXI2XL U20724 ( .A(U0_pipe2[2]), .B(n24576), .S0(n6888), .Y(n4401) );
  NAND2XL U20725 ( .A(n24573), .B(n24572), .Y(n24575) );
  INVXL U20726 ( .A(n24571), .Y(n24573) );
  MXI2XL U20727 ( .A(U0_pipe2[1]), .B(n24580), .S0(n6888), .Y(n4402) );
  INVXL U20728 ( .A(n24984), .Y(n24579) );
  MXI2XL U20729 ( .A(U0_pipe2[0]), .B(n24986), .S0(n6888), .Y(n4403) );
  MXI2XL U20730 ( .A(U0_pipe0[2]), .B(n24982), .S0(n5920), .Y(n4408) );
  NAND2XL U20731 ( .A(n24979), .B(n24978), .Y(n24981) );
  INVXL U20732 ( .A(n24977), .Y(n24979) );
  MXI2XL U20733 ( .A(U0_pipe8[22]), .B(n25546), .S0(n5810), .Y(n4412) );
  XOR2XL U20734 ( .A(n25548), .B(n25547), .Y(n25549) );
  XNOR2X1 U20735 ( .A(n25560), .B(n25559), .Y(n25561) );
  XOR2X1 U20736 ( .A(n25563), .B(n25562), .Y(n25564) );
  XNOR2X1 U20737 ( .A(n25572), .B(n25571), .Y(n25573) );
  XOR2XL U20738 ( .A(n25584), .B(n25583), .Y(n25585) );
  XOR2XL U20739 ( .A(n25589), .B(n25588), .Y(n25590) );
  AOI21XL U20740 ( .A0(n25592), .A1(n25587), .B0(n25586), .Y(n25589) );
  XNOR2XL U20741 ( .A(n25592), .B(n25591), .Y(n25593) );
  XOR2XL U20742 ( .A(n25599), .B(n25598), .Y(n25600) );
  XNOR2XL U20743 ( .A(n25602), .B(n25601), .Y(n25603) );
  XOR2XL U20744 ( .A(n25610), .B(n25609), .Y(n25612) );
  AOI21XL U20745 ( .A0(n25614), .A1(n25608), .B0(n25607), .Y(n25610) );
  INVXL U20746 ( .A(n25606), .Y(n25607) );
  XOR2XL U20747 ( .A(n25623), .B(n25622), .Y(n25624) );
  XOR2XL U20748 ( .A(n25629), .B(n25628), .Y(n25630) );
  AOI21XL U20749 ( .A0(n25632), .A1(n25627), .B0(n25626), .Y(n25629) );
  INVXL U20750 ( .A(n25625), .Y(n25626) );
  MXI2XL U20751 ( .A(U0_pipe8[5]), .B(n25633), .S0(n6888), .Y(n4429) );
  XNOR2XL U20752 ( .A(n25632), .B(n25631), .Y(n25633) );
  MXI2XL U20753 ( .A(U0_pipe8[4]), .B(n25639), .S0(n6888), .Y(n4430) );
  XNOR2XL U20754 ( .A(n25638), .B(n25637), .Y(n25639) );
  MXI2XL U20755 ( .A(U0_pipe8[3]), .B(n25642), .S0(n6888), .Y(n4431) );
  XOR2XL U20756 ( .A(n25641), .B(n25640), .Y(n25642) );
  MXI2XL U20757 ( .A(U0_pipe8[2]), .B(n25645), .S0(n6888), .Y(n4432) );
  MXI2XL U20758 ( .A(U0_pipe8[1]), .B(n25648), .S0(n6888), .Y(n4433) );
  MXI2XL U20759 ( .A(U0_pipe8[0]), .B(n25649), .S0(n6888), .Y(n4434) );
  XOR2X1 U20760 ( .A(n21946), .B(n25286), .Y(n7731) );
  INVXL U20761 ( .A(n22306), .Y(n21964) );
  INVXL U20762 ( .A(n22311), .Y(n21970) );
  INVXL U20763 ( .A(n22314), .Y(n21975) );
  INVXL U20764 ( .A(n22326), .Y(n21987) );
  XOR2X1 U20765 ( .A(n21994), .B(n21993), .Y(n21995) );
  INVXL U20766 ( .A(n22332), .Y(n21993) );
  XNOR2X1 U20767 ( .A(n21998), .B(n21997), .Y(n21999) );
  INVXL U20768 ( .A(n22335), .Y(n21997) );
  NAND2XL U20769 ( .A(n7016), .B(n22005), .Y(n22006) );
  NAND2XL U20770 ( .A(n22016), .B(n22015), .Y(n22017) );
  XNOR2X1 U20771 ( .A(n22022), .B(n22021), .Y(n22023) );
  INVXL U20772 ( .A(n22366), .Y(n22031) );
  AOI21XL U20773 ( .A0(n22036), .A1(n22028), .B0(n22027), .Y(n22032) );
  INVXL U20774 ( .A(n22369), .Y(n22035) );
  INVXL U20775 ( .A(n22377), .Y(n22047) );
  AOI21XL U20776 ( .A0(n22052), .A1(n22043), .B0(n22042), .Y(n22048) );
  INVXL U20777 ( .A(n22380), .Y(n22051) );
  XOR2XL U20778 ( .A(n22056), .B(n22055), .Y(n22057) );
  INVXL U20779 ( .A(n22383), .Y(n22055) );
  XOR2XL U20780 ( .A(n22063), .B(n22062), .Y(n22064) );
  NAND2XL U20781 ( .A(n14514), .B(n22061), .Y(n22062) );
  XOR2XL U20782 ( .A(n22071), .B(n22070), .Y(n22072) );
  NAND2XL U20783 ( .A(n22069), .B(n22068), .Y(n22070) );
  AOI21XL U20784 ( .A0(n22076), .A1(n22074), .B0(n22066), .Y(n22071) );
  XNOR2XL U20785 ( .A(n22076), .B(n22075), .Y(n22077) );
  MXI2XL U20786 ( .A(U0_pipe7[4]), .B(n22086), .S0(n21972), .Y(n4458) );
  NAND2XL U20787 ( .A(n22083), .B(n22082), .Y(n22084) );
  MXI2XL U20788 ( .A(U0_pipe7[3]), .B(n22090), .S0(n21972), .Y(n4459) );
  XOR2XL U20789 ( .A(n22089), .B(n22088), .Y(n22090) );
  INVXL U20790 ( .A(n22415), .Y(n22088) );
  MXI2XL U20791 ( .A(U0_pipe7[2]), .B(n22096), .S0(n21972), .Y(n4460) );
  INVXL U20792 ( .A(n22419), .Y(n22095) );
  MXI2XL U20793 ( .A(U0_pipe7[1]), .B(n22100), .S0(n21972), .Y(n4461) );
  INVXL U20794 ( .A(n22422), .Y(n22099) );
  MXI2XL U20795 ( .A(U0_pipe7[0]), .B(n22424), .S0(n21972), .Y(n4462) );
  INVXL U20796 ( .A(n22181), .Y(n21812) );
  INVXL U20797 ( .A(n22183), .Y(n21819) );
  INVXL U20798 ( .A(n22188), .Y(n21827) );
  INVXL U20799 ( .A(n22193), .Y(n21833) );
  INVXL U20800 ( .A(n22196), .Y(n21836) );
  XNOR2X1 U20801 ( .A(n21849), .B(n21848), .Y(n21850) );
  INVXL U20802 ( .A(n22207), .Y(n21848) );
  INVXL U20803 ( .A(n22213), .Y(n21854) );
  INVXL U20804 ( .A(n22216), .Y(n21857) );
  INVXL U20805 ( .A(n22224), .Y(n21867) );
  XOR2XL U20806 ( .A(n21871), .B(n21870), .Y(n21872) );
  INVXL U20807 ( .A(n22227), .Y(n21870) );
  XOR2XL U20808 ( .A(n21876), .B(n21875), .Y(n21877) );
  INVXL U20809 ( .A(n22232), .Y(n21875) );
  INVXL U20810 ( .A(n22235), .Y(n21878) );
  INVXL U20811 ( .A(n22243), .Y(n21887) );
  AOI21XL U20812 ( .A0(n21892), .A1(n21885), .B0(n21884), .Y(n21888) );
  INVXL U20813 ( .A(n22246), .Y(n21891) );
  INVXL U20814 ( .A(n22255), .Y(n21901) );
  AOI21XL U20815 ( .A0(n21905), .A1(n21899), .B0(n21898), .Y(n21902) );
  INVXL U20816 ( .A(n22258), .Y(n21904) );
  XOR2XL U20817 ( .A(n21908), .B(n21907), .Y(n21909) );
  INVXL U20818 ( .A(n22261), .Y(n21907) );
  XOR2XL U20819 ( .A(n21914), .B(n21913), .Y(n21915) );
  INVXL U20820 ( .A(n22267), .Y(n21913) );
  XOR2XL U20821 ( .A(n21922), .B(n21921), .Y(n21923) );
  INVXL U20822 ( .A(n22273), .Y(n21921) );
  AOI21XL U20823 ( .A0(n21925), .A1(n21919), .B0(n21918), .Y(n21922) );
  XNOR2XL U20824 ( .A(n21925), .B(n21924), .Y(n21926) );
  INVXL U20825 ( .A(n22276), .Y(n21924) );
  MXI2XL U20826 ( .A(U0_pipe6[4]), .B(n21933), .S0(n21972), .Y(n4486) );
  XNOR2XL U20827 ( .A(n21932), .B(n21931), .Y(n21933) );
  INVXL U20828 ( .A(n22282), .Y(n21931) );
  MXI2XL U20829 ( .A(U0_pipe6[3]), .B(n21937), .S0(n21972), .Y(n4487) );
  INVXL U20830 ( .A(n22285), .Y(n21935) );
  MXI2XL U20831 ( .A(U0_pipe6[2]), .B(n21941), .S0(n21972), .Y(n4488) );
  INVXL U20832 ( .A(n22289), .Y(n21940) );
  MXI2XL U20833 ( .A(U0_pipe6[1]), .B(n21945), .S0(n22248), .Y(n4489) );
  INVXL U20834 ( .A(n22292), .Y(n21944) );
  MXI2XL U20835 ( .A(U0_pipe6[0]), .B(n22294), .S0(n22248), .Y(n4490) );
  XOR2XL U20836 ( .A(n22315), .B(n22314), .Y(n22316) );
  XOR2XL U20837 ( .A(n22327), .B(n22326), .Y(n22328) );
  XOR2XL U20838 ( .A(n22331), .B(n22335), .Y(n22336) );
  XOR2XL U20839 ( .A(n22349), .B(n22348), .Y(n22350) );
  NAND2XL U20840 ( .A(n22353), .B(n22352), .Y(n22354) );
  XNOR2X1 U20841 ( .A(n22359), .B(n22358), .Y(n22360) );
  XOR2XL U20842 ( .A(n22367), .B(n22366), .Y(n22368) );
  XNOR2XL U20843 ( .A(n22370), .B(n22369), .Y(n22371) );
  MXI2XL U20844 ( .A(U0_pipe0[1]), .B(n24985), .S0(n25101), .Y(n4508) );
  INVXL U20845 ( .A(n25598), .Y(n25213) );
  INVXL U20846 ( .A(n25601), .Y(n25217) );
  INVXL U20847 ( .A(n25609), .Y(n25228) );
  AOI21XL U20848 ( .A0(n25233), .A1(n25225), .B0(n25224), .Y(n25229) );
  INVXL U20849 ( .A(n25613), .Y(n25232) );
  MXI2XL U20850 ( .A(U0_pipe12[8]), .B(n25238), .S0(n5810), .Y(n4513) );
  XOR2XL U20851 ( .A(n25237), .B(n25236), .Y(n25238) );
  INVXL U20852 ( .A(n25616), .Y(n25236) );
  MXI2XL U20853 ( .A(U0_pipe12[7]), .B(n25246), .S0(n5810), .Y(n4514) );
  XOR2XL U20854 ( .A(n25245), .B(n25244), .Y(n25246) );
  INVXL U20855 ( .A(n25622), .Y(n25244) );
  MXI2XL U20856 ( .A(U0_pipe12[6]), .B(n25255), .S0(n5810), .Y(n4515) );
  XOR2XL U20857 ( .A(n25254), .B(n25253), .Y(n25255) );
  INVXL U20858 ( .A(n25628), .Y(n25253) );
  AOI21XL U20859 ( .A0(n25258), .A1(n25250), .B0(n25249), .Y(n25254) );
  INVXL U20860 ( .A(n25631), .Y(n25257) );
  MXI2XL U20861 ( .A(U0_pipe12[4]), .B(n25268), .S0(n25267), .Y(n4517) );
  XNOR2XL U20862 ( .A(n25266), .B(n25265), .Y(n25268) );
  INVXL U20863 ( .A(n25637), .Y(n25265) );
  MXI2XL U20864 ( .A(U0_pipe12[3]), .B(n25274), .S0(n25273), .Y(n4518) );
  XOR2XL U20865 ( .A(n25272), .B(n25271), .Y(n25274) );
  INVXL U20866 ( .A(n25640), .Y(n25271) );
  MXI2XL U20867 ( .A(U0_pipe12[2]), .B(n25279), .S0(n25318), .Y(n4519) );
  INVXL U20868 ( .A(n25644), .Y(n25278) );
  MXI2XL U20869 ( .A(U0_pipe12[1]), .B(n25284), .S0(n25318), .Y(n4520) );
  INVXL U20870 ( .A(n25647), .Y(n25283) );
  MXI2XL U20871 ( .A(U0_pipe12[0]), .B(n25649), .S0(n25318), .Y(n4521) );
  NAND2XL U20872 ( .A(n22986), .B(n22985), .Y(n22987) );
  INVXL U20873 ( .A(n22991), .Y(n22992) );
  XOR2X1 U20874 ( .A(n22997), .B(n22996), .Y(n22998) );
  INVXL U20875 ( .A(n22995), .Y(n22996) );
  NAND2XL U20876 ( .A(n23010), .B(n23009), .Y(n23011) );
  NAND2XL U20877 ( .A(n23017), .B(n23016), .Y(n23018) );
  NAND2XL U20878 ( .A(n23022), .B(n23021), .Y(n23023) );
  NAND2XL U20879 ( .A(n23032), .B(n23031), .Y(n23033) );
  NAND2XL U20880 ( .A(n23056), .B(n23055), .Y(n23057) );
  NAND2XL U20881 ( .A(n22919), .B(n23060), .Y(n23061) );
  NAND2XL U20882 ( .A(n23070), .B(n23069), .Y(n23071) );
  AOI21XL U20883 ( .A0(n23077), .A1(n23075), .B0(n23067), .Y(n23072) );
  XOR2XL U20884 ( .A(n23081), .B(n23080), .Y(n23082) );
  INVXL U20885 ( .A(n23079), .Y(n23080) );
  XOR2XL U20886 ( .A(n23089), .B(n23088), .Y(n23090) );
  NAND2XL U20887 ( .A(n23087), .B(n23086), .Y(n23088) );
  XOR2XL U20888 ( .A(n23097), .B(n23096), .Y(n23098) );
  NAND2XL U20889 ( .A(n23095), .B(n23094), .Y(n23096) );
  AOI21XL U20890 ( .A0(n23102), .A1(n23100), .B0(n23092), .Y(n23097) );
  XNOR2XL U20891 ( .A(n23102), .B(n23101), .Y(n23103) );
  NAND2XL U20892 ( .A(n23100), .B(n23099), .Y(n23101) );
  XNOR2XL U20893 ( .A(n23109), .B(n23108), .Y(n23110) );
  INVXL U20894 ( .A(n23107), .Y(n23108) );
  MXI2XL U20895 ( .A(U0_pipe11[3]), .B(n23114), .S0(n24784), .Y(n4546) );
  INVXL U20896 ( .A(n23111), .Y(n23112) );
  MXI2XL U20897 ( .A(U0_pipe11[2]), .B(n23118), .S0(n24784), .Y(n4547) );
  INVXL U20898 ( .A(n23115), .Y(n23117) );
  MXI2XL U20899 ( .A(U0_pipe11[1]), .B(n23122), .S0(n24784), .Y(n4548) );
  INVXL U20900 ( .A(n23119), .Y(n23121) );
  MXI2XL U20901 ( .A(U0_pipe11[0]), .B(n23123), .S0(n24784), .Y(n4549) );
  NAND2XL U20902 ( .A(n22740), .B(n22739), .Y(n22741) );
  INVXL U20903 ( .A(n22738), .Y(n22740) );
  INVXL U20904 ( .A(n22747), .Y(n22748) );
  INVXL U20905 ( .A(n22755), .Y(n22756) );
  INVXL U20906 ( .A(n22761), .Y(n22762) );
  INVXL U20907 ( .A(n22765), .Y(n22766) );
  INVXL U20908 ( .A(n14104), .Y(n14105) );
  XNOR2X1 U20909 ( .A(n22771), .B(n22770), .Y(n22772) );
  INVXL U20910 ( .A(n22769), .Y(n22770) );
  INVXL U20911 ( .A(n22775), .Y(n22776) );
  INVXL U20912 ( .A(n22779), .Y(n22780) );
  INVXL U20913 ( .A(n22789), .Y(n22790) );
  INVXL U20914 ( .A(n22793), .Y(n22794) );
  INVXL U20915 ( .A(n22799), .Y(n22800) );
  XNOR2X1 U20916 ( .A(n22805), .B(n22804), .Y(n22806) );
  INVXL U20917 ( .A(n22803), .Y(n22804) );
  INVXL U20918 ( .A(n22812), .Y(n22813) );
  XNOR2XL U20919 ( .A(n22818), .B(n22817), .Y(n22819) );
  INVXL U20920 ( .A(n22816), .Y(n22817) );
  INVXL U20921 ( .A(n22826), .Y(n22827) );
  AOI21XL U20922 ( .A0(n22832), .A1(n22825), .B0(n22824), .Y(n22828) );
  XNOR2XL U20923 ( .A(n22832), .B(n22831), .Y(n22833) );
  INVXL U20924 ( .A(n22830), .Y(n22831) );
  XOR2XL U20925 ( .A(n22836), .B(n22835), .Y(n22837) );
  INVXL U20926 ( .A(n22834), .Y(n22835) );
  XOR2XL U20927 ( .A(n22844), .B(n22843), .Y(n22845) );
  NAND2XL U20928 ( .A(n22842), .B(n22841), .Y(n22843) );
  MXI2XL U20929 ( .A(U0_pipe10[6]), .B(n22854), .S0(n5805), .Y(n4571) );
  XOR2XL U20930 ( .A(n22852), .B(n22851), .Y(n22854) );
  NAND2XL U20931 ( .A(n22850), .B(n22849), .Y(n22851) );
  AOI21XL U20932 ( .A0(n22858), .A1(n22856), .B0(n22847), .Y(n22852) );
  MXI2XL U20933 ( .A(U0_pipe10[5]), .B(n22859), .S0(n5805), .Y(n4572) );
  XNOR2XL U20934 ( .A(n22858), .B(n22857), .Y(n22859) );
  NAND2XL U20935 ( .A(n22856), .B(n22855), .Y(n22857) );
  MXI2XL U20936 ( .A(U0_pipe10[4]), .B(n22866), .S0(n5805), .Y(n4573) );
  XNOR2XL U20937 ( .A(n22865), .B(n22864), .Y(n22866) );
  NAND2XL U20938 ( .A(n22863), .B(n22862), .Y(n22864) );
  MXI2XL U20939 ( .A(U0_pipe10[3]), .B(n22872), .S0(n5805), .Y(n4574) );
  XOR2XL U20940 ( .A(n22871), .B(n22870), .Y(n22872) );
  NAND2XL U20941 ( .A(n22869), .B(n22868), .Y(n22870) );
  INVXL U20942 ( .A(n22867), .Y(n22869) );
  MXI2XL U20943 ( .A(U0_pipe10[2]), .B(n22878), .S0(n5805), .Y(n4575) );
  NAND2XL U20944 ( .A(n22875), .B(n22874), .Y(n22877) );
  INVXL U20945 ( .A(n22873), .Y(n22875) );
  MXI2XL U20946 ( .A(U0_pipe10[1]), .B(n22882), .S0(n24784), .Y(n4576) );
  INVXL U20947 ( .A(n22879), .Y(n22881) );
  MXI2XL U20948 ( .A(U0_pipe10[0]), .B(n22883), .S0(n24784), .Y(n4577) );
  MXI2XL U20949 ( .A(U0_pipe9[21]), .B(n25676), .S0(n25330), .Y(n4584) );
  XOR2X1 U20950 ( .A(n25689), .B(n25688), .Y(n25690) );
  XOR2XL U20951 ( .A(n25693), .B(n25697), .Y(n25698) );
  XOR2XL U20952 ( .A(n25712), .B(n25711), .Y(n25713) );
  NAND2XL U20953 ( .A(n25728), .B(n25727), .Y(n25729) );
  NAND2XL U20954 ( .A(n25743), .B(n25742), .Y(n25744) );
  XOR2XL U20955 ( .A(n25753), .B(n25752), .Y(n25754) );
  XOR2XL U20956 ( .A(n25760), .B(n25759), .Y(n25761) );
  NAND2XL U20957 ( .A(n12087), .B(n25758), .Y(n25759) );
  XOR2XL U20958 ( .A(n25768), .B(n25767), .Y(n25769) );
  NAND2XL U20959 ( .A(n25766), .B(n25765), .Y(n25767) );
  AOI21XL U20960 ( .A0(n25773), .A1(n25771), .B0(n25763), .Y(n25768) );
  XNOR2XL U20961 ( .A(n25773), .B(n25772), .Y(n25774) );
  NAND2XL U20962 ( .A(n25771), .B(n25770), .Y(n25772) );
  MXI2XL U20963 ( .A(U0_pipe9[4]), .B(n25780), .S0(n6887), .Y(n4601) );
  XNOR2XL U20964 ( .A(n25779), .B(n25778), .Y(n25780) );
  MXI2XL U20965 ( .A(U0_pipe9[3]), .B(n25783), .S0(n6887), .Y(n4602) );
  XOR2XL U20966 ( .A(n25782), .B(n25781), .Y(n25783) );
  MXI2XL U20967 ( .A(U0_pipe9[2]), .B(n25786), .S0(n6887), .Y(n4603) );
  MXI2XL U20968 ( .A(U0_pipe9[1]), .B(n25790), .S0(n6887), .Y(n4604) );
  NAND2XL U20969 ( .A(n12118), .B(n25787), .Y(n25789) );
  MXI2XL U20970 ( .A(U0_pipe9[0]), .B(n25791), .S0(n6887), .Y(n4605) );
  XOR2X1 U20971 ( .A(n25528), .B(U2_A_r_d[25]), .Y(n7597) );
  MXI2XL U20972 ( .A(U0_pipe0[0]), .B(n24986), .S0(n25101), .Y(n4608) );
  XOR2X1 U20973 ( .A(n22614), .B(n22995), .Y(n22615) );
  MXI2XL U20974 ( .A(U0_pipe15[17]), .B(n22631), .S0(n25330), .Y(n4619) );
  AOI21XL U20975 ( .A0(n22655), .A1(n12612), .B0(n22647), .Y(n22651) );
  AOI21XL U20976 ( .A0(n22681), .A1(n22679), .B0(n22671), .Y(n22676) );
  XOR2XL U20977 ( .A(n22685), .B(n23079), .Y(n22686) );
  XOR2XL U20978 ( .A(n22692), .B(n22691), .Y(n22693) );
  NAND2BXL U20979 ( .AN(n12481), .B(n22690), .Y(n22691) );
  XOR2XL U20980 ( .A(n22700), .B(n22699), .Y(n22701) );
  NAND2XL U20981 ( .A(n22698), .B(n22697), .Y(n22699) );
  AOI21XL U20982 ( .A0(n22705), .A1(n22703), .B0(n22695), .Y(n22700) );
  XNOR2XL U20983 ( .A(n22705), .B(n22704), .Y(n22706) );
  NAND2XL U20984 ( .A(n22703), .B(n22702), .Y(n22704) );
  MXI2XL U20985 ( .A(U0_pipe15[4]), .B(n22712), .S0(n25330), .Y(n4632) );
  XNOR2XL U20986 ( .A(n22711), .B(n23107), .Y(n22712) );
  MXI2XL U20987 ( .A(U0_pipe15[3]), .B(n22717), .S0(n6887), .Y(n4633) );
  XOR2XL U20988 ( .A(n22716), .B(n23111), .Y(n22717) );
  MXI2XL U20989 ( .A(U0_pipe15[2]), .B(n22722), .S0(n22620), .Y(n4634) );
  XNOR2XL U20990 ( .A(n22721), .B(n23115), .Y(n22722) );
  MXI2XL U20991 ( .A(U0_pipe15[1]), .B(n22726), .S0(n22620), .Y(n4635) );
  MXI2XL U20992 ( .A(U0_pipe15[0]), .B(n23123), .S0(n25330), .Y(n4636) );
  NAND2XL U20993 ( .A(n22464), .B(n22463), .Y(n22465) );
  OAI21XL U20994 ( .A0(n22490), .A1(n22432), .B0(n22488), .Y(n14054) );
  XOR2XL U20995 ( .A(n22490), .B(n22769), .Y(n22491) );
  NAND2XL U20996 ( .A(n7574), .B(n22497), .Y(n22495) );
  XNOR2XL U20997 ( .A(n22498), .B(n22779), .Y(n22499) );
  XOR2XL U20998 ( .A(n22511), .B(n22793), .Y(n22512) );
  XOR2XL U20999 ( .A(n22516), .B(n22799), .Y(n22517) );
  AOI21XL U21000 ( .A0(n5854), .A1(n22519), .B0(n22513), .Y(n22516) );
  XNOR2XL U21001 ( .A(n5854), .B(n22803), .Y(n22520) );
  XNOR2XL U21002 ( .A(n22530), .B(n22816), .Y(n22531) );
  XOR2XL U21003 ( .A(n22538), .B(n22826), .Y(n22539) );
  INVXL U21004 ( .A(n22540), .Y(n22534) );
  MXI2XL U21005 ( .A(U0_pipe14[8]), .B(n22548), .S0(n5805), .Y(n4656) );
  XOR2XL U21006 ( .A(n22547), .B(n22834), .Y(n22548) );
  MXI2XL U21007 ( .A(U0_pipe14[7]), .B(n22555), .S0(n5805), .Y(n4657) );
  XOR2XL U21008 ( .A(n22554), .B(n22553), .Y(n22555) );
  NAND2XL U21009 ( .A(n14015), .B(n22552), .Y(n22553) );
  MXI2XL U21010 ( .A(U0_pipe14[6]), .B(n22563), .S0(n5805), .Y(n4658) );
  XOR2XL U21011 ( .A(n22562), .B(n22561), .Y(n22563) );
  NAND2XL U21012 ( .A(n22560), .B(n22559), .Y(n22561) );
  AOI21XL U21013 ( .A0(n22567), .A1(n22565), .B0(n22557), .Y(n22562) );
  MXI2XL U21014 ( .A(U0_pipe14[5]), .B(n22568), .S0(n5805), .Y(n4659) );
  XNOR2XL U21015 ( .A(n22567), .B(n22566), .Y(n22568) );
  NAND2XL U21016 ( .A(n22565), .B(n22564), .Y(n22566) );
  MXI2XL U21017 ( .A(U0_pipe14[4]), .B(n22575), .S0(n5805), .Y(n4660) );
  XNOR2XL U21018 ( .A(n22574), .B(n22573), .Y(n22575) );
  NAND2XL U21019 ( .A(n22572), .B(n22571), .Y(n22573) );
  MXI2XL U21020 ( .A(U0_pipe14[3]), .B(n22581), .S0(n5805), .Y(n4661) );
  XOR2XL U21021 ( .A(n22580), .B(n22579), .Y(n22581) );
  NAND2XL U21022 ( .A(n22578), .B(n22577), .Y(n22579) );
  INVXL U21023 ( .A(n22576), .Y(n22578) );
  MXI2XL U21024 ( .A(U0_pipe14[2]), .B(n22587), .S0(n22620), .Y(n4662) );
  NAND2XL U21025 ( .A(n22584), .B(n22583), .Y(n22586) );
  INVXL U21026 ( .A(n22582), .Y(n22584) );
  MXI2XL U21027 ( .A(U0_pipe14[1]), .B(n22590), .S0(n22620), .Y(n4663) );
  MXI2XL U21028 ( .A(U0_pipe14[0]), .B(n22883), .S0(n22620), .Y(n4664) );
  XOR2X1 U21029 ( .A(n25317), .B(n25316), .Y(n25319) );
  INVXL U21030 ( .A(n25674), .Y(n25316) );
  INVXL U21031 ( .A(n25688), .Y(n25333) );
  INVXL U21032 ( .A(n25697), .Y(n25344) );
  NAND2XL U21033 ( .A(n25364), .B(n25363), .Y(n25365) );
  MXI2XL U21034 ( .A(U0_pipe13[13]), .B(n25371), .S0(n25330), .Y(n4679) );
  NAND2XL U21035 ( .A(n25377), .B(n25376), .Y(n25378) );
  NAND2XL U21036 ( .A(n25391), .B(n25390), .Y(n25392) );
  MXI2XL U21037 ( .A(U0_pipe13[9]), .B(n25399), .S0(U1_valid[0]), .Y(n4683) );
  NAND2XL U21038 ( .A(n25396), .B(n25395), .Y(n25397) );
  XOR2XL U21039 ( .A(n25402), .B(n25401), .Y(n25403) );
  INVXL U21040 ( .A(n25752), .Y(n25401) );
  XOR2XL U21041 ( .A(n25409), .B(n25408), .Y(n25410) );
  NAND2XL U21042 ( .A(n12362), .B(n25407), .Y(n25408) );
  AOI21XL U21043 ( .A0(n25422), .A1(n25406), .B0(n25405), .Y(n25409) );
  XOR2XL U21044 ( .A(n25417), .B(n25416), .Y(n25418) );
  NAND2XL U21045 ( .A(n25415), .B(n25414), .Y(n25416) );
  XNOR2XL U21046 ( .A(n25422), .B(n25421), .Y(n25423) );
  NAND2XL U21047 ( .A(n25420), .B(n25419), .Y(n25421) );
  MXI2XL U21048 ( .A(U0_pipe13[4]), .B(n25432), .S0(n6887), .Y(n4688) );
  XNOR2XL U21049 ( .A(n25431), .B(n25430), .Y(n25432) );
  INVXL U21050 ( .A(n25778), .Y(n25430) );
  MXI2XL U21051 ( .A(U0_pipe13[3]), .B(n25436), .S0(n6887), .Y(n4689) );
  XOR2XL U21052 ( .A(n25435), .B(n25434), .Y(n25436) );
  INVXL U21053 ( .A(n25781), .Y(n25434) );
  MXI2XL U21054 ( .A(U0_pipe13[2]), .B(n25442), .S0(n6887), .Y(n4690) );
  INVXL U21055 ( .A(n25785), .Y(n25441) );
  MXI2XL U21056 ( .A(U0_pipe13[1]), .B(n25447), .S0(n6887), .Y(n4691) );
  NAND2XL U21057 ( .A(n25444), .B(n25443), .Y(n25446) );
  MXI2XL U21058 ( .A(U0_pipe13[0]), .B(n25791), .S0(n6887), .Y(n4692) );
  MXI2XL U21059 ( .A(U0_pipe12[25]), .B(n25128), .S0(n5810), .Y(n4695) );
  INVXL U21060 ( .A(n25530), .Y(n25126) );
  INVXL U21061 ( .A(n25539), .Y(n25142) );
  INVXL U21062 ( .A(n25544), .Y(n25148) );
  MXI2XL U21063 ( .A(U0_pipe12[21]), .B(n25154), .S0(n5810), .Y(n4699) );
  INVXL U21064 ( .A(n25547), .Y(n25152) );
  INVXL U21065 ( .A(n25559), .Y(n25163) );
  MXI2XL U21066 ( .A(U0_pipe12[19]), .B(n25169), .S0(n5810), .Y(n4701) );
  XNOR2X1 U21067 ( .A(n25168), .B(n25167), .Y(n25169) );
  INVXL U21068 ( .A(n25562), .Y(n25167) );
  INVXL U21069 ( .A(n25568), .Y(n25175) );
  INVXL U21070 ( .A(n25571), .Y(n25179) );
  INVXL U21071 ( .A(n25580), .Y(n25190) );
  XOR2XL U21072 ( .A(n25195), .B(n25194), .Y(n25196) );
  INVXL U21073 ( .A(n25583), .Y(n25194) );
  XOR2XL U21074 ( .A(n25201), .B(n25200), .Y(n25202) );
  INVXL U21075 ( .A(n25588), .Y(n25200) );
  INVXL U21076 ( .A(n25591), .Y(n25204) );
  MXI2XL U21077 ( .A(U1_pipe12[13]), .B(n19871), .S0(n25330), .Y(n4708) );
  XNOR2XL U21078 ( .A(n19870), .B(n19869), .Y(n19871) );
  INVXL U21079 ( .A(n20250), .Y(n19869) );
  MXI2XL U21080 ( .A(U1_pipe12[14]), .B(n19867), .S0(n25330), .Y(n4709) );
  XOR2XL U21081 ( .A(n19866), .B(n19865), .Y(n19867) );
  INVXL U21082 ( .A(n20247), .Y(n19865) );
  MXI2XL U21083 ( .A(U1_pipe12[15]), .B(n19861), .S0(n25330), .Y(n4710) );
  XOR2XL U21084 ( .A(n19860), .B(n19859), .Y(n19861) );
  INVXL U21085 ( .A(n20242), .Y(n19859) );
  MXI2XL U21086 ( .A(U1_pipe12[16]), .B(n19857), .S0(n25330), .Y(n4711) );
  INVXL U21087 ( .A(n20238), .Y(n19855) );
  MXI2XL U21088 ( .A(U1_pipe12[17]), .B(n19846), .S0(n25330), .Y(n4712) );
  XNOR2XL U21089 ( .A(n19845), .B(n19844), .Y(n19846) );
  INVXL U21090 ( .A(n20229), .Y(n19844) );
  MXI2XL U21091 ( .A(U1_pipe12[18]), .B(n19842), .S0(n25330), .Y(n4713) );
  XOR2XL U21092 ( .A(n19841), .B(n19840), .Y(n19842) );
  INVXL U21093 ( .A(n20226), .Y(n19840) );
  MXI2XL U21094 ( .A(U1_pipe12[19]), .B(n19834), .S0(n25330), .Y(n4714) );
  XOR2XL U21095 ( .A(n7528), .B(n20220), .Y(n19834) );
  INVXL U21096 ( .A(n20217), .Y(n19830) );
  XOR2X1 U21097 ( .A(n19820), .B(n19819), .Y(n19821) );
  INVXL U21098 ( .A(n20205), .Y(n19819) );
  INVXL U21099 ( .A(n20202), .Y(n19815) );
  INVXL U21100 ( .A(n20197), .Y(n19808) );
  XNOR2XL U21101 ( .A(n19790), .B(U1_A_r_d0[25]), .Y(n7527) );
  MXI2XL U21102 ( .A(U1_pipe13[0]), .B(n20458), .S0(n20240), .Y(n4723) );
  MXI2XL U21103 ( .A(U1_pipe13[1]), .B(n20178), .S0(n20240), .Y(n4724) );
  INVXL U21104 ( .A(n20456), .Y(n20177) );
  MXI2XL U21105 ( .A(U1_pipe13[2]), .B(n20174), .S0(n20025), .Y(n4725) );
  INVXL U21106 ( .A(n20453), .Y(n20173) );
  MXI2XL U21107 ( .A(U1_pipe13[3]), .B(n20168), .S0(n20025), .Y(n4726) );
  INVXL U21108 ( .A(n20449), .Y(n20166) );
  MXI2XL U21109 ( .A(U1_pipe13[4]), .B(n20164), .S0(n20025), .Y(n4727) );
  NAND2XL U21110 ( .A(n20161), .B(n20160), .Y(n20162) );
  MXI2XL U21111 ( .A(U1_pipe13[5]), .B(n20155), .S0(n20025), .Y(n4728) );
  XNOR2XL U21112 ( .A(n20154), .B(n20153), .Y(n20155) );
  NAND2XL U21113 ( .A(n20152), .B(n20151), .Y(n20153) );
  XOR2XL U21114 ( .A(n20149), .B(n20148), .Y(n20150) );
  NAND2XL U21115 ( .A(n20147), .B(n20146), .Y(n20148) );
  AOI21XL U21116 ( .A0(n20154), .A1(n20152), .B0(n20144), .Y(n20149) );
  XOR2XL U21117 ( .A(n20141), .B(n20140), .Y(n20142) );
  NAND2XL U21118 ( .A(n19950), .B(n20139), .Y(n20140) );
  XOR2XL U21119 ( .A(n20134), .B(n20133), .Y(n20135) );
  INVXL U21120 ( .A(n20416), .Y(n20133) );
  NAND2XL U21121 ( .A(n20123), .B(n20122), .Y(n20124) );
  AOI21XL U21122 ( .A0(n20130), .A1(n20128), .B0(n20120), .Y(n20125) );
  NAND2XL U21123 ( .A(n20108), .B(n20107), .Y(n20109) );
  NAND2XL U21124 ( .A(n20090), .B(n20089), .Y(n20091) );
  NAND2XL U21125 ( .A(n20085), .B(n20084), .Y(n20086) );
  INVXL U21126 ( .A(n20360), .Y(n20076) );
  INVXL U21127 ( .A(n20357), .Y(n20073) );
  INVXL U21128 ( .A(n20352), .Y(n20066) );
  NAND2XL U21129 ( .A(n20061), .B(n20060), .Y(n20062) );
  INVXL U21130 ( .A(n20349), .Y(n20052) );
  MXI2XL U21131 ( .A(U1_pipe14[0]), .B(n17595), .S0(n5809), .Y(n4751) );
  MXI2XL U21132 ( .A(U1_pipe14[1]), .B(n17295), .S0(n22853), .Y(n4752) );
  MXI2XL U21133 ( .A(U1_pipe14[2]), .B(n17292), .S0(n22853), .Y(n4753) );
  MXI2XL U21134 ( .A(U1_pipe14[3]), .B(n17287), .S0(n22853), .Y(n4754) );
  XOR2XL U21135 ( .A(n17286), .B(n17583), .Y(n17287) );
  MXI2XL U21136 ( .A(U1_pipe14[4]), .B(n17282), .S0(n22853), .Y(n4755) );
  XNOR2XL U21137 ( .A(n17281), .B(n17579), .Y(n17282) );
  MXI2XL U21138 ( .A(U1_pipe14[5]), .B(n17276), .S0(n22853), .Y(n4756) );
  XNOR2XL U21139 ( .A(n17275), .B(n17572), .Y(n17276) );
  XOR2XL U21140 ( .A(n17271), .B(n17568), .Y(n17272) );
  AOI21XL U21141 ( .A0(n17275), .A1(n17274), .B0(n17267), .Y(n17271) );
  INVXL U21142 ( .A(n17273), .Y(n17267) );
  XOR2XL U21143 ( .A(n17264), .B(n17560), .Y(n17265) );
  XOR2XL U21144 ( .A(n17257), .B(n17553), .Y(n17258) );
  XNOR2XL U21145 ( .A(n17253), .B(n17549), .Y(n17254) );
  AOI21XL U21146 ( .A0(n17253), .A1(n17252), .B0(n17244), .Y(n17248) );
  XNOR2XL U21147 ( .A(n17240), .B(n17535), .Y(n17241) );
  XOR2XL U21148 ( .A(n17237), .B(n17531), .Y(n17238) );
  MXI2XL U21149 ( .A(U1_pipe14[13]), .B(n17231), .S0(n5809), .Y(n4764) );
  XNOR2XL U21150 ( .A(n17230), .B(n17522), .Y(n17231) );
  XOR2XL U21151 ( .A(n17226), .B(n17518), .Y(n17227) );
  AOI21XL U21152 ( .A0(n17230), .A1(n17229), .B0(n17224), .Y(n17226) );
  XOR2XL U21153 ( .A(n17222), .B(n17512), .Y(n17223) );
  OAI21XL U21154 ( .A0(n17222), .A1(n17215), .B0(n17220), .Y(n17218) );
  XNOR2XL U21155 ( .A(n17209), .B(n17498), .Y(n17210) );
  INVX1 U21156 ( .A(n17209), .Y(n17203) );
  XOR2XL U21157 ( .A(n17200), .B(n17487), .Y(n17201) );
  XNOR2X1 U21158 ( .A(n13729), .B(n17483), .Y(n13730) );
  XOR2X1 U21159 ( .A(n17196), .B(n17475), .Y(n17197) );
  XOR2XL U21160 ( .A(n7320), .B(n17458), .Y(n17179) );
  AOI21XL U21161 ( .A0(n17180), .A1(n9604), .B0(n9603), .Y(n7320) );
  MXI2XL U21162 ( .A(U1_pipe15[0]), .B(n17742), .S0(n5805), .Y(n4779) );
  MXI2XL U21163 ( .A(U1_pipe15[1]), .B(n17445), .S0(n6887), .Y(n4780) );
  NAND2XL U21164 ( .A(n17442), .B(n17441), .Y(n17444) );
  MXI2XL U21165 ( .A(U1_pipe15[2]), .B(n17440), .S0(n6887), .Y(n4781) );
  NAND2XL U21166 ( .A(n13535), .B(n17437), .Y(n17438) );
  MXI2XL U21167 ( .A(U1_pipe15[3]), .B(n17435), .S0(n22853), .Y(n4782) );
  XOR2XL U21168 ( .A(n17434), .B(n17433), .Y(n17435) );
  NAND2XL U21169 ( .A(n17432), .B(n17431), .Y(n17433) );
  INVXL U21170 ( .A(n17430), .Y(n17432) );
  XNOR2XL U21171 ( .A(n17428), .B(n17427), .Y(n17429) );
  NAND2XL U21172 ( .A(n17426), .B(n17425), .Y(n17427) );
  XNOR2XL U21173 ( .A(n17421), .B(n17420), .Y(n17422) );
  NAND2XL U21174 ( .A(n17419), .B(n17418), .Y(n17420) );
  XOR2XL U21175 ( .A(n17416), .B(n17415), .Y(n17417) );
  NAND2XL U21176 ( .A(n17414), .B(n17413), .Y(n17415) );
  AOI21XL U21177 ( .A0(n17421), .A1(n17419), .B0(n17411), .Y(n17416) );
  XOR2XL U21178 ( .A(n17408), .B(n17407), .Y(n17409) );
  NAND2XL U21179 ( .A(n13534), .B(n17406), .Y(n17407) );
  MXI2XL U21180 ( .A(U1_pipe15[8]), .B(n17402), .S0(n25330), .Y(n4787) );
  XOR2XL U21181 ( .A(n17401), .B(n17695), .Y(n17402) );
  NAND2XL U21182 ( .A(n17390), .B(n17389), .Y(n17391) );
  AOI21XL U21183 ( .A0(n17397), .A1(n17395), .B0(n17387), .Y(n17392) );
  NAND2XL U21184 ( .A(n17377), .B(n17376), .Y(n17378) );
  NAND2XL U21185 ( .A(n17364), .B(n17363), .Y(n17365) );
  XOR2X1 U21186 ( .A(n17360), .B(n17653), .Y(n17361) );
  INVXL U21187 ( .A(n17359), .Y(n17353) );
  NAND2X1 U21188 ( .A(n17304), .B(n7552), .Y(n7551) );
  MXI2XL U21189 ( .A(n7505), .B(U1_pipe15[27]), .S0(n17032), .Y(n4806) );
  MXI2XL U21190 ( .A(U1_pipe0[0]), .B(n19504), .S0(n19405), .Y(n4807) );
  MXI2XL U21191 ( .A(U1_pipe9[0]), .B(n20458), .S0(n20438), .Y(n4810) );
  MXI2XL U21192 ( .A(U1_pipe9[1]), .B(n20457), .S0(n20438), .Y(n4811) );
  MXI2XL U21193 ( .A(U1_pipe9[2]), .B(n20454), .S0(n20438), .Y(n4812) );
  MXI2XL U21194 ( .A(U1_pipe9[3]), .B(n20451), .S0(n20438), .Y(n4813) );
  XOR2XL U21195 ( .A(n20450), .B(n20449), .Y(n20451) );
  MXI2XL U21196 ( .A(U1_pipe9[4]), .B(n20448), .S0(n20438), .Y(n4814) );
  NAND2XL U21197 ( .A(n20445), .B(n20444), .Y(n20446) );
  MXI2XL U21198 ( .A(U1_pipe9[5]), .B(n20439), .S0(n20438), .Y(n4815) );
  XNOR2XL U21199 ( .A(n20437), .B(n20436), .Y(n20439) );
  NAND2XL U21200 ( .A(n20435), .B(n20434), .Y(n20436) );
  XOR2XL U21201 ( .A(n20432), .B(n20431), .Y(n20433) );
  NAND2XL U21202 ( .A(n20430), .B(n20429), .Y(n20431) );
  AOI21XL U21203 ( .A0(n20437), .A1(n20435), .B0(n20427), .Y(n20432) );
  XOR2XL U21204 ( .A(n20424), .B(n20423), .Y(n20425) );
  NAND2XL U21205 ( .A(n14865), .B(n20422), .Y(n20423) );
  XOR2XL U21206 ( .A(n20417), .B(n20416), .Y(n20418) );
  NAND2XL U21207 ( .A(n20407), .B(n20406), .Y(n20408) );
  AOI21XL U21208 ( .A0(n20414), .A1(n20412), .B0(n20404), .Y(n20409) );
  NAND2XL U21209 ( .A(n20393), .B(n20392), .Y(n20394) );
  XNOR2XL U21210 ( .A(n20386), .B(n20385), .Y(n20387) );
  NAND2XL U21211 ( .A(n20384), .B(n20383), .Y(n20385) );
  XOR2XL U21212 ( .A(n20381), .B(n20380), .Y(n20382) );
  NAND2XL U21213 ( .A(n20379), .B(n20378), .Y(n20380) );
  AOI21XL U21214 ( .A0(n20386), .A1(n20384), .B0(n20377), .Y(n20381) );
  XOR2XL U21215 ( .A(n20375), .B(n20374), .Y(n20376) );
  XNOR2XL U21216 ( .A(n20361), .B(n20360), .Y(n20362) );
  NAND2XL U21217 ( .A(n20361), .B(n20356), .Y(n7444) );
  XOR2X1 U21218 ( .A(n20353), .B(n20352), .Y(n20354) );
  INVXL U21219 ( .A(n7478), .Y(n7436) );
  MXI2XL U21220 ( .A(U1_pipe10[0]), .B(n17595), .S0(n5812), .Y(n4838) );
  MXI2XL U21221 ( .A(U1_pipe10[1]), .B(n17594), .S0(n17641), .Y(n4839) );
  INVXL U21222 ( .A(n17591), .Y(n17593) );
  MXI2XL U21223 ( .A(U1_pipe10[2]), .B(n17590), .S0(n5809), .Y(n4840) );
  INVXL U21224 ( .A(n17587), .Y(n17589) );
  MXI2XL U21225 ( .A(U1_pipe10[3]), .B(n17586), .S0(n5809), .Y(n4841) );
  XOR2XL U21226 ( .A(n17585), .B(n17584), .Y(n17586) );
  INVXL U21227 ( .A(n17583), .Y(n17584) );
  MXI2XL U21228 ( .A(U1_pipe10[4]), .B(n17582), .S0(n5809), .Y(n4842) );
  XNOR2XL U21229 ( .A(n17581), .B(n17580), .Y(n17582) );
  INVXL U21230 ( .A(n17579), .Y(n17580) );
  MXI2XL U21231 ( .A(U1_pipe10[5]), .B(n17575), .S0(n5809), .Y(n4843) );
  XNOR2XL U21232 ( .A(n17574), .B(n17573), .Y(n17575) );
  INVXL U21233 ( .A(n17572), .Y(n17573) );
  MXI2XL U21234 ( .A(U1_pipe10[6]), .B(n17571), .S0(n5809), .Y(n4844) );
  INVXL U21235 ( .A(n17568), .Y(n17569) );
  AOI21XL U21236 ( .A0(n17574), .A1(n17567), .B0(n17566), .Y(n17570) );
  MXI2XL U21237 ( .A(U1_pipe10[7]), .B(n17563), .S0(n5809), .Y(n4845) );
  XOR2XL U21238 ( .A(n17562), .B(n17561), .Y(n17563) );
  INVXL U21239 ( .A(n17560), .Y(n17561) );
  MXI2XL U21240 ( .A(U1_pipe10[8]), .B(n17556), .S0(n5809), .Y(n4846) );
  XOR2XL U21241 ( .A(n17555), .B(n17554), .Y(n17556) );
  INVXL U21242 ( .A(n17553), .Y(n17554) );
  INVXL U21243 ( .A(n17549), .Y(n17550) );
  INVXL U21244 ( .A(n17545), .Y(n17546) );
  AOI21XL U21245 ( .A0(n17551), .A1(n17544), .B0(n17543), .Y(n17547) );
  INVXL U21246 ( .A(n17535), .Y(n17536) );
  INVXL U21247 ( .A(n17531), .Y(n17532) );
  AOI21XL U21248 ( .A0(n17537), .A1(n17530), .B0(n17529), .Y(n17533) );
  MXI2XL U21249 ( .A(U1_pipe10[13]), .B(n17525), .S0(n5809), .Y(n4851) );
  XNOR2XL U21250 ( .A(n17524), .B(n17523), .Y(n17525) );
  INVXL U21251 ( .A(n17522), .Y(n17523) );
  XOR2XL U21252 ( .A(n17520), .B(n17519), .Y(n17521) );
  INVXL U21253 ( .A(n17518), .Y(n17519) );
  XOR2XL U21254 ( .A(n17514), .B(n17513), .Y(n17515) );
  INVXL U21255 ( .A(n17512), .Y(n17513) );
  INVXL U21256 ( .A(n17508), .Y(n17509) );
  OAI21XL U21257 ( .A0(n17514), .A1(n17507), .B0(n17506), .Y(n17510) );
  INVXL U21258 ( .A(n17498), .Y(n17499) );
  INVXL U21259 ( .A(n17494), .Y(n17495) );
  INVXL U21260 ( .A(n17483), .Y(n17484) );
  MXI2XL U21261 ( .A(U1_pipe11[0]), .B(n17742), .S0(n24784), .Y(n4866) );
  MXI2XL U21262 ( .A(U1_pipe11[1]), .B(n17741), .S0(n5812), .Y(n4867) );
  NAND2XL U21263 ( .A(n12860), .B(n17738), .Y(n17740) );
  MXI2XL U21264 ( .A(U1_pipe11[2]), .B(n17737), .S0(n24784), .Y(n4868) );
  NAND2XL U21265 ( .A(n17734), .B(n17733), .Y(n17736) );
  INVXL U21266 ( .A(n17732), .Y(n17734) );
  MXI2XL U21267 ( .A(U1_pipe11[3]), .B(n17731), .S0(n25330), .Y(n4869) );
  XOR2XL U21268 ( .A(n17730), .B(n17729), .Y(n17731) );
  NAND2XL U21269 ( .A(n17728), .B(n17727), .Y(n17729) );
  INVXL U21270 ( .A(n17726), .Y(n17728) );
  MXI2XL U21271 ( .A(U1_pipe11[4]), .B(n17725), .S0(n5812), .Y(n4870) );
  XNOR2XL U21272 ( .A(n17724), .B(n17723), .Y(n17725) );
  NAND2XL U21273 ( .A(n17722), .B(n17721), .Y(n17723) );
  MXI2XL U21274 ( .A(U1_pipe11[5]), .B(n17718), .S0(n5812), .Y(n4871) );
  XNOR2XL U21275 ( .A(n17717), .B(n17716), .Y(n17718) );
  NAND2XL U21276 ( .A(n17715), .B(n17714), .Y(n17716) );
  XOR2XL U21277 ( .A(n17712), .B(n17711), .Y(n17713) );
  NAND2XL U21278 ( .A(n17710), .B(n17709), .Y(n17711) );
  AOI21XL U21279 ( .A0(n17717), .A1(n17715), .B0(n17707), .Y(n17712) );
  MXI2XL U21280 ( .A(U1_pipe11[7]), .B(n17705), .S0(n25330), .Y(n4873) );
  XOR2XL U21281 ( .A(n17704), .B(n17703), .Y(n17705) );
  NAND2XL U21282 ( .A(n12795), .B(n17702), .Y(n17703) );
  AOI21XL U21283 ( .A0(n17717), .A1(n17701), .B0(n17700), .Y(n17704) );
  MXI2XL U21284 ( .A(U1_pipe11[8]), .B(n17698), .S0(n5812), .Y(n4874) );
  XOR2XL U21285 ( .A(n17697), .B(n17696), .Y(n17698) );
  INVXL U21286 ( .A(n17695), .Y(n17696) );
  NAND2XL U21287 ( .A(n17691), .B(n17690), .Y(n17692) );
  NAND2XL U21288 ( .A(n17686), .B(n17685), .Y(n17687) );
  AOI21XL U21289 ( .A0(n17693), .A1(n17691), .B0(n17683), .Y(n17688) );
  NAND2XL U21290 ( .A(n17676), .B(n17675), .Y(n17677) );
  NAND2XL U21291 ( .A(n17671), .B(n17670), .Y(n17672) );
  NAND2XL U21292 ( .A(n13034), .B(n17662), .Y(n17663) );
  INVXL U21293 ( .A(n17653), .Y(n17654) );
  INVXL U21294 ( .A(n17649), .Y(n17650) );
  NAND2XL U21295 ( .A(n17639), .B(n17638), .Y(n17640) );
  INVXL U21296 ( .A(n17634), .Y(n17635) );
  NAND2XL U21297 ( .A(n17623), .B(n17622), .Y(n17624) );
  INVXL U21298 ( .A(n17617), .Y(n17618) );
  INVXL U21299 ( .A(n17613), .Y(n17614) );
  MXI2XL U21300 ( .A(U1_pipe12[0]), .B(n20307), .S0(n20240), .Y(n4894) );
  MXI2XL U21301 ( .A(U1_pipe12[1]), .B(n19949), .S0(n20240), .Y(n4895) );
  INVXL U21302 ( .A(n20305), .Y(n19948) );
  MXI2XL U21303 ( .A(U1_pipe12[2]), .B(n19945), .S0(n20240), .Y(n4896) );
  INVXL U21304 ( .A(n20302), .Y(n19944) );
  MXI2XL U21305 ( .A(U1_pipe12[3]), .B(n19939), .S0(n20240), .Y(n4897) );
  XOR2XL U21306 ( .A(n19938), .B(n19937), .Y(n19939) );
  INVXL U21307 ( .A(n20298), .Y(n19937) );
  MXI2XL U21308 ( .A(U1_pipe12[4]), .B(n19935), .S0(n20240), .Y(n4898) );
  XNOR2XL U21309 ( .A(n19934), .B(n19933), .Y(n19935) );
  INVXL U21310 ( .A(n20295), .Y(n19933) );
  MXI2XL U21311 ( .A(U1_pipe12[5]), .B(n19926), .S0(n20240), .Y(n4899) );
  XNOR2XL U21312 ( .A(n19925), .B(n19924), .Y(n19926) );
  INVXL U21313 ( .A(n20289), .Y(n19924) );
  MXI2XL U21314 ( .A(U1_pipe12[6]), .B(n19922), .S0(n20240), .Y(n4900) );
  XOR2XL U21315 ( .A(n19921), .B(n19920), .Y(n19922) );
  INVXL U21316 ( .A(n20286), .Y(n19920) );
  AOI21XL U21317 ( .A0(n19925), .A1(n19916), .B0(n19915), .Y(n19921) );
  MXI2XL U21318 ( .A(U1_pipe12[7]), .B(n19912), .S0(n20240), .Y(n4901) );
  XOR2XL U21319 ( .A(n19911), .B(n19910), .Y(n19912) );
  INVXL U21320 ( .A(n20280), .Y(n19910) );
  MXI2XL U21321 ( .A(U1_pipe12[8]), .B(n19905), .S0(n20240), .Y(n4902) );
  XOR2XL U21322 ( .A(n19904), .B(n19903), .Y(n19905) );
  INVXL U21323 ( .A(n20274), .Y(n19903) );
  INVXL U21324 ( .A(n20271), .Y(n19899) );
  INVXL U21325 ( .A(n20268), .Y(n19895) );
  AOI21XL U21326 ( .A0(n19900), .A1(n19891), .B0(n19890), .Y(n19896) );
  INVXL U21327 ( .A(n20260), .Y(n19883) );
  INVXL U21328 ( .A(n20257), .Y(n19879) );
  MXI2XL U21329 ( .A(U1_pipe0[1]), .B(n19503), .S0(n19405), .Y(n4907) );
  XOR2XL U21330 ( .A(n17112), .B(n17111), .Y(n17113) );
  AOI21XL U21331 ( .A0(n17115), .A1(n13881), .B0(n17110), .Y(n17112) );
  XNOR2X1 U21332 ( .A(n5966), .B(n17105), .Y(n17106) );
  NAND2XL U21333 ( .A(n17099), .B(n17098), .Y(n17100) );
  XNOR2XL U21334 ( .A(n17081), .B(n17080), .Y(n17082) );
  XOR2XL U21335 ( .A(n17072), .B(n17071), .Y(n17073) );
  MXI2XL U21336 ( .A(U1_pipe6[0]), .B(n17049), .S0(n25330), .Y(n4925) );
  MXI2XL U21337 ( .A(U1_pipe6[1]), .B(n16779), .S0(n25267), .Y(n4926) );
  INVXL U21338 ( .A(n17047), .Y(n16778) );
  MXI2XL U21339 ( .A(U1_pipe6[2]), .B(n16775), .S0(n25330), .Y(n4927) );
  INVXL U21340 ( .A(n17044), .Y(n16774) );
  MXI2XL U21341 ( .A(U1_pipe6[3]), .B(n16769), .S0(n5812), .Y(n4928) );
  XOR2XL U21342 ( .A(n16768), .B(n16767), .Y(n16769) );
  INVXL U21343 ( .A(n17040), .Y(n16767) );
  MXI2XL U21344 ( .A(U1_pipe6[4]), .B(n16765), .S0(n25330), .Y(n4929) );
  XNOR2XL U21345 ( .A(n16764), .B(n16763), .Y(n16765) );
  INVXL U21346 ( .A(n17037), .Y(n16763) );
  MXI2XL U21347 ( .A(U1_pipe6[5]), .B(n16756), .S0(n5812), .Y(n4930) );
  XNOR2XL U21348 ( .A(n16755), .B(n16754), .Y(n16756) );
  INVXL U21349 ( .A(n17030), .Y(n16754) );
  MXI2XL U21350 ( .A(U1_pipe6[6]), .B(n16752), .S0(n25330), .Y(n4931) );
  XOR2XL U21351 ( .A(n16751), .B(n16750), .Y(n16752) );
  INVXL U21352 ( .A(n17027), .Y(n16750) );
  AOI21XL U21353 ( .A0(n16755), .A1(n16747), .B0(n16746), .Y(n16751) );
  MXI2XL U21354 ( .A(U1_pipe6[7]), .B(n16743), .S0(n25330), .Y(n4932) );
  XOR2XL U21355 ( .A(n16742), .B(n16741), .Y(n16743) );
  INVXL U21356 ( .A(n17021), .Y(n16741) );
  AOI21XL U21357 ( .A0(n16755), .A1(n16738), .B0(n16737), .Y(n16742) );
  MXI2XL U21358 ( .A(U1_pipe6[8]), .B(n16735), .S0(n5812), .Y(n4933) );
  XOR2XL U21359 ( .A(n16734), .B(n16733), .Y(n16735) );
  INVXL U21360 ( .A(n17015), .Y(n16733) );
  MXI2XL U21361 ( .A(U1_pipe6[9]), .B(n16731), .S0(n25330), .Y(n4934) );
  INVXL U21362 ( .A(n17012), .Y(n16729) );
  INVXL U21363 ( .A(n17009), .Y(n16725) );
  AOI21XL U21364 ( .A0(n16730), .A1(n16721), .B0(n16720), .Y(n16726) );
  MXI2XL U21365 ( .A(U1_pipe6[11]), .B(n16715), .S0(n25330), .Y(n4936) );
  INVXL U21366 ( .A(n17001), .Y(n16713) );
  INVXL U21367 ( .A(n16998), .Y(n16709) );
  AOI21XL U21368 ( .A0(n16714), .A1(n16706), .B0(n16705), .Y(n16710) );
  MXI2XL U21369 ( .A(U1_pipe6[13]), .B(n16701), .S0(n25330), .Y(n4938) );
  XNOR2XL U21370 ( .A(n16700), .B(n16699), .Y(n16701) );
  INVXL U21371 ( .A(n16992), .Y(n16699) );
  XOR2XL U21372 ( .A(n16696), .B(n16695), .Y(n16697) );
  INVXL U21373 ( .A(n16989), .Y(n16695) );
  XOR2XL U21374 ( .A(n16690), .B(n16689), .Y(n16691) );
  INVXL U21375 ( .A(n16984), .Y(n16689) );
  INVXL U21376 ( .A(n16981), .Y(n16685) );
  INVXL U21377 ( .A(n16973), .Y(n16675) );
  INVXL U21378 ( .A(n16970), .Y(n16671) );
  MXI2XL U21379 ( .A(U1_pipe6[20]), .B(n16664), .S0(n25330), .Y(n4945) );
  INVXL U21380 ( .A(n16962), .Y(n16662) );
  MXI2XL U21381 ( .A(U1_pipe6[21]), .B(n16653), .S0(n25330), .Y(n4946) );
  INVXL U21382 ( .A(n16955), .Y(n16651) );
  MXI2XL U21383 ( .A(U1_pipe6[24]), .B(n16639), .S0(n25330), .Y(n4949) );
  NAND2XL U21384 ( .A(n7167), .B(n7401), .Y(n16638) );
  MXI2XL U21385 ( .A(U1_pipe6[25]), .B(n16632), .S0(n25330), .Y(n4950) );
  MXI2XL U21386 ( .A(U1_pipe7[0]), .B(n17166), .S0(n5812), .Y(n4953) );
  MXI2XL U21387 ( .A(U1_pipe7[1]), .B(n16931), .S0(n17641), .Y(n4954) );
  INVXL U21388 ( .A(n17164), .Y(n16930) );
  MXI2XL U21389 ( .A(U1_pipe7[2]), .B(n16927), .S0(n5812), .Y(n4955) );
  INVXL U21390 ( .A(n17161), .Y(n16926) );
  MXI2XL U21391 ( .A(U1_pipe7[3]), .B(n16921), .S0(n24784), .Y(n4956) );
  XOR2XL U21392 ( .A(n16920), .B(n16919), .Y(n16921) );
  INVXL U21393 ( .A(n17157), .Y(n16919) );
  MXI2XL U21394 ( .A(U1_pipe7[4]), .B(n16917), .S0(n5804), .Y(n4957) );
  XNOR2XL U21395 ( .A(n16916), .B(n16915), .Y(n16917) );
  INVXL U21396 ( .A(n17154), .Y(n16915) );
  MXI2XL U21397 ( .A(U1_pipe7[5]), .B(n16908), .S0(n5804), .Y(n4958) );
  XNOR2XL U21398 ( .A(n16907), .B(n16906), .Y(n16908) );
  NAND2XL U21399 ( .A(n16905), .B(n16904), .Y(n16906) );
  MXI2XL U21400 ( .A(U1_pipe7[6]), .B(n16903), .S0(n5804), .Y(n4959) );
  XOR2XL U21401 ( .A(n16902), .B(n16901), .Y(n16903) );
  NAND2XL U21402 ( .A(n16900), .B(n16899), .Y(n16901) );
  AOI21XL U21403 ( .A0(n16907), .A1(n16905), .B0(n16897), .Y(n16902) );
  MXI2XL U21404 ( .A(U1_pipe7[7]), .B(n16895), .S0(n5804), .Y(n4960) );
  XOR2XL U21405 ( .A(n16894), .B(n16893), .Y(n16895) );
  NAND2XL U21406 ( .A(n14903), .B(n16892), .Y(n16893) );
  MXI2XL U21407 ( .A(U1_pipe7[8]), .B(n16888), .S0(n5804), .Y(n4961) );
  XOR2XL U21408 ( .A(n16887), .B(n16886), .Y(n16888) );
  INVXL U21409 ( .A(n17128), .Y(n16886) );
  INVXL U21410 ( .A(n17125), .Y(n16882) );
  INVXL U21411 ( .A(n17122), .Y(n16878) );
  AOI21XL U21412 ( .A0(n16883), .A1(n16874), .B0(n16873), .Y(n16879) );
  INVXL U21413 ( .A(n17114), .Y(n16866) );
  INVXL U21414 ( .A(n17111), .Y(n16862) );
  NAND2XL U21415 ( .A(n16849), .B(n16848), .Y(n16850) );
  NAND2XL U21416 ( .A(n16843), .B(n16842), .Y(n16844) );
  NAND2XL U21417 ( .A(n16838), .B(n16837), .Y(n16839) );
  MXI2XL U21418 ( .A(U1_pipe7[17]), .B(n16833), .S0(n25330), .Y(n4970) );
  INVXL U21419 ( .A(n17080), .Y(n16831) );
  MXI2XL U21420 ( .A(U1_pipe7[18]), .B(n16829), .S0(n25330), .Y(n4971) );
  INVXL U21421 ( .A(n17077), .Y(n16827) );
  MXI2XL U21422 ( .A(U1_pipe7[19]), .B(n16822), .S0(n25330), .Y(n4972) );
  INVXL U21423 ( .A(n17071), .Y(n16820) );
  INVXL U21424 ( .A(n16814), .Y(n16815) );
  INVXL U21425 ( .A(n17068), .Y(n16805) );
  MXI2XL U21426 ( .A(U1_pipe8[0]), .B(n20307), .S0(n20240), .Y(n4981) );
  MXI2XL U21427 ( .A(U1_pipe8[1]), .B(n20306), .S0(n20240), .Y(n4982) );
  MXI2XL U21428 ( .A(U1_pipe8[2]), .B(n20303), .S0(n20240), .Y(n4983) );
  MXI2XL U21429 ( .A(U1_pipe8[3]), .B(n20300), .S0(n20240), .Y(n4984) );
  XOR2XL U21430 ( .A(n20299), .B(n20298), .Y(n20300) );
  MXI2XL U21431 ( .A(U1_pipe8[4]), .B(n20297), .S0(n20240), .Y(n4985) );
  XNOR2XL U21432 ( .A(n20296), .B(n20295), .Y(n20297) );
  MXI2XL U21433 ( .A(U1_pipe8[5]), .B(n20291), .S0(n20240), .Y(n4986) );
  XNOR2XL U21434 ( .A(n20290), .B(n20289), .Y(n20291) );
  MXI2XL U21435 ( .A(U1_pipe8[6]), .B(n20288), .S0(n20240), .Y(n4987) );
  XOR2XL U21436 ( .A(n20287), .B(n20286), .Y(n20288) );
  AOI21XL U21437 ( .A0(n20290), .A1(n20285), .B0(n20284), .Y(n20287) );
  INVXL U21438 ( .A(n20283), .Y(n20284) );
  MXI2XL U21439 ( .A(U1_pipe8[7]), .B(n20282), .S0(n20240), .Y(n4988) );
  XOR2XL U21440 ( .A(n20281), .B(n20280), .Y(n20282) );
  AOI21XL U21441 ( .A0(n20290), .A1(n20279), .B0(n20278), .Y(n20281) );
  MXI2XL U21442 ( .A(U1_pipe8[8]), .B(n20276), .S0(n20240), .Y(n4989) );
  XOR2XL U21443 ( .A(n20275), .B(n20274), .Y(n20276) );
  XNOR2XL U21444 ( .A(n20272), .B(n20271), .Y(n20273) );
  XOR2XL U21445 ( .A(n20269), .B(n20268), .Y(n20270) );
  AOI21XL U21446 ( .A0(n20272), .A1(n20267), .B0(n20266), .Y(n20269) );
  INVXL U21447 ( .A(n20265), .Y(n20266) );
  XNOR2XL U21448 ( .A(n20261), .B(n20260), .Y(n20262) );
  XOR2XL U21449 ( .A(n20258), .B(n20257), .Y(n20259) );
  XNOR2XL U21450 ( .A(n20251), .B(n20250), .Y(n20252) );
  XOR2XL U21451 ( .A(n20248), .B(n20247), .Y(n20249) );
  AOI21XL U21452 ( .A0(n20251), .A1(n20246), .B0(n20245), .Y(n20248) );
  XOR2XL U21453 ( .A(n20243), .B(n20242), .Y(n20244) );
  XNOR2XL U21454 ( .A(n20230), .B(n20229), .Y(n20231) );
  XOR2XL U21455 ( .A(n20221), .B(n20220), .Y(n20222) );
  XOR2XL U21456 ( .A(n20206), .B(n20205), .Y(n20207) );
  XOR2XL U21457 ( .A(n7304), .B(n20192), .Y(n20193) );
  MXI2XL U21458 ( .A(U1_pipe0[2]), .B(n19500), .S0(n19405), .Y(n5007) );
  MXI2XL U21459 ( .A(U1_pipe2[0]), .B(n19504), .S0(n19215), .Y(n5012) );
  MXI2XL U21460 ( .A(U1_pipe2[1]), .B(n19230), .S0(n19215), .Y(n5013) );
  INVXL U21461 ( .A(n19502), .Y(n19229) );
  MXI2XL U21462 ( .A(U1_pipe2[2]), .B(n19226), .S0(n19215), .Y(n5014) );
  INVXL U21463 ( .A(n19499), .Y(n19225) );
  MXI2XL U21464 ( .A(U1_pipe2[3]), .B(n19220), .S0(n19215), .Y(n5015) );
  XOR2XL U21465 ( .A(n19219), .B(n19218), .Y(n19220) );
  INVXL U21466 ( .A(n19495), .Y(n19218) );
  MXI2XL U21467 ( .A(U1_pipe2[4]), .B(n19216), .S0(n19215), .Y(n5016) );
  XNOR2XL U21468 ( .A(n19214), .B(n19213), .Y(n19216) );
  INVXL U21469 ( .A(n19492), .Y(n19213) );
  XNOR2XL U21470 ( .A(n19205), .B(n19204), .Y(n19206) );
  INVXL U21471 ( .A(n19486), .Y(n19204) );
  XOR2XL U21472 ( .A(n19201), .B(n19200), .Y(n19202) );
  INVXL U21473 ( .A(n19483), .Y(n19200) );
  AOI21XL U21474 ( .A0(n19205), .A1(n19196), .B0(n19195), .Y(n19201) );
  XOR2XL U21475 ( .A(n19191), .B(n19190), .Y(n19192) );
  INVXL U21476 ( .A(n19477), .Y(n19190) );
  XOR2XL U21477 ( .A(n19184), .B(n19183), .Y(n19185) );
  INVXL U21478 ( .A(n19471), .Y(n19183) );
  INVXL U21479 ( .A(n19468), .Y(n19179) );
  INVXL U21480 ( .A(n19465), .Y(n19175) );
  AOI21XL U21481 ( .A0(n19180), .A1(n19171), .B0(n19170), .Y(n19176) );
  INVXL U21482 ( .A(n19457), .Y(n19163) );
  INVXL U21483 ( .A(n19454), .Y(n19159) );
  AOI21XL U21484 ( .A0(n19164), .A1(n19156), .B0(n19155), .Y(n19160) );
  INVXL U21485 ( .A(n19448), .Y(n19149) );
  XOR2XL U21486 ( .A(n19146), .B(n19145), .Y(n19147) );
  INVXL U21487 ( .A(n19445), .Y(n19145) );
  XOR2XL U21488 ( .A(n19140), .B(n19139), .Y(n19141) );
  INVXL U21489 ( .A(n19440), .Y(n19139) );
  INVXL U21490 ( .A(n19437), .Y(n19135) );
  INVXL U21491 ( .A(n19428), .Y(n19124) );
  INVXL U21492 ( .A(n19425), .Y(n19120) );
  INVXL U21493 ( .A(n19416), .Y(n19109) );
  XOR2X1 U21494 ( .A(n19100), .B(n19099), .Y(n19101) );
  MXI2XL U21495 ( .A(U1_pipe3[0]), .B(n19701), .S0(n19405), .Y(n5040) );
  MXI2XL U21496 ( .A(U1_pipe3[1]), .B(n19376), .S0(n19405), .Y(n5041) );
  INVXL U21497 ( .A(n19699), .Y(n19375) );
  MXI2XL U21498 ( .A(U1_pipe3[2]), .B(n19372), .S0(n19405), .Y(n5042) );
  INVXL U21499 ( .A(n19695), .Y(n19371) );
  MXI2XL U21500 ( .A(U1_pipe3[3]), .B(n19367), .S0(n19405), .Y(n5043) );
  XOR2XL U21501 ( .A(n19366), .B(n19365), .Y(n19367) );
  INVXL U21502 ( .A(n19690), .Y(n19365) );
  INVXL U21503 ( .A(n19687), .Y(n19360) );
  XNOR2XL U21504 ( .A(n19353), .B(n19352), .Y(n19354) );
  NAND2XL U21505 ( .A(n19351), .B(n19350), .Y(n19352) );
  XOR2XL U21506 ( .A(n19348), .B(n19347), .Y(n19349) );
  NAND2XL U21507 ( .A(n19346), .B(n19345), .Y(n19347) );
  AOI21XL U21508 ( .A0(n19353), .A1(n19351), .B0(n19343), .Y(n19348) );
  XOR2XL U21509 ( .A(n19340), .B(n19339), .Y(n19341) );
  NAND2XL U21510 ( .A(n19338), .B(n19337), .Y(n19339) );
  XOR2XL U21511 ( .A(n19332), .B(n19331), .Y(n19333) );
  INVXL U21512 ( .A(n19661), .Y(n19331) );
  INVXL U21513 ( .A(n19658), .Y(n19327) );
  INVXL U21514 ( .A(n19655), .Y(n19323) );
  AOI21XL U21515 ( .A0(n19328), .A1(n19320), .B0(n19319), .Y(n19324) );
  INVXL U21516 ( .A(n19647), .Y(n19312) );
  NAND2XL U21517 ( .A(n19306), .B(n19305), .Y(n19307) );
  NAND2XL U21518 ( .A(n14824), .B(n19297), .Y(n19298) );
  XOR2XL U21519 ( .A(n19295), .B(n19294), .Y(n19296) );
  NAND2XL U21520 ( .A(n19293), .B(n19292), .Y(n19294) );
  XOR2XL U21521 ( .A(n19289), .B(n19288), .Y(n19290) );
  MXI2XL U21522 ( .A(U1_pipe4[0]), .B(n17049), .S0(n5804), .Y(n5068) );
  MXI2XL U21523 ( .A(U1_pipe4[1]), .B(n17048), .S0(n5804), .Y(n5069) );
  MXI2XL U21524 ( .A(U1_pipe4[2]), .B(n17045), .S0(n5804), .Y(n5070) );
  MXI2XL U21525 ( .A(U1_pipe4[3]), .B(n17042), .S0(n5804), .Y(n5071) );
  XOR2XL U21526 ( .A(n17041), .B(n17040), .Y(n17042) );
  MXI2XL U21527 ( .A(U1_pipe4[4]), .B(n17039), .S0(n5804), .Y(n5072) );
  XNOR2XL U21528 ( .A(n17038), .B(n17037), .Y(n17039) );
  MXI2XL U21529 ( .A(U1_pipe4[5]), .B(n17033), .S0(n5804), .Y(n5073) );
  XNOR2XL U21530 ( .A(n17031), .B(n17030), .Y(n17033) );
  MXI2XL U21531 ( .A(U1_pipe4[6]), .B(n17029), .S0(n5812), .Y(n5074) );
  XOR2XL U21532 ( .A(n17028), .B(n17027), .Y(n17029) );
  AOI21XL U21533 ( .A0(n17031), .A1(n17026), .B0(n17025), .Y(n17028) );
  INVXL U21534 ( .A(n17024), .Y(n17025) );
  MXI2XL U21535 ( .A(U1_pipe4[7]), .B(n17023), .S0(n7095), .Y(n5075) );
  XOR2XL U21536 ( .A(n17022), .B(n17021), .Y(n17023) );
  MXI2XL U21537 ( .A(U1_pipe4[8]), .B(n17017), .S0(n5812), .Y(n5076) );
  XOR2XL U21538 ( .A(n17016), .B(n17015), .Y(n17017) );
  XNOR2XL U21539 ( .A(n17013), .B(n17012), .Y(n17014) );
  XOR2XL U21540 ( .A(n17010), .B(n17009), .Y(n17011) );
  AOI21XL U21541 ( .A0(n17013), .A1(n17008), .B0(n17007), .Y(n17010) );
  INVXL U21542 ( .A(n17006), .Y(n17007) );
  MXI2XL U21543 ( .A(U1_pipe4[11]), .B(n17003), .S0(U1_valid[0]), .Y(n5079) );
  XNOR2XL U21544 ( .A(n17002), .B(n17001), .Y(n17003) );
  MXI2XL U21545 ( .A(U1_pipe4[12]), .B(n17000), .S0(U1_valid[0]), .Y(n5080) );
  XOR2XL U21546 ( .A(n16999), .B(n16998), .Y(n17000) );
  MXI2XL U21547 ( .A(U1_pipe4[13]), .B(n16994), .S0(U1_valid[0]), .Y(n5081) );
  XNOR2XL U21548 ( .A(n16993), .B(n16992), .Y(n16994) );
  MXI2XL U21549 ( .A(U1_pipe4[14]), .B(n16991), .S0(U1_valid[0]), .Y(n5082) );
  XOR2XL U21550 ( .A(n16990), .B(n16989), .Y(n16991) );
  AOI21XL U21551 ( .A0(n16993), .A1(n16988), .B0(n16987), .Y(n16990) );
  MXI2XL U21552 ( .A(U1_pipe4[15]), .B(n16986), .S0(U1_valid[0]), .Y(n5083) );
  XOR2XL U21553 ( .A(n16985), .B(n16984), .Y(n16986) );
  MXI2XL U21554 ( .A(U1_pipe4[16]), .B(n16983), .S0(U1_valid[0]), .Y(n5084) );
  MXI2XL U21555 ( .A(U1_pipe4[17]), .B(n16974), .S0(U1_valid[0]), .Y(n5085) );
  XOR2XL U21556 ( .A(n16969), .B(n16973), .Y(n16974) );
  MXI2XL U21557 ( .A(U1_pipe4[18]), .B(n16972), .S0(U1_valid[0]), .Y(n5086) );
  XNOR2XL U21558 ( .A(n16963), .B(n16962), .Y(n16964) );
  XOR2XL U21559 ( .A(n16942), .B(n16941), .Y(n16943) );
  MXI2XL U21560 ( .A(U1_pipe5[0]), .B(n17166), .S0(n17187), .Y(n5096) );
  MXI2XL U21561 ( .A(U1_pipe5[1]), .B(n17165), .S0(n5804), .Y(n5097) );
  MXI2XL U21562 ( .A(U1_pipe5[2]), .B(n17162), .S0(n5804), .Y(n5098) );
  MXI2XL U21563 ( .A(U1_pipe5[3]), .B(n17159), .S0(n5804), .Y(n5099) );
  XOR2XL U21564 ( .A(n17158), .B(n17157), .Y(n17159) );
  MXI2XL U21565 ( .A(U1_pipe5[4]), .B(n17156), .S0(n5804), .Y(n5100) );
  MXI2XL U21566 ( .A(U1_pipe5[5]), .B(n17150), .S0(n5804), .Y(n5101) );
  XNOR2XL U21567 ( .A(n17149), .B(n17148), .Y(n17150) );
  NAND2XL U21568 ( .A(n17147), .B(n17146), .Y(n17148) );
  MXI2XL U21569 ( .A(U1_pipe5[6]), .B(n17145), .S0(n5804), .Y(n5102) );
  XOR2XL U21570 ( .A(n17144), .B(n17143), .Y(n17145) );
  NAND2XL U21571 ( .A(n17142), .B(n17141), .Y(n17143) );
  AOI21XL U21572 ( .A0(n17149), .A1(n17147), .B0(n17139), .Y(n17144) );
  MXI2XL U21573 ( .A(U1_pipe5[7]), .B(n17137), .S0(n5804), .Y(n5103) );
  XOR2XL U21574 ( .A(n17136), .B(n17135), .Y(n17137) );
  NAND2XL U21575 ( .A(n13801), .B(n17134), .Y(n17135) );
  MXI2XL U21576 ( .A(U1_pipe5[8]), .B(n17130), .S0(n5804), .Y(n5104) );
  XOR2XL U21577 ( .A(n17129), .B(n17128), .Y(n17130) );
  XNOR2XL U21578 ( .A(n17126), .B(n17125), .Y(n17127) );
  XOR2XL U21579 ( .A(n17123), .B(n17122), .Y(n17124) );
  AOI21XL U21580 ( .A0(n17126), .A1(n17121), .B0(n17120), .Y(n17123) );
  MXI2XL U21581 ( .A(U1_pipe0[3]), .B(n19497), .S0(n19405), .Y(n5107) );
  XOR2XL U21582 ( .A(n19496), .B(n19495), .Y(n19497) );
  MXI2XL U21583 ( .A(U1_pipe0[5]), .B(n19488), .S0(n19215), .Y(n5108) );
  XOR2XL U21584 ( .A(n19484), .B(n19483), .Y(n19485) );
  AOI21XL U21585 ( .A0(n19487), .A1(n19482), .B0(n19481), .Y(n19484) );
  INVXL U21586 ( .A(n19480), .Y(n19481) );
  XOR2XL U21587 ( .A(n19478), .B(n19477), .Y(n19479) );
  XOR2XL U21588 ( .A(n19472), .B(n19471), .Y(n19473) );
  XNOR2XL U21589 ( .A(n19469), .B(n19468), .Y(n19470) );
  XOR2XL U21590 ( .A(n19466), .B(n19465), .Y(n19467) );
  AOI21XL U21591 ( .A0(n19469), .A1(n19464), .B0(n19463), .Y(n19466) );
  XNOR2XL U21592 ( .A(n19458), .B(n19457), .Y(n19459) );
  XOR2XL U21593 ( .A(n19455), .B(n19454), .Y(n19456) );
  XNOR2XL U21594 ( .A(n7685), .B(n19448), .Y(n19449) );
  XOR2XL U21595 ( .A(n19446), .B(n19445), .Y(n19447) );
  XOR2XL U21596 ( .A(n19441), .B(n19440), .Y(n19442) );
  XNOR2XL U21597 ( .A(n19429), .B(n19428), .Y(n19430) );
  XNOR2X1 U21598 ( .A(n19417), .B(n19416), .Y(n19418) );
  XOR2XL U21599 ( .A(n19404), .B(n19403), .Y(n19406) );
  XNOR2XL U21600 ( .A(n19396), .B(n19395), .Y(n19397) );
  MXI2XL U21601 ( .A(U1_pipe1[0]), .B(n19701), .S0(n25330), .Y(n5131) );
  MXI2XL U21602 ( .A(U1_pipe1[1]), .B(n19700), .S0(n25330), .Y(n5132) );
  MXI2XL U21603 ( .A(U1_pipe1[2]), .B(n19697), .S0(n25330), .Y(n5133) );
  MXI2XL U21604 ( .A(U1_pipe1[3]), .B(n19692), .S0(n25330), .Y(n5134) );
  XOR2XL U21605 ( .A(n19691), .B(n19690), .Y(n19692) );
  MXI2XL U21606 ( .A(U1_pipe1[4]), .B(n19689), .S0(n25330), .Y(n5135) );
  XNOR2XL U21607 ( .A(n19688), .B(n19687), .Y(n19689) );
  MXI2XL U21608 ( .A(U1_pipe1[5]), .B(n19683), .S0(n25330), .Y(n5136) );
  XNOR2XL U21609 ( .A(n19682), .B(n19681), .Y(n19683) );
  NAND2XL U21610 ( .A(n19680), .B(n19679), .Y(n19681) );
  MXI2XL U21611 ( .A(U1_pipe1[6]), .B(n19678), .S0(n25330), .Y(n5137) );
  XOR2XL U21612 ( .A(n19677), .B(n19676), .Y(n19678) );
  NAND2XL U21613 ( .A(n19675), .B(n19674), .Y(n19676) );
  AOI21XL U21614 ( .A0(n19682), .A1(n19680), .B0(n19672), .Y(n19677) );
  MXI2XL U21615 ( .A(U1_pipe1[7]), .B(n19670), .S0(n25330), .Y(n5138) );
  XOR2XL U21616 ( .A(n19669), .B(n19668), .Y(n19670) );
  NAND2XL U21617 ( .A(n19505), .B(n19667), .Y(n19668) );
  MXI2XL U21618 ( .A(U1_pipe1[8]), .B(n19663), .S0(n25330), .Y(n5139) );
  MXI2XL U21619 ( .A(U1_pipe1[9]), .B(n19660), .S0(n25330), .Y(n5140) );
  XNOR2XL U21620 ( .A(n19659), .B(n19658), .Y(n19660) );
  MXI2XL U21621 ( .A(U1_pipe1[10]), .B(n19657), .S0(n25330), .Y(n5141) );
  XOR2XL U21622 ( .A(n19656), .B(n19655), .Y(n19657) );
  AOI21XL U21623 ( .A0(n19659), .A1(n19654), .B0(n19653), .Y(n19656) );
  INVXL U21624 ( .A(n19652), .Y(n19653) );
  XNOR2XL U21625 ( .A(n19648), .B(n19647), .Y(n19649) );
  NAND2XL U21626 ( .A(n5788), .B(n19643), .Y(n19644) );
  XOR2XL U21627 ( .A(n19633), .B(n19632), .Y(n19634) );
  AOI21XL U21628 ( .A0(n19540), .A1(n19637), .B0(n19629), .Y(n19633) );
  MXI2XL U21629 ( .A(U1_pipe1[19]), .B(n19608), .S0(n25330), .Y(n5150) );
  MXI2XL U21630 ( .A(U1_pipe0[4]), .B(n19494), .S0(n19215), .Y(n5155) );
  XNOR2XL U21631 ( .A(n19493), .B(n19492), .Y(n19494) );
  AOI22XL U21632 ( .A0(in_valid), .A1(D_im[0]), .B0(buffer[0]), .B1(n29099), 
        .Y(n5157) );
  AOI22XL U21633 ( .A0(in_valid), .A1(D_im[1]), .B0(buffer[1]), .B1(n29099), 
        .Y(n5158) );
  AOI22XL U21634 ( .A0(in_valid), .A1(D_im[2]), .B0(buffer[2]), .B1(n11971), 
        .Y(n5159) );
  AOI22XL U21635 ( .A0(in_valid), .A1(D_im[3]), .B0(buffer[3]), .B1(n29099), 
        .Y(n5160) );
  AOI22XL U21636 ( .A0(in_valid), .A1(D_im[4]), .B0(buffer[4]), .B1(n11971), 
        .Y(n5161) );
  AOI22XL U21637 ( .A0(in_valid), .A1(D_im[5]), .B0(buffer[5]), .B1(n11971), 
        .Y(n5162) );
  AOI22XL U21638 ( .A0(in_valid), .A1(D_im[6]), .B0(buffer[6]), .B1(n11971), 
        .Y(n5163) );
  AOI22XL U21639 ( .A0(in_valid), .A1(D_im[7]), .B0(buffer[7]), .B1(n11971), 
        .Y(n5164) );
  AOI22XL U21640 ( .A0(in_valid), .A1(D_im[8]), .B0(buffer[8]), .B1(n29099), 
        .Y(n5165) );
  AOI22XL U21641 ( .A0(in_valid), .A1(D_im[9]), .B0(buffer[9]), .B1(n11971), 
        .Y(n5166) );
  AOI22XL U21642 ( .A0(in_valid), .A1(D_im[10]), .B0(buffer[10]), .B1(n11971), 
        .Y(n5167) );
  AOI22XL U21643 ( .A0(in_valid), .A1(D_im[11]), .B0(buffer[11]), .B1(n11971), 
        .Y(n5168) );
  AOI22XL U21644 ( .A0(in_valid), .A1(D_im[12]), .B0(buffer[12]), .B1(n11971), 
        .Y(n5169) );
  AOI22XL U21645 ( .A0(in_valid), .A1(D_im[13]), .B0(buffer[13]), .B1(n11971), 
        .Y(n5170) );
  AOI22XL U21646 ( .A0(in_valid), .A1(D_im[14]), .B0(buffer[14]), .B1(n11971), 
        .Y(n5171) );
  AOI22XL U21647 ( .A0(in_valid), .A1(D_im[15]), .B0(buffer[15]), .B1(n29099), 
        .Y(n5172) );
  AOI22XL U21648 ( .A0(in_valid), .A1(D_re[0]), .B0(buffer[16]), .B1(n11971), 
        .Y(n5173) );
  AOI22XL U21649 ( .A0(in_valid), .A1(D_re[1]), .B0(buffer[17]), .B1(n11971), 
        .Y(n5174) );
  AOI22XL U21650 ( .A0(in_valid), .A1(D_re[2]), .B0(buffer[18]), .B1(n11971), 
        .Y(n5175) );
  AOI22XL U21651 ( .A0(in_valid), .A1(D_re[3]), .B0(buffer[19]), .B1(n29099), 
        .Y(n5176) );
  AOI22XL U21652 ( .A0(in_valid), .A1(D_re[4]), .B0(buffer[20]), .B1(n11971), 
        .Y(n5177) );
  AOI22XL U21653 ( .A0(in_valid), .A1(D_re[5]), .B0(buffer[21]), .B1(n29099), 
        .Y(n5178) );
  AOI22XL U21654 ( .A0(in_valid), .A1(D_re[6]), .B0(buffer[22]), .B1(n11971), 
        .Y(n5179) );
  AOI22XL U21655 ( .A0(in_valid), .A1(D_re[7]), .B0(buffer[23]), .B1(n11971), 
        .Y(n5180) );
  AOI22XL U21656 ( .A0(in_valid), .A1(D_re[8]), .B0(buffer[24]), .B1(n11971), 
        .Y(n5181) );
  AOI22XL U21657 ( .A0(in_valid), .A1(D_re[9]), .B0(buffer[25]), .B1(n11971), 
        .Y(n5182) );
  AOI22XL U21658 ( .A0(in_valid), .A1(D_re[10]), .B0(buffer[26]), .B1(n11971), 
        .Y(n5183) );
  AOI22XL U21659 ( .A0(in_valid), .A1(D_re[11]), .B0(buffer[27]), .B1(n11971), 
        .Y(n5184) );
  AOI22XL U21660 ( .A0(in_valid), .A1(D_re[12]), .B0(buffer[28]), .B1(n29099), 
        .Y(n5185) );
  AOI22XL U21661 ( .A0(in_valid), .A1(D_re[13]), .B0(buffer[29]), .B1(n11971), 
        .Y(n5186) );
  AOI22XL U21662 ( .A0(in_valid), .A1(D_re[14]), .B0(buffer[30]), .B1(n11971), 
        .Y(n5187) );
  AOI22XL U21663 ( .A0(in_valid), .A1(D_re[15]), .B0(buffer[31]), .B1(n11971), 
        .Y(n5188) );
  AOI22XL U21664 ( .A0(B5_q[0]), .A1(n11864), .B0(B6_q[0]), .B1(n5801), .Y(
        n11718) );
  AOI22XL U21665 ( .A0(B4_q[0]), .A1(n5802), .B0(B0_q[0]), .B1(n5828), .Y(
        n11717) );
  AOI22XL U21666 ( .A0(B2_q[0]), .A1(n5831), .B0(B1_q[0]), .B1(n5832), .Y(
        n11716) );
  AOI22XL U21667 ( .A0(B7_q[10]), .A1(n5803), .B0(B0_q[10]), .B1(n5828), .Y(
        n11727) );
  AOI22XL U21668 ( .A0(B4_q[10]), .A1(n5802), .B0(B2_q[10]), .B1(n5831), .Y(
        n11726) );
  AOI22XL U21669 ( .A0(B6_q[10]), .A1(n5801), .B0(B3_q[10]), .B1(n5833), .Y(
        n11725) );
  AOI22XL U21670 ( .A0(B4_q[11]), .A1(n5802), .B0(B6_q[11]), .B1(n5801), .Y(
        n11791) );
  AOI22XL U21671 ( .A0(B5_q[11]), .A1(n11864), .B0(B1_q[11]), .B1(n5832), .Y(
        n11790) );
  AOI22XL U21672 ( .A0(B7_q[11]), .A1(n5803), .B0(B2_q[11]), .B1(n5831), .Y(
        n11789) );
  AOI22XL U21673 ( .A0(B6_q[12]), .A1(n5801), .B0(B1_q[12]), .B1(n5832), .Y(
        n11835) );
  AOI22XL U21674 ( .A0(B4_q[12]), .A1(n5802), .B0(B3_q[12]), .B1(n5833), .Y(
        n11834) );
  AOI22XL U21675 ( .A0(B7_q[12]), .A1(n5803), .B0(B2_q[12]), .B1(n5831), .Y(
        n11833) );
  AOI22XL U21676 ( .A0(B0_q[13]), .A1(n5828), .B0(B3_q[13]), .B1(n5833), .Y(
        n11743) );
  AOI22XL U21677 ( .A0(B1_q[13]), .A1(n5832), .B0(B2_q[13]), .B1(n5831), .Y(
        n11742) );
  AOI22XL U21678 ( .A0(B4_q[13]), .A1(n5802), .B0(B7_q[13]), .B1(n5803), .Y(
        n11741) );
  AOI22XL U21679 ( .A0(B4_q[14]), .A1(n5802), .B0(B2_q[14]), .B1(n5831), .Y(
        n11714) );
  AOI22XL U21680 ( .A0(B7_q[14]), .A1(n5803), .B0(B0_q[14]), .B1(n5828), .Y(
        n11713) );
  AOI22XL U21681 ( .A0(B5_q[14]), .A1(n11864), .B0(B6_q[14]), .B1(n5801), .Y(
        n11712) );
  AOI22XL U21682 ( .A0(B5_q[15]), .A1(n11676), .B0(B4_q[15]), .B1(n5802), .Y(
        n11872) );
  AOI22XL U21683 ( .A0(B3_q[15]), .A1(n5833), .B0(B1_q[15]), .B1(n5832), .Y(
        n11871) );
  AOI22XL U21684 ( .A0(B6_q[15]), .A1(n5801), .B0(B2_q[15]), .B1(n5831), .Y(
        n11870) );
  AOI22XL U21685 ( .A0(B4_q[16]), .A1(n5802), .B0(B1_q[16]), .B1(n5832), .Y(
        n11868) );
  AOI22XL U21686 ( .A0(B5_q[16]), .A1(n11864), .B0(B3_q[16]), .B1(n5833), .Y(
        n11867) );
  AOI22XL U21687 ( .A0(B7_q[16]), .A1(n5803), .B0(B2_q[16]), .B1(n5831), .Y(
        n11866) );
  AOI22XL U21688 ( .A0(B6_q[17]), .A1(n5801), .B0(B3_q[17]), .B1(n5833), .Y(
        n11803) );
  AOI22XL U21689 ( .A0(B7_q[17]), .A1(n5803), .B0(B2_q[17]), .B1(n5831), .Y(
        n11802) );
  AOI22XL U21690 ( .A0(B5_q[17]), .A1(n11676), .B0(B4_q[17]), .B1(n5802), .Y(
        n11801) );
  AOI22XL U21691 ( .A0(B4_q[18]), .A1(n5802), .B0(B3_q[18]), .B1(n5833), .Y(
        n11863) );
  AOI22XL U21692 ( .A0(B5_q[18]), .A1(n11864), .B0(B2_q[18]), .B1(n5831), .Y(
        n11862) );
  AOI22XL U21693 ( .A0(B6_q[18]), .A1(n5801), .B0(B0_q[18]), .B1(n5828), .Y(
        n11861) );
  AOI22XL U21694 ( .A0(B4_q[19]), .A1(n5802), .B0(B0_q[19]), .B1(n5828), .Y(
        n11815) );
  AOI22XL U21695 ( .A0(B5_q[19]), .A1(n11864), .B0(B1_q[19]), .B1(n5832), .Y(
        n11814) );
  AOI22XL U21696 ( .A0(B3_q[19]), .A1(n5833), .B0(B2_q[19]), .B1(n5831), .Y(
        n11813) );
  AOI22XL U21697 ( .A0(B5_q[1]), .A1(n11864), .B0(B0_q[1]), .B1(n5828), .Y(
        n11671) );
  AOI22XL U21698 ( .A0(B7_q[1]), .A1(n5803), .B0(B6_q[1]), .B1(n5801), .Y(
        n11670) );
  AOI22XL U21699 ( .A0(B3_q[1]), .A1(n5833), .B0(B2_q[1]), .B1(n5831), .Y(
        n11669) );
  AOI22XL U21700 ( .A0(B2_q[20]), .A1(n5831), .B0(B1_q[20]), .B1(n5832), .Y(
        n11843) );
  AOI22XL U21701 ( .A0(B7_q[20]), .A1(n5803), .B0(B0_q[20]), .B1(n5828), .Y(
        n11842) );
  AOI22XL U21702 ( .A0(B4_q[20]), .A1(n5802), .B0(B5_q[20]), .B1(n11676), .Y(
        n11841) );
  AOI22XL U21703 ( .A0(B7_q[21]), .A1(n5803), .B0(B1_q[21]), .B1(n5832), .Y(
        n11811) );
  AOI22XL U21704 ( .A0(B5_q[21]), .A1(n11864), .B0(B3_q[21]), .B1(n5833), .Y(
        n11810) );
  AOI22XL U21705 ( .A0(B4_q[21]), .A1(n5802), .B0(B6_q[21]), .B1(n5801), .Y(
        n11809) );
  AND4XL U21706 ( .A(n11723), .B(n11722), .C(n11721), .D(n11720), .Y(n5217) );
  AOI22XL U21707 ( .A0(B6_q[22]), .A1(n5801), .B0(B2_q[22]), .B1(n5831), .Y(
        n11723) );
  AOI22XL U21708 ( .A0(B0_q[22]), .A1(n5828), .B0(B3_q[22]), .B1(n5833), .Y(
        n11722) );
  AOI22XL U21709 ( .A0(B4_q[22]), .A1(n5802), .B0(B5_q[22]), .B1(n11676), .Y(
        n11721) );
  AOI22XL U21710 ( .A0(B5_q[23]), .A1(n11676), .B0(B3_q[23]), .B1(n5833), .Y(
        n11807) );
  AOI22XL U21711 ( .A0(B4_q[23]), .A1(n5802), .B0(B1_q[23]), .B1(n5832), .Y(
        n11806) );
  AOI22XL U21712 ( .A0(B6_q[23]), .A1(n5801), .B0(B7_q[23]), .B1(n5803), .Y(
        n11805) );
  AOI22XL U21713 ( .A0(B5_q[24]), .A1(n11676), .B0(B2_q[24]), .B1(n5831), .Y(
        n11839) );
  AOI22XL U21714 ( .A0(B7_q[24]), .A1(n5803), .B0(B6_q[24]), .B1(n5801), .Y(
        n11838) );
  AOI22XL U21715 ( .A0(B4_q[24]), .A1(n5802), .B0(B1_q[24]), .B1(n5832), .Y(
        n11837) );
  AOI22XL U21716 ( .A0(B6_q[25]), .A1(n5801), .B0(B3_q[25]), .B1(n5833), .Y(
        n11783) );
  AOI22XL U21717 ( .A0(B5_q[25]), .A1(n11676), .B0(B4_q[25]), .B1(n5802), .Y(
        n11782) );
  AOI22XL U21718 ( .A0(B7_q[25]), .A1(n5803), .B0(B0_q[25]), .B1(n5828), .Y(
        n11781) );
  AOI22XL U21719 ( .A0(B5_q[26]), .A1(n11676), .B0(B1_q[26]), .B1(n5832), .Y(
        n11859) );
  AOI22XL U21720 ( .A0(B2_q[26]), .A1(n5831), .B0(B3_q[26]), .B1(n5833), .Y(
        n11858) );
  AOI22XL U21721 ( .A0(B7_q[26]), .A1(n5803), .B0(B0_q[26]), .B1(n5828), .Y(
        n11857) );
  AOI22XL U21722 ( .A0(B5_q[27]), .A1(n11676), .B0(B2_q[27]), .B1(n5831), .Y(
        n11739) );
  AOI22XL U21723 ( .A0(B6_q[27]), .A1(n5801), .B0(B0_q[27]), .B1(n5828), .Y(
        n11738) );
  AOI22XL U21724 ( .A0(B7_q[27]), .A1(n5803), .B0(B3_q[27]), .B1(n5833), .Y(
        n11737) );
  AOI22XL U21725 ( .A0(B7_q[28]), .A1(n5803), .B0(B0_q[28]), .B1(n5828), .Y(
        n11688) );
  AOI22XL U21726 ( .A0(B2_q[28]), .A1(n5831), .B0(B1_q[28]), .B1(n5832), .Y(
        n11687) );
  AOI22XL U21727 ( .A0(B6_q[28]), .A1(n5801), .B0(B5_q[28]), .B1(n11676), .Y(
        n11686) );
  AOI22XL U21728 ( .A0(B7_q[29]), .A1(n5803), .B0(B2_q[29]), .B1(n5831), .Y(
        n11696) );
  AOI22XL U21729 ( .A0(B6_q[29]), .A1(n5801), .B0(B1_q[29]), .B1(n5832), .Y(
        n11695) );
  AOI22XL U21730 ( .A0(B5_q[29]), .A1(n11676), .B0(B3_q[29]), .B1(n5833), .Y(
        n11694) );
  AOI22XL U21731 ( .A0(B7_q[2]), .A1(n5803), .B0(B5_q[2]), .B1(n11676), .Y(
        n11779) );
  AOI22XL U21732 ( .A0(B4_q[2]), .A1(n5802), .B0(B3_q[2]), .B1(n5833), .Y(
        n11778) );
  AOI22XL U21733 ( .A0(B6_q[2]), .A1(n5801), .B0(B2_q[2]), .B1(n5831), .Y(
        n11777) );
  AOI22XL U21734 ( .A0(B7_q[30]), .A1(n5803), .B0(B3_q[30]), .B1(n5833), .Y(
        n11795) );
  AOI22XL U21735 ( .A0(B4_q[30]), .A1(n5802), .B0(B1_q[30]), .B1(n5832), .Y(
        n11794) );
  AOI22XL U21736 ( .A0(B5_q[30]), .A1(n11676), .B0(B6_q[30]), .B1(n5801), .Y(
        n11793) );
  AOI22XL U21737 ( .A0(B7_q[31]), .A1(n5803), .B0(B3_q[31]), .B1(n5833), .Y(
        n11759) );
  AOI22XL U21738 ( .A0(B6_q[31]), .A1(n5801), .B0(B1_q[31]), .B1(n5832), .Y(
        n11758) );
  AOI22XL U21739 ( .A0(B4_q[31]), .A1(n5802), .B0(B2_q[31]), .B1(n5831), .Y(
        n11757) );
  AOI22XL U21740 ( .A0(B3_q[32]), .A1(n5833), .B0(B2_q[32]), .B1(n5831), .Y(
        n11747) );
  AOI22XL U21741 ( .A0(B6_q[32]), .A1(n5801), .B0(B1_q[32]), .B1(n5832), .Y(
        n11746) );
  AOI22XL U21742 ( .A0(B5_q[32]), .A1(n11676), .B0(B0_q[32]), .B1(n5828), .Y(
        n11745) );
  AOI22XL U21743 ( .A0(B5_q[33]), .A1(n11676), .B0(B3_q[33]), .B1(n5833), .Y(
        n11683) );
  AOI22XL U21744 ( .A0(B6_q[33]), .A1(n5801), .B0(B0_q[33]), .B1(n5828), .Y(
        n11682) );
  AOI22XL U21745 ( .A0(B4_q[33]), .A1(n5802), .B0(B2_q[33]), .B1(n5831), .Y(
        n11681) );
  AOI22XL U21746 ( .A0(B1_q[34]), .A1(n5832), .B0(B3_q[34]), .B1(n5833), .Y(
        n11731) );
  AOI22XL U21747 ( .A0(B4_q[34]), .A1(n5802), .B0(B0_q[34]), .B1(n5828), .Y(
        n11730) );
  AOI22XL U21748 ( .A0(B7_q[34]), .A1(n5803), .B0(B2_q[34]), .B1(n5831), .Y(
        n11729) );
  AOI22XL U21749 ( .A0(B7_q[35]), .A1(n5803), .B0(B4_q[35]), .B1(n5802), .Y(
        n11847) );
  AOI22XL U21750 ( .A0(B1_q[35]), .A1(n5832), .B0(B3_q[35]), .B1(n5833), .Y(
        n11846) );
  AOI22XL U21751 ( .A0(B6_q[35]), .A1(n5801), .B0(B0_q[35]), .B1(n5828), .Y(
        n11845) );
  AND4XL U21752 ( .A(n11819), .B(n11818), .C(n11817), .D(n11816), .Y(n5247) );
  AOI22XL U21753 ( .A0(B6_q[36]), .A1(n5801), .B0(B0_q[36]), .B1(n5828), .Y(
        n11819) );
  AOI22XL U21754 ( .A0(B2_q[36]), .A1(n5831), .B0(B3_q[36]), .B1(n5833), .Y(
        n11818) );
  AOI22XL U21755 ( .A0(B5_q[36]), .A1(n11676), .B0(B7_q[36]), .B1(n5803), .Y(
        n11817) );
  AOI22XL U21756 ( .A0(B5_q[37]), .A1(n11676), .B0(B4_q[37]), .B1(n5802), .Y(
        n11767) );
  AOI22XL U21757 ( .A0(B6_q[37]), .A1(n5801), .B0(B2_q[37]), .B1(n5831), .Y(
        n11766) );
  AOI22XL U21758 ( .A0(B0_q[37]), .A1(n5828), .B0(B3_q[37]), .B1(n5833), .Y(
        n11765) );
  AOI22XL U21759 ( .A0(B4_q[38]), .A1(n5802), .B0(B6_q[38]), .B1(n5801), .Y(
        n11751) );
  AOI22XL U21760 ( .A0(B2_q[38]), .A1(n5831), .B0(B1_q[38]), .B1(n5832), .Y(
        n11750) );
  AOI22XL U21761 ( .A0(B5_q[38]), .A1(n11864), .B0(B0_q[38]), .B1(n5828), .Y(
        n11749) );
  AOI22XL U21762 ( .A0(B7_q[39]), .A1(n5803), .B0(B2_q[39]), .B1(n5831), .Y(
        n11675) );
  AOI22XL U21763 ( .A0(B4_q[39]), .A1(n5802), .B0(B6_q[39]), .B1(n5801), .Y(
        n11674) );
  AOI22XL U21764 ( .A0(B5_q[39]), .A1(n11864), .B0(B0_q[39]), .B1(n5828), .Y(
        n11673) );
  AOI22XL U21765 ( .A0(B4_q[3]), .A1(n5802), .B0(B0_q[3]), .B1(n5828), .Y(
        n11827) );
  AOI22XL U21766 ( .A0(B1_q[3]), .A1(n5832), .B0(B3_q[3]), .B1(n5833), .Y(
        n11826) );
  AOI22XL U21767 ( .A0(B7_q[3]), .A1(n5803), .B0(B2_q[3]), .B1(n5831), .Y(
        n11825) );
  AOI22XL U21768 ( .A0(B5_q[40]), .A1(n11676), .B0(B6_q[40]), .B1(n5801), .Y(
        n11787) );
  AOI22XL U21769 ( .A0(B2_q[40]), .A1(n5831), .B0(B1_q[40]), .B1(n5832), .Y(
        n11786) );
  AOI22XL U21770 ( .A0(B4_q[40]), .A1(n5802), .B0(B3_q[40]), .B1(n5833), .Y(
        n11785) );
  AOI22XL U21771 ( .A0(B5_q[41]), .A1(n11864), .B0(B0_q[41]), .B1(n5828), .Y(
        n11855) );
  AOI22XL U21772 ( .A0(B6_q[41]), .A1(n5801), .B0(B1_q[41]), .B1(n5832), .Y(
        n11854) );
  AOI22XL U21773 ( .A0(B7_q[41]), .A1(n5803), .B0(B3_q[41]), .B1(n5833), .Y(
        n11853) );
  AOI22XL U21774 ( .A0(B2_q[42]), .A1(n5831), .B0(B3_q[42]), .B1(n5833), .Y(
        n11663) );
  AOI22XL U21775 ( .A0(B6_q[42]), .A1(n5801), .B0(B7_q[42]), .B1(n5803), .Y(
        n11662) );
  AOI22XL U21776 ( .A0(B5_q[42]), .A1(n11864), .B0(B0_q[42]), .B1(n5828), .Y(
        n11661) );
  AOI22XL U21777 ( .A0(B6_q[43]), .A1(n5801), .B0(B3_q[43]), .B1(n5833), .Y(
        n11823) );
  AOI22XL U21778 ( .A0(B5_q[43]), .A1(n11864), .B0(B7_q[43]), .B1(n5803), .Y(
        n11822) );
  AOI22XL U21779 ( .A0(B4_q[43]), .A1(n5802), .B0(B2_q[43]), .B1(n5831), .Y(
        n11821) );
  AOI22XL U21780 ( .A0(B6_q[44]), .A1(n5801), .B0(B2_q[44]), .B1(n5831), .Y(
        n11763) );
  AOI22XL U21781 ( .A0(B5_q[44]), .A1(n11864), .B0(B7_q[44]), .B1(n5803), .Y(
        n11762) );
  AOI22XL U21782 ( .A0(B4_q[44]), .A1(n5802), .B0(B1_q[44]), .B1(n5832), .Y(
        n11761) );
  AOI22XL U21783 ( .A0(B0_q[45]), .A1(n5828), .B0(B3_q[45]), .B1(n5833), .Y(
        n11704) );
  AOI22XL U21784 ( .A0(B5_q[45]), .A1(n11676), .B0(B6_q[45]), .B1(n5801), .Y(
        n11703) );
  AOI22XL U21785 ( .A0(B2_q[45]), .A1(n5831), .B0(B1_q[45]), .B1(n5832), .Y(
        n11702) );
  AOI22XL U21786 ( .A0(B7_q[46]), .A1(n5803), .B0(B3_q[46]), .B1(n5833), .Y(
        n11708) );
  AOI22XL U21787 ( .A0(B4_q[46]), .A1(n5802), .B0(B2_q[46]), .B1(n5831), .Y(
        n11707) );
  AOI22XL U21788 ( .A0(B5_q[46]), .A1(n11864), .B0(B0_q[46]), .B1(n5828), .Y(
        n11706) );
  AOI22XL U21789 ( .A0(B7_q[47]), .A1(n5803), .B0(B0_q[47]), .B1(n5828), .Y(
        n11659) );
  AOI22XL U21790 ( .A0(B4_q[47]), .A1(n5802), .B0(B3_q[47]), .B1(n5833), .Y(
        n11658) );
  AOI22XL U21791 ( .A0(B6_q[47]), .A1(n5801), .B0(B2_q[47]), .B1(n5831), .Y(
        n11657) );
  AOI22XL U21792 ( .A0(B6_q[48]), .A1(n5801), .B0(B3_q[48]), .B1(n5833), .Y(
        n11692) );
  AOI22XL U21793 ( .A0(B4_q[48]), .A1(n5802), .B0(B2_q[48]), .B1(n5831), .Y(
        n11691) );
  AOI22XL U21794 ( .A0(B7_q[48]), .A1(n5803), .B0(B0_q[48]), .B1(n5828), .Y(
        n11690) );
  AOI22XL U21795 ( .A0(B0_q[49]), .A1(n5828), .B0(B3_q[49]), .B1(n5833), .Y(
        n11755) );
  AOI22XL U21796 ( .A0(B6_q[49]), .A1(n5801), .B0(B2_q[49]), .B1(n5831), .Y(
        n11754) );
  AOI22XL U21797 ( .A0(B4_q[49]), .A1(n5802), .B0(B1_q[49]), .B1(n5832), .Y(
        n11753) );
  AND4XL U21798 ( .A(n11735), .B(n11734), .C(n11733), .D(n11732), .Y(n5277) );
  AOI22XL U21799 ( .A0(B2_q[4]), .A1(n5831), .B0(B3_q[4]), .B1(n5833), .Y(
        n11735) );
  AOI22XL U21800 ( .A0(B4_q[4]), .A1(n5802), .B0(B1_q[4]), .B1(n5832), .Y(
        n11734) );
  AOI22XL U21801 ( .A0(B6_q[4]), .A1(n5801), .B0(B0_q[4]), .B1(n5828), .Y(
        n11733) );
  AOI22XL U21802 ( .A0(B6_q[50]), .A1(n5801), .B0(B7_q[50]), .B1(n5803), .Y(
        n11700) );
  AOI22XL U21803 ( .A0(B2_q[50]), .A1(n5831), .B0(B0_q[50]), .B1(n5828), .Y(
        n11699) );
  AOI22XL U21804 ( .A0(B4_q[50]), .A1(n5802), .B0(B3_q[50]), .B1(n5833), .Y(
        n11698) );
  AOI22XL U21805 ( .A0(B5_q[51]), .A1(n11676), .B0(B4_q[51]), .B1(n5802), .Y(
        n11771) );
  AOI22XL U21806 ( .A0(B2_q[51]), .A1(n5831), .B0(B1_q[51]), .B1(n5832), .Y(
        n11770) );
  AOI22XL U21807 ( .A0(B0_q[51]), .A1(n5828), .B0(B3_q[51]), .B1(n5833), .Y(
        n11769) );
  AOI22XL U21808 ( .A0(B6_q[5]), .A1(n5801), .B0(B3_q[5]), .B1(n5833), .Y(
        n11799) );
  AOI22XL U21809 ( .A0(B7_q[5]), .A1(n5803), .B0(B4_q[5]), .B1(n5802), .Y(
        n11798) );
  AOI22XL U21810 ( .A0(B5_q[5]), .A1(n11676), .B0(B1_q[5]), .B1(n5832), .Y(
        n11797) );
  AOI22XL U21811 ( .A0(B7_q[6]), .A1(n5803), .B0(B1_q[6]), .B1(n5832), .Y(
        n11851) );
  AOI22XL U21812 ( .A0(B5_q[6]), .A1(n11676), .B0(B2_q[6]), .B1(n5831), .Y(
        n11850) );
  AOI22XL U21813 ( .A0(B3_q[6]), .A1(n5833), .B0(B0_q[6]), .B1(n5828), .Y(
        n11849) );
  AOI22XL U21814 ( .A0(B6_q[7]), .A1(n5801), .B0(B3_q[7]), .B1(n5833), .Y(
        n11667) );
  AOI22XL U21815 ( .A0(B2_q[7]), .A1(n5831), .B0(B0_q[7]), .B1(n5828), .Y(
        n11666) );
  AOI22XL U21816 ( .A0(B7_q[7]), .A1(n5803), .B0(B4_q[7]), .B1(n5802), .Y(
        n11665) );
  AOI22XL U21817 ( .A0(B7_q[8]), .A1(n5803), .B0(B0_q[8]), .B1(n5828), .Y(
        n11775) );
  AOI22XL U21818 ( .A0(B4_q[8]), .A1(n5802), .B0(B3_q[8]), .B1(n5833), .Y(
        n11774) );
  AOI22XL U21819 ( .A0(B6_q[8]), .A1(n5801), .B0(B1_q[8]), .B1(n5832), .Y(
        n11773) );
  AOI22XL U21820 ( .A0(B6_q[9]), .A1(n5801), .B0(B7_q[9]), .B1(n5803), .Y(
        n11831) );
  AOI22XL U21821 ( .A0(B4_q[9]), .A1(n5802), .B0(B0_q[9]), .B1(n5828), .Y(
        n11830) );
  AOI22XL U21822 ( .A0(B5_q[9]), .A1(n11864), .B0(B3_q[9]), .B1(n5833), .Y(
        n11829) );
  AOI22XL U21823 ( .A0(n5834), .A1(Q2_addr[15]), .B0(Q2_addr[7]), .B1(n5830), 
        .Y(n5345) );
  AOI22XL U21824 ( .A0(n5911), .A1(Q2_addr[23]), .B0(Q2_addr[15]), .B1(n11958), 
        .Y(n5346) );
  AOI22XL U21825 ( .A0(n11956), .A1(Q2_addr[31]), .B0(Q2_addr[23]), .B1(n5808), 
        .Y(n5347) );
  AOI22XL U21826 ( .A0(n5834), .A1(Q2_addr[39]), .B0(Q2_addr[31]), .B1(n5830), 
        .Y(n5348) );
  AOI22XL U21827 ( .A0(n5834), .A1(Q3_addr[15]), .B0(Q3_addr[7]), .B1(n11958), 
        .Y(n5350) );
  AOI22XL U21828 ( .A0(n5834), .A1(Q3_addr[23]), .B0(Q3_addr[15]), .B1(n5830), 
        .Y(n5351) );
  AOI22XL U21829 ( .A0(n5834), .A1(Q3_addr[31]), .B0(Q3_addr[23]), .B1(n5808), 
        .Y(n5352) );
  AOI22XL U21830 ( .A0(n5834), .A1(Q3_addr[39]), .B0(Q3_addr[31]), .B1(n5808), 
        .Y(n5353) );
  AOI22XL U21831 ( .A0(n5834), .A1(Q2_addr[14]), .B0(Q2_addr[6]), .B1(n5808), 
        .Y(n5355) );
  AOI22XL U21832 ( .A0(n5834), .A1(Q2_addr[22]), .B0(Q2_addr[14]), .B1(n5808), 
        .Y(n5356) );
  AOI22XL U21833 ( .A0(n5834), .A1(Q2_addr[30]), .B0(Q2_addr[22]), .B1(n5808), 
        .Y(n5357) );
  AOI22XL U21834 ( .A0(n5834), .A1(Q2_addr[38]), .B0(Q2_addr[30]), .B1(n11954), 
        .Y(n5358) );
  AOI22XL U21835 ( .A0(n5834), .A1(Q0_addr[14]), .B0(Q0_addr[6]), .B1(n5808), 
        .Y(n5360) );
  AOI22XL U21836 ( .A0(n5834), .A1(Q0_addr[22]), .B0(Q0_addr[14]), .B1(n11954), 
        .Y(n5361) );
  AOI22XL U21837 ( .A0(n5911), .A1(Q0_addr[30]), .B0(Q0_addr[22]), .B1(n11957), 
        .Y(n5362) );
  AOI22XL U21838 ( .A0(n5911), .A1(Q0_addr[38]), .B0(Q0_addr[30]), .B1(n11954), 
        .Y(n5363) );
  AOI22XL U21839 ( .A0(n5911), .A1(Q2_addr[12]), .B0(Q2_addr[4]), .B1(n11958), 
        .Y(n5365) );
  AOI22XL U21840 ( .A0(n11956), .A1(Q2_addr[20]), .B0(Q2_addr[12]), .B1(n11954), .Y(n5366) );
  AOI22XL U21841 ( .A0(n5911), .A1(Q2_addr[28]), .B0(Q2_addr[20]), .B1(n11954), 
        .Y(n5367) );
  AOI22XL U21842 ( .A0(n11956), .A1(Q2_addr[36]), .B0(Q2_addr[28]), .B1(n5808), 
        .Y(n5368) );
  AOI22XL U21843 ( .A0(n5911), .A1(Q0_addr[12]), .B0(Q0_addr[4]), .B1(n11957), 
        .Y(n5370) );
  AOI22XL U21844 ( .A0(n11956), .A1(Q0_addr[20]), .B0(Q0_addr[12]), .B1(n5808), 
        .Y(n5371) );
  AOI22XL U21845 ( .A0(n5911), .A1(Q0_addr[28]), .B0(Q0_addr[20]), .B1(n11958), 
        .Y(n5372) );
  AOI22XL U21846 ( .A0(n11956), .A1(Q0_addr[36]), .B0(Q0_addr[28]), .B1(n5830), 
        .Y(n5373) );
  AOI22XL U21847 ( .A0(n5911), .A1(Q0_addr[13]), .B0(Q0_addr[5]), .B1(n5830), 
        .Y(n5375) );
  AOI22XL U21848 ( .A0(n5911), .A1(Q0_addr[21]), .B0(Q0_addr[13]), .B1(n5830), 
        .Y(n5376) );
  AOI22XL U21849 ( .A0(n5911), .A1(Q0_addr[29]), .B0(Q0_addr[21]), .B1(n5830), 
        .Y(n5377) );
  AOI22XL U21850 ( .A0(n11953), .A1(Q0_addr[37]), .B0(Q0_addr[29]), .B1(n11952), .Y(n5378) );
  AOI22XL U21851 ( .A0(n5911), .A1(Q1_addr[13]), .B0(Q1_addr[5]), .B1(n11952), 
        .Y(n5380) );
  AOI22XL U21852 ( .A0(n11956), .A1(Q1_addr[21]), .B0(Q1_addr[13]), .B1(n11957), .Y(n5381) );
  AOI22XL U21853 ( .A0(n5911), .A1(Q1_addr[29]), .B0(Q1_addr[21]), .B1(n5808), 
        .Y(n5382) );
  AOI22XL U21854 ( .A0(n11956), .A1(Q1_addr[37]), .B0(Q1_addr[29]), .B1(n5808), 
        .Y(n5383) );
  AOI22XL U21855 ( .A0(n5911), .A1(Q0_addr[15]), .B0(Q0_addr[7]), .B1(n5808), 
        .Y(n5385) );
  AOI22XL U21856 ( .A0(n11956), .A1(Q0_addr[23]), .B0(Q0_addr[15]), .B1(n5808), 
        .Y(n5386) );
  AOI22XL U21857 ( .A0(n5911), .A1(Q0_addr[31]), .B0(Q0_addr[23]), .B1(n5808), 
        .Y(n5387) );
  AOI22XL U21858 ( .A0(n11956), .A1(Q0_addr[39]), .B0(Q0_addr[31]), .B1(n5808), 
        .Y(n5388) );
  AOI22XL U21859 ( .A0(n5911), .A1(Q1_addr[15]), .B0(Q1_addr[7]), .B1(n5808), 
        .Y(n5390) );
  AOI22XL U21860 ( .A0(n11956), .A1(Q1_addr[23]), .B0(Q1_addr[15]), .B1(n5808), 
        .Y(n5391) );
  AOI22XL U21861 ( .A0(n5911), .A1(Q1_addr[31]), .B0(Q1_addr[23]), .B1(n11952), 
        .Y(n5392) );
  AOI22XL U21862 ( .A0(n11956), .A1(Q1_addr[39]), .B0(Q1_addr[31]), .B1(n5830), 
        .Y(n5393) );
  AOI22XL U21863 ( .A0(n5834), .A1(Q1_addr[14]), .B0(Q1_addr[6]), .B1(n11954), 
        .Y(n5395) );
  AOI22XL U21864 ( .A0(n5834), .A1(Q1_addr[22]), .B0(Q1_addr[14]), .B1(n11952), 
        .Y(n5396) );
  AOI22XL U21865 ( .A0(n11953), .A1(Q1_addr[30]), .B0(Q1_addr[22]), .B1(n11957), .Y(n5397) );
  AOI22XL U21866 ( .A0(n11953), .A1(Q1_addr[38]), .B0(Q1_addr[30]), .B1(n11957), .Y(n5398) );
  AOI22XL U21867 ( .A0(n11953), .A1(Q3_addr[14]), .B0(Q3_addr[6]), .B1(n11958), 
        .Y(n5400) );
  AOI22XL U21868 ( .A0(n11953), .A1(Q3_addr[22]), .B0(Q3_addr[14]), .B1(n11957), .Y(n5401) );
  AOI22XL U21869 ( .A0(n11953), .A1(Q3_addr[30]), .B0(Q3_addr[22]), .B1(n11957), .Y(n5402) );
  AOI22XL U21870 ( .A0(n11953), .A1(Q3_addr[38]), .B0(Q3_addr[30]), .B1(n11954), .Y(n5403) );
  AOI22XL U21871 ( .A0(n11997), .A1(C_sel_reg[1]), .B0(C_sel_reg[3]), .B1(
        n5829), .Y(n5407) );
  AOI22XL U21872 ( .A0(n11997), .A1(C_sel_reg[3]), .B0(C_sel_reg[5]), .B1(
        n5829), .Y(n5408) );
  AOI22XL U21873 ( .A0(n11997), .A1(C_sel_reg[5]), .B0(C_sel_reg[7]), .B1(
        n5829), .Y(n5409) );
  AOI22XL U21874 ( .A0(n11997), .A1(C_sel_reg[7]), .B0(C_sel_reg[9]), .B1(
        n5829), .Y(n5410) );
  AOI22XL U21875 ( .A0(n12000), .A1(C_sel_reg[9]), .B0(n11999), .B1(n5829), 
        .Y(n5411) );
  AOI22XL U21876 ( .A0(n12000), .A1(C_sel_reg[2]), .B0(C_sel_reg[4]), .B1(
        n5829), .Y(n5413) );
  AOI22XL U21877 ( .A0(n12000), .A1(C_sel_reg[4]), .B0(C_sel_reg[6]), .B1(
        n5829), .Y(n5414) );
  AOI22XL U21878 ( .A0(n12000), .A1(C_sel_reg[6]), .B0(C_sel_reg[8]), .B1(
        n5829), .Y(n5415) );
  AOI22XL U21879 ( .A0(n12000), .A1(A_sel_reg[1]), .B0(A_sel_reg[2]), .B1(
        n5829), .Y(n5418) );
  AOI22XL U21880 ( .A0(n12000), .A1(A_sel_reg[2]), .B0(A_sel_reg[3]), .B1(
        n5829), .Y(n5419) );
  AOI22XL U21881 ( .A0(n12000), .A1(A_sel_reg[3]), .B0(A_sel_reg[4]), .B1(
        n5829), .Y(n5420) );
  AOI22XL U21882 ( .A0(n12000), .A1(A_sel_reg[4]), .B0(n11998), .B1(n5829), 
        .Y(n5421) );
  AOI22XL U21883 ( .A0(n12000), .A1(B_sel_reg[0]), .B0(B_sel_reg[1]), .B1(
        n5829), .Y(n5422) );
  AOI22XL U21884 ( .A0(n12000), .A1(B_sel_reg[1]), .B0(B_sel_reg[2]), .B1(
        n5829), .Y(n5423) );
  AOI22XL U21885 ( .A0(n11997), .A1(B_sel_reg[2]), .B0(B_sel_reg[3]), .B1(
        n5829), .Y(n5424) );
  AOI22XL U21886 ( .A0(n11997), .A1(B_sel_reg[3]), .B0(D_sel_reg_4__0_), .B1(
        n5829), .Y(n5425) );
  AOI22XL U21887 ( .A0(n11997), .A1(D_sel_reg_4__0_), .B0(n11984), .B1(n5829), 
        .Y(n5426) );
  AOI22XL U21888 ( .A0(n11997), .A1(ram_sel_reg[1]), .B0(ram_sel_reg[3]), .B1(
        n5829), .Y(n5427) );
  AOI22XL U21889 ( .A0(n11997), .A1(ram_sel_reg[3]), .B0(ram_sel_reg[5]), .B1(
        n5829), .Y(n5428) );
  AOI22XL U21890 ( .A0(n11997), .A1(ram_sel_reg[5]), .B0(ram_sel_reg[7]), .B1(
        n5829), .Y(n5429) );
  AOI22XL U21891 ( .A0(n11997), .A1(ram_sel_reg[7]), .B0(ram_sel_reg[9]), .B1(
        n5829), .Y(n5430) );
  AOI22XL U21892 ( .A0(n11997), .A1(ram_sel_reg[9]), .B0(n11993), .B1(n5829), 
        .Y(n5431) );
  AOI22XL U21893 ( .A0(n11997), .A1(ram_sel_reg[0]), .B0(ram_sel_reg[2]), .B1(
        n5829), .Y(n5432) );
  AOI22XL U21894 ( .A0(n11997), .A1(ram_sel_reg[2]), .B0(ram_sel_reg[4]), .B1(
        n5829), .Y(n5433) );
  AOI22XL U21895 ( .A0(n11997), .A1(ram_sel_reg[4]), .B0(ram_sel_reg[6]), .B1(
        n5829), .Y(n5434) );
  AOI22XL U21896 ( .A0(n11997), .A1(ram_sel_reg[6]), .B0(ram_sel_reg[8]), .B1(
        n5829), .Y(n5435) );
  AOI22XL U21897 ( .A0(n11997), .A1(ram_sel_reg[8]), .B0(n11992), .B1(n5829), 
        .Y(n5436) );
  AOI22XL U21898 ( .A0(n11953), .A1(Q0_addr[11]), .B0(Q0_addr[3]), .B1(n5830), 
        .Y(n5437) );
  AOI22XL U21899 ( .A0(n11953), .A1(Q0_addr[19]), .B0(Q0_addr[11]), .B1(n5830), 
        .Y(n5438) );
  AOI22XL U21900 ( .A0(n11953), .A1(Q0_addr[27]), .B0(Q0_addr[19]), .B1(n11954), .Y(n5439) );
  AOI22XL U21901 ( .A0(n11953), .A1(Q0_addr[10]), .B0(Q0_addr[2]), .B1(n11958), 
        .Y(n5440) );
  AOI22XL U21902 ( .A0(n11953), .A1(Q0_addr[18]), .B0(Q0_addr[10]), .B1(n11957), .Y(n5441) );
  AOI22XL U21903 ( .A0(n5834), .A1(Q0_addr[26]), .B0(Q0_addr[18]), .B1(n11957), 
        .Y(n5442) );
  AOI22XL U21904 ( .A0(n5834), .A1(Q0_addr[9]), .B0(Q0_addr[1]), .B1(n11952), 
        .Y(n5443) );
  AOI22XL U21905 ( .A0(n5834), .A1(Q0_addr[17]), .B0(Q0_addr[9]), .B1(n11952), 
        .Y(n5444) );
  AOI22XL U21906 ( .A0(n5834), .A1(Q0_addr[25]), .B0(Q0_addr[17]), .B1(n11958), 
        .Y(n5445) );
  AOI22XL U21907 ( .A0(n5834), .A1(Q0_addr[8]), .B0(Q0_addr[0]), .B1(n11958), 
        .Y(n5446) );
  AOI22XL U21908 ( .A0(n5834), .A1(Q0_addr[16]), .B0(Q0_addr[8]), .B1(n11958), 
        .Y(n5447) );
  AOI22XL U21909 ( .A0(n5834), .A1(Q0_addr[24]), .B0(Q0_addr[16]), .B1(n5830), 
        .Y(n5448) );
  AOI22XL U21910 ( .A0(n5834), .A1(Q2_addr[13]), .B0(Q2_addr[5]), .B1(n11952), 
        .Y(n5449) );
  AOI22XL U21911 ( .A0(n5834), .A1(Q2_addr[21]), .B0(Q2_addr[13]), .B1(n11954), 
        .Y(n5450) );
  AOI22XL U21912 ( .A0(n5834), .A1(Q2_addr[29]), .B0(Q2_addr[21]), .B1(n11952), 
        .Y(n5451) );
  AOI22XL U21913 ( .A0(n5834), .A1(Q2_addr[37]), .B0(Q2_addr[29]), .B1(n11954), 
        .Y(n5452) );
  AOI22XL U21914 ( .A0(n5911), .A1(Q2_addr[11]), .B0(Q2_addr[3]), .B1(n5830), 
        .Y(n5454) );
  AOI22XL U21915 ( .A0(n5834), .A1(Q2_addr[19]), .B0(Q2_addr[11]), .B1(n11958), 
        .Y(n5455) );
  AOI22XL U21916 ( .A0(n5834), .A1(Q2_addr[27]), .B0(Q2_addr[19]), .B1(n11957), 
        .Y(n5456) );
  AOI22XL U21917 ( .A0(n5834), .A1(Q2_addr[35]), .B0(Q2_addr[27]), .B1(n11954), 
        .Y(n5457) );
  AOI22XL U21918 ( .A0(n5834), .A1(Q2_addr[10]), .B0(Q2_addr[2]), .B1(n11957), 
        .Y(n5459) );
  AOI22XL U21919 ( .A0(n5834), .A1(Q2_addr[18]), .B0(Q2_addr[10]), .B1(n11958), 
        .Y(n5460) );
  AOI22XL U21920 ( .A0(n5834), .A1(Q2_addr[26]), .B0(Q2_addr[18]), .B1(n11952), 
        .Y(n5461) );
  AOI22XL U21921 ( .A0(n5834), .A1(Q2_addr[34]), .B0(Q2_addr[26]), .B1(n11952), 
        .Y(n5462) );
  AOI22XL U21922 ( .A0(n5834), .A1(Q2_addr[9]), .B0(Q2_addr[1]), .B1(n11958), 
        .Y(n5464) );
  AOI22XL U21923 ( .A0(n5834), .A1(Q2_addr[17]), .B0(Q2_addr[9]), .B1(n11954), 
        .Y(n5465) );
  AOI22XL U21924 ( .A0(n5834), .A1(Q2_addr[25]), .B0(Q2_addr[17]), .B1(n11957), 
        .Y(n5466) );
  AOI22XL U21925 ( .A0(n5834), .A1(Q2_addr[33]), .B0(Q2_addr[25]), .B1(n5830), 
        .Y(n5467) );
  AOI22XL U21926 ( .A0(n11956), .A1(Q2_addr[8]), .B0(Q2_addr[0]), .B1(n11952), 
        .Y(n5469) );
  AOI22XL U21927 ( .A0(n5834), .A1(Q2_addr[16]), .B0(Q2_addr[8]), .B1(n11957), 
        .Y(n5470) );
  AOI22XL U21928 ( .A0(n5911), .A1(Q2_addr[24]), .B0(Q2_addr[16]), .B1(n11952), 
        .Y(n5471) );
  AOI22XL U21929 ( .A0(n5911), .A1(Q2_addr[32]), .B0(Q2_addr[24]), .B1(n11957), 
        .Y(n5472) );
  AOI22XL U21930 ( .A0(n5911), .A1(Q3_addr[13]), .B0(Q3_addr[5]), .B1(n11952), 
        .Y(n5474) );
  AOI22XL U21931 ( .A0(n5911), .A1(Q3_addr[21]), .B0(Q3_addr[13]), .B1(n11958), 
        .Y(n5475) );
  AOI22XL U21932 ( .A0(n5911), .A1(Q3_addr[29]), .B0(Q3_addr[21]), .B1(n11952), 
        .Y(n5476) );
  AOI22XL U21933 ( .A0(n5911), .A1(Q3_addr[37]), .B0(Q3_addr[29]), .B1(n5830), 
        .Y(n5477) );
  AOI22XL U21934 ( .A0(n5911), .A1(Q3_addr[12]), .B0(Q3_addr[4]), .B1(n11957), 
        .Y(n5478) );
  AOI22XL U21935 ( .A0(n5834), .A1(Q3_addr[20]), .B0(Q3_addr[12]), .B1(n5808), 
        .Y(n5479) );
  AOI22XL U21936 ( .A0(n5834), .A1(Q3_addr[36]), .B0(Q3_addr[28]), .B1(n5808), 
        .Y(n5481) );
  AOI22XL U21937 ( .A0(n11956), .A1(Q3_addr[11]), .B0(Q3_addr[3]), .B1(n5808), 
        .Y(n5482) );
  AOI22XL U21938 ( .A0(n5834), .A1(Q3_addr[19]), .B0(Q3_addr[11]), .B1(n5808), 
        .Y(n5483) );
  AOI22XL U21939 ( .A0(n5911), .A1(Q3_addr[27]), .B0(Q3_addr[19]), .B1(n5808), 
        .Y(n5484) );
  AOI22XL U21940 ( .A0(n5834), .A1(Q3_addr[35]), .B0(Q3_addr[27]), .B1(n5808), 
        .Y(n5485) );
  AOI22XL U21941 ( .A0(n11956), .A1(Q3_addr[10]), .B0(Q3_addr[2]), .B1(n5808), 
        .Y(n5486) );
  AOI22XL U21942 ( .A0(n11956), .A1(Q3_addr[18]), .B0(Q3_addr[10]), .B1(n5808), 
        .Y(n5487) );
  AOI22XL U21943 ( .A0(n11956), .A1(Q3_addr[26]), .B0(Q3_addr[18]), .B1(n5808), 
        .Y(n5488) );
  AOI22XL U21944 ( .A0(n5911), .A1(Q3_addr[34]), .B0(Q3_addr[26]), .B1(n5808), 
        .Y(n5489) );
  AOI22XL U21945 ( .A0(n5834), .A1(Q3_addr[9]), .B0(Q3_addr[1]), .B1(n5808), 
        .Y(n5490) );
  AOI22XL U21946 ( .A0(n11956), .A1(Q3_addr[17]), .B0(Q3_addr[9]), .B1(n5808), 
        .Y(n5491) );
  AOI22XL U21947 ( .A0(n5911), .A1(Q3_addr[25]), .B0(Q3_addr[17]), .B1(n5808), 
        .Y(n5492) );
  AOI22XL U21948 ( .A0(n11956), .A1(Q3_addr[33]), .B0(Q3_addr[25]), .B1(n5808), 
        .Y(n5493) );
  AOI22XL U21949 ( .A0(n11953), .A1(Q3_addr[8]), .B0(Q3_addr[0]), .B1(n11957), 
        .Y(n5494) );
  AOI22XL U21950 ( .A0(n11956), .A1(Q3_addr[16]), .B0(Q3_addr[8]), .B1(n5808), 
        .Y(n5495) );
  AOI22XL U21951 ( .A0(n5911), .A1(Q3_addr[24]), .B0(Q3_addr[16]), .B1(n5808), 
        .Y(n5496) );
  AOI22XL U21952 ( .A0(n11956), .A1(Q3_addr[32]), .B0(Q3_addr[24]), .B1(n5830), 
        .Y(n5497) );
  AOI22XL U21953 ( .A0(n11953), .A1(Q0_addr[35]), .B0(Q0_addr[27]), .B1(n11954), .Y(n5498) );
  AOI22XL U21954 ( .A0(n5911), .A1(Q0_addr[34]), .B0(Q0_addr[26]), .B1(n5830), 
        .Y(n5500) );
  AOI22XL U21955 ( .A0(n5834), .A1(Q0_addr[33]), .B0(Q0_addr[25]), .B1(n11954), 
        .Y(n5502) );
  AOI22XL U21956 ( .A0(n11956), .A1(Q0_addr[32]), .B0(Q0_addr[24]), .B1(n11954), .Y(n5504) );
  AOI22XL U21957 ( .A0(n5834), .A1(Q1_addr[12]), .B0(Q1_addr[4]), .B1(n11954), 
        .Y(n5506) );
  AOI22XL U21958 ( .A0(n5834), .A1(Q1_addr[20]), .B0(Q1_addr[12]), .B1(n5830), 
        .Y(n5507) );
  AOI22XL U21959 ( .A0(n5911), .A1(Q1_addr[28]), .B0(Q1_addr[20]), .B1(n11957), 
        .Y(n5508) );
  AOI22XL U21960 ( .A0(n11956), .A1(Q1_addr[36]), .B0(Q1_addr[28]), .B1(n5808), 
        .Y(n5509) );
  AOI22XL U21961 ( .A0(n11953), .A1(Q1_addr[11]), .B0(Q1_addr[3]), .B1(n11954), 
        .Y(n5511) );
  AOI22XL U21962 ( .A0(n5911), .A1(Q1_addr[19]), .B0(Q1_addr[11]), .B1(n5808), 
        .Y(n5512) );
  AOI22XL U21963 ( .A0(n5911), .A1(Q1_addr[27]), .B0(Q1_addr[19]), .B1(n5808), 
        .Y(n5513) );
  AOI22XL U21964 ( .A0(n5911), .A1(Q1_addr[35]), .B0(Q1_addr[27]), .B1(n11954), 
        .Y(n5514) );
  AOI22XL U21965 ( .A0(n11956), .A1(Q1_addr[18]), .B0(Q1_addr[10]), .B1(n5808), 
        .Y(n5517) );
  AOI22XL U21966 ( .A0(n5834), .A1(Q1_addr[26]), .B0(Q1_addr[18]), .B1(n5808), 
        .Y(n5518) );
  AOI22XL U21967 ( .A0(n11956), .A1(Q1_addr[9]), .B0(Q1_addr[1]), .B1(n5808), 
        .Y(n5521) );
  AOI22XL U21968 ( .A0(n11953), .A1(Q1_addr[17]), .B0(Q1_addr[9]), .B1(n5808), 
        .Y(n5522) );
  AOI22XL U21969 ( .A0(n11956), .A1(Q1_addr[25]), .B0(Q1_addr[17]), .B1(n5808), 
        .Y(n5523) );
  AOI22XL U21970 ( .A0(n5834), .A1(Q1_addr[8]), .B0(Q1_addr[0]), .B1(n11957), 
        .Y(n5526) );
  AOI22XL U21971 ( .A0(n11628), .A1(Q1_addr[16]), .B0(Q1_addr[8]), .B1(n5808), 
        .Y(n5527) );
  AOI22XL U21972 ( .A0(n5911), .A1(Q1_addr[24]), .B0(Q1_addr[16]), .B1(n5830), 
        .Y(n5528) );
  AOI22XL U21973 ( .A0(n5834), .A1(Q1_addr[32]), .B0(Q1_addr[24]), .B1(n11958), 
        .Y(n5529) );
  INVXL U21974 ( .A(T1_rom2_q[0]), .Y(n29176) );
  INVXL U21975 ( .A(T1_rom2_q[10]), .Y(n29175) );
  INVXL U21976 ( .A(T1_rom2_q[11]), .Y(n29174) );
  INVXL U21977 ( .A(T1_rom2_q[12]), .Y(n29173) );
  INVXL U21978 ( .A(T1_rom2_q[13]), .Y(n29172) );
  INVXL U21979 ( .A(T1_rom2_q[14]), .Y(n29171) );
  INVXL U21980 ( .A(T1_rom2_q[16]), .Y(n29169) );
  INVXL U21981 ( .A(T1_rom2_q[17]), .Y(n29168) );
  INVXL U21982 ( .A(T1_rom2_q[18]), .Y(n29167) );
  INVXL U21983 ( .A(T1_rom2_q[19]), .Y(n29166) );
  INVXL U21984 ( .A(T1_rom2_q[1]), .Y(n29165) );
  INVXL U21985 ( .A(T1_rom2_q[20]), .Y(n29164) );
  INVXL U21986 ( .A(T1_rom2_q[21]), .Y(n29163) );
  INVXL U21987 ( .A(T1_rom2_q[22]), .Y(n29162) );
  INVXL U21988 ( .A(T1_rom2_q[24]), .Y(n29160) );
  INVXL U21989 ( .A(T1_rom2_q[25]), .Y(n29159) );
  INVXL U21990 ( .A(T1_rom2_q[28]), .Y(n29156) );
  INVXL U21991 ( .A(T1_rom2_q[29]), .Y(n29155) );
  INVXL U21992 ( .A(T1_rom2_q[2]), .Y(n29154) );
  INVXL U21993 ( .A(T1_rom2_q[30]), .Y(n29153) );
  INVXL U21994 ( .A(T1_rom2_q[31]), .Y(n29152) );
  INVXL U21995 ( .A(T1_rom2_q[3]), .Y(n29151) );
  INVXL U21996 ( .A(T1_rom2_q[4]), .Y(n29150) );
  INVXL U21997 ( .A(T1_rom2_q[5]), .Y(n29149) );
  INVXL U21998 ( .A(T1_rom2_q[6]), .Y(n29148) );
  INVXL U21999 ( .A(T1_rom2_q[7]), .Y(n29147) );
  INVXL U22000 ( .A(T1_rom2_q[8]), .Y(n29146) );
  INVXL U22001 ( .A(T1_rom2_q[9]), .Y(n29145) );
  INVXL U22002 ( .A(T1_rom1_q[0]), .Y(n29208) );
  INVXL U22003 ( .A(T1_rom1_q[10]), .Y(n29207) );
  INVXL U22004 ( .A(T1_rom1_q[12]), .Y(n29205) );
  INVXL U22005 ( .A(T1_rom1_q[13]), .Y(n29204) );
  INVXL U22006 ( .A(T1_rom1_q[14]), .Y(n29203) );
  INVXL U22007 ( .A(T1_rom1_q[15]), .Y(n29202) );
  INVXL U22008 ( .A(T1_rom1_q[16]), .Y(n29201) );
  INVXL U22009 ( .A(T1_rom1_q[17]), .Y(n29200) );
  INVXL U22010 ( .A(T1_rom1_q[1]), .Y(n29197) );
  INVXL U22011 ( .A(T1_rom1_q[20]), .Y(n29196) );
  INVXL U22012 ( .A(T1_rom1_q[21]), .Y(n29195) );
  INVXL U22013 ( .A(T1_rom1_q[22]), .Y(n29194) );
  INVXL U22014 ( .A(T1_rom1_q[24]), .Y(n29192) );
  INVXL U22015 ( .A(T1_rom1_q[26]), .Y(n29190) );
  INVXL U22016 ( .A(T1_rom1_q[28]), .Y(n29188) );
  INVXL U22017 ( .A(T1_rom1_q[29]), .Y(n29187) );
  INVXL U22018 ( .A(T1_rom1_q[2]), .Y(n29186) );
  INVXL U22019 ( .A(T1_rom1_q[30]), .Y(n29185) );
  INVXL U22020 ( .A(T1_rom1_q[31]), .Y(n29184) );
  INVXL U22021 ( .A(T1_rom1_q[3]), .Y(n29183) );
  INVXL U22022 ( .A(T1_rom1_q[4]), .Y(n29182) );
  INVXL U22023 ( .A(T1_rom1_q[5]), .Y(n29181) );
  INVXL U22024 ( .A(T1_rom1_q[6]), .Y(n29180) );
  INVXL U22025 ( .A(T1_rom1_q[7]), .Y(n29179) );
  INVXL U22026 ( .A(T1_rom1_q[8]), .Y(n29178) );
  INVXL U22027 ( .A(T1_rom0_q[0]), .Y(n29240) );
  INVXL U22028 ( .A(T1_rom0_q[10]), .Y(n29239) );
  INVXL U22029 ( .A(T1_rom0_q[11]), .Y(n29238) );
  INVXL U22030 ( .A(T1_rom0_q[12]), .Y(n29237) );
  INVXL U22031 ( .A(T1_rom0_q[13]), .Y(n29236) );
  INVXL U22032 ( .A(T1_rom0_q[14]), .Y(n29235) );
  INVXL U22033 ( .A(T1_rom0_q[15]), .Y(n29234) );
  INVXL U22034 ( .A(T1_rom0_q[16]), .Y(n29233) );
  INVXL U22035 ( .A(T1_rom0_q[17]), .Y(n29232) );
  INVXL U22036 ( .A(T1_rom0_q[18]), .Y(n29231) );
  INVXL U22037 ( .A(T1_rom0_q[1]), .Y(n29229) );
  INVXL U22038 ( .A(T1_rom0_q[20]), .Y(n29228) );
  INVXL U22039 ( .A(T1_rom0_q[21]), .Y(n29227) );
  INVXL U22040 ( .A(T1_rom0_q[22]), .Y(n29226) );
  INVXL U22041 ( .A(T1_rom0_q[24]), .Y(n29224) );
  INVXL U22042 ( .A(T1_rom0_q[26]), .Y(n29222) );
  INVXL U22043 ( .A(T1_rom0_q[27]), .Y(n29221) );
  INVXL U22044 ( .A(T1_rom0_q[28]), .Y(n29220) );
  INVXL U22045 ( .A(T1_rom0_q[29]), .Y(n29219) );
  INVXL U22046 ( .A(T1_rom0_q[2]), .Y(n29218) );
  INVXL U22047 ( .A(T1_rom0_q[30]), .Y(n29217) );
  INVXL U22048 ( .A(T1_rom0_q[31]), .Y(n29216) );
  INVXL U22049 ( .A(T1_rom0_q[3]), .Y(n29215) );
  INVXL U22050 ( .A(T1_rom0_q[4]), .Y(n29214) );
  INVXL U22051 ( .A(T1_rom0_q[5]), .Y(n29213) );
  INVXL U22052 ( .A(T1_rom0_q[6]), .Y(n29212) );
  INVXL U22053 ( .A(T1_rom0_q[7]), .Y(n29211) );
  INVXL U22054 ( .A(T1_rom0_q[8]), .Y(n29210) );
  INVXL U22055 ( .A(T1_rom0_q[9]), .Y(n29209) );
  AOI22XL U22056 ( .A0(cnt[9]), .A1(n28634), .B0(n11996), .B1(n28758), .Y(
        n5638) );
  INVXL U22057 ( .A(T1_rom3_q[0]), .Y(n29144) );
  INVXL U22058 ( .A(T1_rom3_q[10]), .Y(n29143) );
  INVXL U22059 ( .A(T1_rom3_q[12]), .Y(n29141) );
  INVXL U22060 ( .A(T1_rom3_q[14]), .Y(n29139) );
  INVXL U22061 ( .A(T1_rom3_q[16]), .Y(n29137) );
  INVXL U22062 ( .A(T1_rom3_q[17]), .Y(n29136) );
  INVXL U22063 ( .A(T1_rom3_q[18]), .Y(n29135) );
  INVXL U22064 ( .A(T1_rom3_q[19]), .Y(n29134) );
  INVXL U22065 ( .A(T1_rom3_q[1]), .Y(n29133) );
  INVXL U22066 ( .A(T1_rom3_q[20]), .Y(n29132) );
  INVXL U22067 ( .A(T1_rom3_q[21]), .Y(n29131) );
  INVXL U22068 ( .A(T1_rom3_q[22]), .Y(n29130) );
  INVXL U22069 ( .A(T1_rom3_q[23]), .Y(n29129) );
  INVXL U22070 ( .A(T1_rom3_q[24]), .Y(n29128) );
  INVXL U22071 ( .A(T1_rom3_q[26]), .Y(n29126) );
  INVXL U22072 ( .A(T1_rom3_q[27]), .Y(n29125) );
  INVXL U22073 ( .A(T1_rom3_q[28]), .Y(n29124) );
  INVXL U22074 ( .A(T1_rom3_q[29]), .Y(n29123) );
  INVXL U22075 ( .A(T1_rom3_q[2]), .Y(n29122) );
  INVXL U22076 ( .A(T1_rom3_q[30]), .Y(n29121) );
  INVXL U22077 ( .A(T1_rom3_q[31]), .Y(n29120) );
  INVXL U22078 ( .A(T1_rom3_q[3]), .Y(n29119) );
  INVXL U22079 ( .A(T1_rom3_q[4]), .Y(n29118) );
  INVXL U22080 ( .A(T1_rom3_q[5]), .Y(n29117) );
  INVXL U22081 ( .A(T1_rom3_q[6]), .Y(n29116) );
  INVXL U22082 ( .A(T1_rom3_q[9]), .Y(n29113) );
  NAND2XL U22083 ( .A(n28633), .B(n11955), .Y(n5678) );
  AOI22XL U22084 ( .A0(n11980), .A1(cnt[11]), .B0(n11979), .B1(n11978), .Y(
        n5680) );
  NOR2XL U22085 ( .A(cnt[11]), .B(n28635), .Y(n11978) );
  INVXL U22086 ( .A(n11948), .Y(n11629) );
  INVXL U22087 ( .A(n11946), .Y(n11947) );
  NAND2XL U22088 ( .A(n11951), .B(n11873), .Y(n5694) );
  NAND2XL U22089 ( .A(n11980), .B(n11977), .Y(n5688) );
  NAND2XL U22090 ( .A(n11644), .B(n11643), .Y(T1_rom_addr[7]) );
  AOI22XL U22091 ( .A0(cnt[7]), .A1(n11648), .B0(cnt[3]), .B1(n11979), .Y(
        n11644) );
  AOI22XL U22092 ( .A0(cnt[5]), .A1(n11647), .B0(cnt[1]), .B1(n11652), .Y(
        n11643) );
  AOI22XL U22093 ( .A0(cnt[6]), .A1(n11648), .B0(cnt[2]), .B1(n11979), .Y(
        n11649) );
  AOI22XL U22094 ( .A0(cnt[4]), .A1(n11647), .B0(cnt[0]), .B1(n11652), .Y(
        n11650) );
  NOR2XL U22095 ( .A(n28704), .B(n14977), .Y(n7134) );
  NOR2XL U22096 ( .A(n28680), .B(n14979), .Y(n7133) );
  NOR2XL U22097 ( .A(n11991), .B(n11987), .Y(A7_WEN) );
  AOI211XL U22098 ( .A0(n5826), .A1(n27555), .B0(n28349), .C0(n27116), .Y(
        n27117) );
  OAI22XL U22099 ( .A0(n27959), .A1(n27553), .B0(n7140), .B1(n27552), .Y(
        n27116) );
  AOI211XL U22100 ( .A0(n5826), .A1(n27549), .B0(n28342), .C0(n27113), .Y(
        n27114) );
  OAI22XL U22101 ( .A0(n27959), .A1(n27547), .B0(n7140), .B1(n27546), .Y(
        n27113) );
  AOI211XL U22102 ( .A0(n27162), .A1(n27543), .B0(n28335), .C0(n27110), .Y(
        n27111) );
  OAI22XL U22103 ( .A0(n27959), .A1(n27541), .B0(n27540), .B1(n5823), .Y(
        n27110) );
  AOI211XL U22104 ( .A0(n27162), .A1(n27537), .B0(n28328), .C0(n27107), .Y(
        n27108) );
  OAI22XL U22105 ( .A0(n27959), .A1(n27535), .B0(n7140), .B1(n27534), .Y(
        n27107) );
  OAI22XL U22106 ( .A0(n27959), .A1(n27529), .B0(n7140), .B1(n27528), .Y(
        n27104) );
  AOI211XL U22107 ( .A0(n27162), .A1(n27811), .B0(n28625), .C0(n27279), .Y(
        n27280) );
  OAI22XL U22108 ( .A0(n27959), .A1(n27809), .B0(n27813), .B1(n28054), .Y(
        n27279) );
  AOI211XL U22109 ( .A0(n27162), .A1(n27805), .B0(n28625), .C0(n27275), .Y(
        n27276) );
  OAI22XL U22110 ( .A0(n27959), .A1(n27803), .B0(n27807), .B1(n5823), .Y(
        n27275) );
  OAI22XL U22111 ( .A0(n27959), .A1(n27523), .B0(n27522), .B1(n5823), .Y(
        n27101) );
  AOI211XL U22112 ( .A0(n27162), .A1(n27799), .B0(n28625), .C0(n27271), .Y(
        n27272) );
  OAI22XL U22113 ( .A0(n27959), .A1(n27797), .B0(n27801), .B1(n5823), .Y(
        n27271) );
  OAI22XL U22114 ( .A0(n27959), .A1(n27791), .B0(n28050), .B1(n27795), .Y(
        n27267) );
  OAI22XL U22115 ( .A0(n27959), .A1(n27785), .B0(n7140), .B1(n27784), .Y(
        n27262) );
  AOI211XL U22116 ( .A0(n27162), .A1(n27781), .B0(n28625), .C0(n27258), .Y(
        n27259) );
  OAI22XL U22117 ( .A0(n27959), .A1(n27779), .B0(n7140), .B1(n27783), .Y(
        n27258) );
  OAI22XL U22118 ( .A0(n27959), .A1(n27773), .B0(n27777), .B1(n5823), .Y(
        n27254) );
  AOI211XL U22119 ( .A0(n27162), .A1(n27768), .B0(n28625), .C0(n27250), .Y(
        n27251) );
  OAI22XL U22120 ( .A0(n27959), .A1(n27766), .B0(n27765), .B1(n5823), .Y(
        n27250) );
  AOI211XL U22121 ( .A0(n27162), .A1(n27762), .B0(n28625), .C0(n27246), .Y(
        n27247) );
  OAI22XL U22122 ( .A0(n27959), .A1(n27760), .B0(n27759), .B1(n5823), .Y(
        n27246) );
  AOI211XL U22123 ( .A0(n5826), .A1(n27756), .B0(n28625), .C0(n27242), .Y(
        n27243) );
  OAI22XL U22124 ( .A0(n27959), .A1(n27754), .B0(n7140), .B1(n27758), .Y(
        n27242) );
  AOI211XL U22125 ( .A0(n27162), .A1(n27750), .B0(n28625), .C0(n27238), .Y(
        n27239) );
  OAI22XL U22126 ( .A0(n27959), .A1(n27748), .B0(n27747), .B1(n28054), .Y(
        n27238) );
  AOI211XL U22127 ( .A0(n27162), .A1(n27744), .B0(n28557), .C0(n27233), .Y(
        n27234) );
  OAI22XL U22128 ( .A0(n27959), .A1(n27742), .B0(n7140), .B1(n27746), .Y(
        n27233) );
  AOI211XL U22129 ( .A0(n27162), .A1(n27519), .B0(n28306), .C0(n27098), .Y(
        n27099) );
  OAI22XL U22130 ( .A0(n27959), .A1(n27517), .B0(n7140), .B1(n27521), .Y(
        n27098) );
  AOI211XL U22131 ( .A0(n5826), .A1(n27738), .B0(n28550), .C0(n27229), .Y(
        n27230) );
  OAI22XL U22132 ( .A0(n27959), .A1(n27736), .B0(n7140), .B1(n27735), .Y(
        n27229) );
  AOI211XL U22133 ( .A0(n27162), .A1(n27732), .B0(n28543), .C0(n27225), .Y(
        n27226) );
  OAI22XL U22134 ( .A0(n27959), .A1(n27730), .B0(n7140), .B1(n7104), .Y(n27225) );
  AOI211XL U22135 ( .A0(n27162), .A1(n27726), .B0(n28536), .C0(n27221), .Y(
        n27222) );
  OAI22XL U22136 ( .A0(n27959), .A1(n27724), .B0(n7140), .B1(n27728), .Y(
        n27221) );
  AOI211XL U22137 ( .A0(n27162), .A1(n27720), .B0(n28529), .C0(n27217), .Y(
        n27218) );
  OAI22XL U22138 ( .A0(n27959), .A1(n27718), .B0(n7140), .B1(n27717), .Y(
        n27217) );
  OAI22XL U22139 ( .A0(n27959), .A1(n27712), .B0(n28050), .B1(n27716), .Y(
        n27214) );
  AOI211XL U22140 ( .A0(n27162), .A1(n27708), .B0(n28515), .C0(n27209), .Y(
        n27210) );
  OAI22XL U22141 ( .A0(n27959), .A1(n27706), .B0(n7140), .B1(n27710), .Y(
        n27209) );
  OAI22XL U22142 ( .A0(n27959), .A1(n27700), .B0(n27704), .B1(n5823), .Y(
        n27206) );
  OAI22XL U22143 ( .A0(n27959), .A1(n27694), .B0(n27693), .B1(n5823), .Y(
        n27202) );
  AOI211XL U22144 ( .A0(n5826), .A1(n27690), .B0(n28494), .C0(n27199), .Y(
        n27200) );
  OAI22XL U22145 ( .A0(n27959), .A1(n27688), .B0(n7140), .B1(n27692), .Y(
        n27199) );
  AOI211XL U22146 ( .A0(n27162), .A1(n27683), .B0(n28487), .C0(n27196), .Y(
        n27197) );
  OAI22XL U22147 ( .A0(n27959), .A1(n27681), .B0(n7140), .B1(n27680), .Y(
        n27196) );
  OAI22XL U22148 ( .A0(n27959), .A1(n27511), .B0(n7140), .B1(n27515), .Y(
        n27095) );
  AOI211XL U22149 ( .A0(n27162), .A1(n27677), .B0(n28480), .C0(n27193), .Y(
        n27194) );
  OAI22XL U22150 ( .A0(n27959), .A1(n27675), .B0(n27679), .B1(n5823), .Y(
        n27193) );
  AOI211XL U22151 ( .A0(n5826), .A1(n27671), .B0(n28473), .C0(n27190), .Y(
        n27191) );
  OAI22XL U22152 ( .A0(n27959), .A1(n27669), .B0(n7140), .B1(n27673), .Y(
        n27190) );
  OAI22XL U22153 ( .A0(n27959), .A1(n27663), .B0(n7140), .B1(n27667), .Y(
        n27187) );
  OAI22XL U22154 ( .A0(n27959), .A1(n27657), .B0(n7140), .B1(n27656), .Y(
        n27184) );
  OAI22XL U22155 ( .A0(n27959), .A1(n27651), .B0(n27650), .B1(n5823), .Y(
        n27181) );
  OAI22XL U22156 ( .A0(n27959), .A1(n27645), .B0(n7140), .B1(n27644), .Y(
        n27177) );
  AOI211XL U22157 ( .A0(n27162), .A1(n27641), .B0(n28452), .C0(n27173), .Y(
        n27174) );
  OAI22XL U22158 ( .A0(n27959), .A1(n27639), .B0(n7140), .B1(n27643), .Y(
        n27173) );
  OAI22XL U22159 ( .A0(n27959), .A1(n27633), .B0(n7140), .B1(n27632), .Y(
        n27169) );
  AOI211XL U22160 ( .A0(n27162), .A1(n27628), .B0(n28452), .C0(n27165), .Y(
        n27166) );
  OAI22XL U22161 ( .A0(n27959), .A1(n27626), .B0(n7140), .B1(n27625), .Y(
        n27165) );
  AOI211XL U22162 ( .A0(n27162), .A1(n27622), .B0(n28452), .C0(n27160), .Y(
        n27161) );
  OAI22XL U22163 ( .A0(n27959), .A1(n27620), .B0(n27619), .B1(n5823), .Y(
        n27160) );
  OAI22XL U22164 ( .A0(n27959), .A1(n27505), .B0(n7140), .B1(n27509), .Y(
        n27092) );
  AOI211XL U22165 ( .A0(n27162), .A1(n27616), .B0(n28452), .C0(n27156), .Y(
        n27157) );
  OAI22XL U22166 ( .A0(n27959), .A1(n27614), .B0(n7140), .B1(n27613), .Y(
        n27156) );
  AOI211XL U22167 ( .A0(n27162), .A1(n27610), .B0(n28452), .C0(n27152), .Y(
        n27153) );
  OAI22XL U22168 ( .A0(n27959), .A1(n27608), .B0(n7140), .B1(n7102), .Y(n27152) );
  AOI211XL U22169 ( .A0(n27162), .A1(n27604), .B0(n28452), .C0(n27148), .Y(
        n27149) );
  OAI22XL U22170 ( .A0(n27959), .A1(n27602), .B0(n7114), .B1(n5823), .Y(n27148) );
  AOI211XL U22171 ( .A0(n27162), .A1(n27598), .B0(n28452), .C0(n27144), .Y(
        n27145) );
  OAI22XL U22172 ( .A0(n27959), .A1(n27596), .B0(n7140), .B1(n27600), .Y(
        n27144) );
  AOI211XL U22173 ( .A0(n27162), .A1(n27592), .B0(n28452), .C0(n27140), .Y(
        n27141) );
  OAI22XL U22174 ( .A0(n27959), .A1(n27590), .B0(n27589), .B1(n5823), .Y(
        n27140) );
  OAI22XL U22175 ( .A0(n27959), .A1(n27584), .B0(n7112), .B1(n5823), .Y(n27136) );
  OAI22XL U22176 ( .A0(n27959), .A1(n27578), .B0(n7140), .B1(n27582), .Y(
        n27132) );
  OAI22XL U22177 ( .A0(n27959), .A1(n27572), .B0(n27571), .B1(n5823), .Y(
        n27128) );
  AOI211XL U22178 ( .A0(n27162), .A1(n27568), .B0(n28364), .C0(n27124), .Y(
        n27125) );
  OAI22XL U22179 ( .A0(n27959), .A1(n27566), .B0(n27565), .B1(n5823), .Y(
        n27124) );
  AOI211XL U22180 ( .A0(n27162), .A1(n27562), .B0(n28357), .C0(n27119), .Y(
        n27120) );
  OAI22XL U22181 ( .A0(n27959), .A1(n27559), .B0(n27564), .B1(n5823), .Y(
        n27119) );
  AOI211XL U22182 ( .A0(n27162), .A1(n27501), .B0(n7120), .C0(n27089), .Y(
        n27090) );
  OAI22XL U22183 ( .A0(n27959), .A1(n27499), .B0(n7140), .B1(n27498), .Y(
        n27089) );
  NOR2XL U22184 ( .A(n11991), .B(n11981), .Y(A6_WEN) );
  AOI211XL U22185 ( .A0(n5921), .A1(n27555), .B0(n28349), .C0(n27301), .Y(
        n27302) );
  OAI22XL U22186 ( .A0(n28125), .A1(n27553), .B0(n27379), .B1(n27552), .Y(
        n27301) );
  AOI211XL U22187 ( .A0(n5921), .A1(n27549), .B0(n28342), .C0(n27299), .Y(
        n27300) );
  OAI22XL U22188 ( .A0(n28125), .A1(n27547), .B0(n27551), .B1(n28138), .Y(
        n27299) );
  AOI211XL U22189 ( .A0(n28143), .A1(n27543), .B0(n28335), .C0(n27296), .Y(
        n27297) );
  OAI22XL U22190 ( .A0(n28125), .A1(n27541), .B0(n27379), .B1(n27545), .Y(
        n27296) );
  AOI211XL U22191 ( .A0(n28143), .A1(n27537), .B0(n28328), .C0(n27294), .Y(
        n27295) );
  OAI22XL U22192 ( .A0(n28125), .A1(n27535), .B0(n27379), .B1(n27534), .Y(
        n27294) );
  OAI22XL U22193 ( .A0(n28125), .A1(n27529), .B0(n27533), .B1(n28093), .Y(
        n27292) );
  AOI211XL U22194 ( .A0(n28143), .A1(n27811), .B0(n28625), .C0(n27387), .Y(
        n27388) );
  OAI22XL U22195 ( .A0(n28125), .A1(n27809), .B0(n27813), .B1(n27386), .Y(
        n27387) );
  AOI211XL U22196 ( .A0(n28143), .A1(n27805), .B0(n28625), .C0(n27384), .Y(
        n27385) );
  OAI22XL U22197 ( .A0(n28125), .A1(n27803), .B0(n27807), .B1(n27386), .Y(
        n27384) );
  OAI22XL U22198 ( .A0(n28125), .A1(n27523), .B0(n27379), .B1(n27527), .Y(
        n27290) );
  AOI211XL U22199 ( .A0(n28143), .A1(n27799), .B0(n28625), .C0(n27382), .Y(
        n27383) );
  OAI22XL U22200 ( .A0(n28125), .A1(n27797), .B0(n28068), .B1(n27796), .Y(
        n27382) );
  OAI22XL U22201 ( .A0(n28125), .A1(n27791), .B0(n27379), .B1(n27795), .Y(
        n27380) );
  AOI211XL U22202 ( .A0(n28143), .A1(n27787), .B0(n28625), .C0(n27377), .Y(
        n27378) );
  OAI22XL U22203 ( .A0(n28125), .A1(n27785), .B0(n27789), .B1(n28118), .Y(
        n27377) );
  AOI211XL U22204 ( .A0(n28143), .A1(n27781), .B0(n28625), .C0(n27375), .Y(
        n27376) );
  OAI22XL U22205 ( .A0(n28125), .A1(n27779), .B0(n27778), .B1(n28093), .Y(
        n27375) );
  AOI211XL U22206 ( .A0(n28143), .A1(n27775), .B0(n28625), .C0(n27373), .Y(
        n27374) );
  OAI22XL U22207 ( .A0(n28125), .A1(n27773), .B0(n27777), .B1(n28138), .Y(
        n27373) );
  AOI211XL U22208 ( .A0(n28143), .A1(n27768), .B0(n28625), .C0(n27371), .Y(
        n27372) );
  OAI22XL U22209 ( .A0(n28125), .A1(n27766), .B0(n27765), .B1(n28093), .Y(
        n27371) );
  AOI211XL U22210 ( .A0(n28143), .A1(n27762), .B0(n28625), .C0(n27369), .Y(
        n27370) );
  OAI22XL U22211 ( .A0(n28125), .A1(n27760), .B0(n27759), .B1(n28093), .Y(
        n27369) );
  AOI211XL U22212 ( .A0(n28143), .A1(n27756), .B0(n28625), .C0(n27367), .Y(
        n27368) );
  OAI22XL U22213 ( .A0(n28125), .A1(n27754), .B0(n27753), .B1(n28158), .Y(
        n27367) );
  AOI211XL U22214 ( .A0(n28143), .A1(n27750), .B0(n28625), .C0(n27365), .Y(
        n27366) );
  OAI22XL U22215 ( .A0(n28125), .A1(n27748), .B0(n27747), .B1(n28165), .Y(
        n27365) );
  AOI211XL U22216 ( .A0(n5921), .A1(n27744), .B0(n28557), .C0(n27363), .Y(
        n27364) );
  OAI22XL U22217 ( .A0(n28125), .A1(n27742), .B0(n27379), .B1(n27746), .Y(
        n27363) );
  AOI211XL U22218 ( .A0(n28143), .A1(n27519), .B0(n28306), .C0(n27288), .Y(
        n27289) );
  OAI22XL U22219 ( .A0(n28125), .A1(n27517), .B0(n27516), .B1(n28093), .Y(
        n27288) );
  AOI211XL U22220 ( .A0(n28143), .A1(n27738), .B0(n28550), .C0(n27361), .Y(
        n27362) );
  OAI22XL U22221 ( .A0(n28125), .A1(n27736), .B0(n28068), .B1(n27735), .Y(
        n27361) );
  AOI211XL U22222 ( .A0(n5921), .A1(n27732), .B0(n28543), .C0(n27359), .Y(
        n27360) );
  OAI22XL U22223 ( .A0(n28125), .A1(n27730), .B0(n27729), .B1(n27386), .Y(
        n27359) );
  AOI211XL U22224 ( .A0(n28143), .A1(n27726), .B0(n28536), .C0(n27357), .Y(
        n27358) );
  OAI22XL U22225 ( .A0(n28125), .A1(n27724), .B0(n27723), .B1(n28138), .Y(
        n27357) );
  AOI211XL U22226 ( .A0(n5921), .A1(n27720), .B0(n28529), .C0(n27355), .Y(
        n27356) );
  OAI22XL U22227 ( .A0(n28125), .A1(n27718), .B0(n28068), .B1(n27717), .Y(
        n27355) );
  OAI22XL U22228 ( .A0(n28125), .A1(n27712), .B0(n28068), .B1(n27716), .Y(
        n27353) );
  AOI211XL U22229 ( .A0(n5921), .A1(n27708), .B0(n28515), .C0(n27351), .Y(
        n27352) );
  OAI22XL U22230 ( .A0(n28125), .A1(n27706), .B0(n27705), .B1(n28138), .Y(
        n27351) );
  OAI22XL U22231 ( .A0(n28125), .A1(n27700), .B0(n27704), .B1(n28138), .Y(
        n27349) );
  OAI22XL U22232 ( .A0(n28125), .A1(n27694), .B0(n27693), .B1(n28138), .Y(
        n27347) );
  AOI211XL U22233 ( .A0(n28143), .A1(n27690), .B0(n28494), .C0(n27345), .Y(
        n27346) );
  OAI22XL U22234 ( .A0(n28125), .A1(n27688), .B0(n27687), .B1(n28138), .Y(
        n27345) );
  AOI211XL U22235 ( .A0(n28143), .A1(n27683), .B0(n28487), .C0(n27343), .Y(
        n27344) );
  OAI22XL U22236 ( .A0(n28125), .A1(n27681), .B0(n27379), .B1(n27680), .Y(
        n27343) );
  OAI22XL U22237 ( .A0(n28125), .A1(n27511), .B0(n27379), .B1(n27515), .Y(
        n27286) );
  AOI211XL U22238 ( .A0(n28143), .A1(n27677), .B0(n28480), .C0(n27341), .Y(
        n27342) );
  OAI22XL U22239 ( .A0(n28125), .A1(n27675), .B0(n27679), .B1(n28138), .Y(
        n27341) );
  AOI211XL U22240 ( .A0(n28143), .A1(n27671), .B0(n28473), .C0(n27339), .Y(
        n27340) );
  OAI22XL U22241 ( .A0(n28125), .A1(n27669), .B0(n27379), .B1(n27673), .Y(
        n27339) );
  OAI22XL U22242 ( .A0(n28125), .A1(n27663), .B0(n27662), .B1(n28138), .Y(
        n27337) );
  OAI22XL U22243 ( .A0(n28125), .A1(n27657), .B0(n27661), .B1(n28093), .Y(
        n27335) );
  AOI211XL U22244 ( .A0(n28143), .A1(n27653), .B0(n28452), .C0(n27333), .Y(
        n27334) );
  OAI22XL U22245 ( .A0(n28125), .A1(n27651), .B0(n27650), .B1(n28093), .Y(
        n27333) );
  AOI211XL U22246 ( .A0(n28143), .A1(n27647), .B0(n28452), .C0(n27331), .Y(
        n27332) );
  OAI22XL U22247 ( .A0(n28125), .A1(n27645), .B0(n27379), .B1(n27644), .Y(
        n27331) );
  AOI211XL U22248 ( .A0(n28143), .A1(n27641), .B0(n28452), .C0(n27329), .Y(
        n27330) );
  OAI22XL U22249 ( .A0(n28125), .A1(n27639), .B0(n28068), .B1(n27643), .Y(
        n27329) );
  AOI211XL U22250 ( .A0(n28143), .A1(n27635), .B0(n28452), .C0(n27327), .Y(
        n27328) );
  OAI22XL U22251 ( .A0(n28125), .A1(n27633), .B0(n27637), .B1(n28138), .Y(
        n27327) );
  AOI211XL U22252 ( .A0(n28143), .A1(n27628), .B0(n28452), .C0(n27325), .Y(
        n27326) );
  OAI22XL U22253 ( .A0(n28125), .A1(n27626), .B0(n27630), .B1(n28093), .Y(
        n27325) );
  AOI211XL U22254 ( .A0(n28143), .A1(n27622), .B0(n28452), .C0(n27323), .Y(
        n27324) );
  OAI22XL U22255 ( .A0(n28125), .A1(n27620), .B0(n27619), .B1(n28138), .Y(
        n27323) );
  OAI22XL U22256 ( .A0(n28125), .A1(n27505), .B0(n27379), .B1(n27509), .Y(
        n27284) );
  AOI211XL U22257 ( .A0(n5921), .A1(n27616), .B0(n28452), .C0(n27321), .Y(
        n27322) );
  OAI22XL U22258 ( .A0(n28125), .A1(n27614), .B0(n27379), .B1(n27613), .Y(
        n27321) );
  AOI211XL U22259 ( .A0(n5921), .A1(n27610), .B0(n28452), .C0(n27319), .Y(
        n27320) );
  OAI22XL U22260 ( .A0(n28125), .A1(n27608), .B0(n27607), .B1(n28093), .Y(
        n27319) );
  AOI211XL U22261 ( .A0(n5921), .A1(n27604), .B0(n28452), .C0(n27317), .Y(
        n27318) );
  OAI22XL U22262 ( .A0(n28125), .A1(n27602), .B0(n27379), .B1(n27601), .Y(
        n27317) );
  AOI211XL U22263 ( .A0(n5921), .A1(n27598), .B0(n28452), .C0(n27315), .Y(
        n27316) );
  OAI22XL U22264 ( .A0(n28125), .A1(n27596), .B0(n27379), .B1(n27600), .Y(
        n27315) );
  AOI211XL U22265 ( .A0(n5921), .A1(n27592), .B0(n28452), .C0(n27313), .Y(
        n27314) );
  OAI22XL U22266 ( .A0(n28125), .A1(n27590), .B0(n27379), .B1(n7100), .Y(
        n27313) );
  OAI22XL U22267 ( .A0(n28125), .A1(n27584), .B0(n27379), .B1(n27583), .Y(
        n27311) );
  OAI22XL U22268 ( .A0(n28125), .A1(n27578), .B0(n27577), .B1(n28138), .Y(
        n27309) );
  OAI22XL U22269 ( .A0(n28125), .A1(n27572), .B0(n27571), .B1(n28093), .Y(
        n27307) );
  AOI211XL U22270 ( .A0(n5921), .A1(n27568), .B0(n28364), .C0(n27305), .Y(
        n27306) );
  OAI22XL U22271 ( .A0(n28125), .A1(n27566), .B0(n27379), .B1(n7098), .Y(
        n27305) );
  AOI211XL U22272 ( .A0(n5921), .A1(n27562), .B0(n28357), .C0(n27303), .Y(
        n27304) );
  OAI22XL U22273 ( .A0(n28125), .A1(n27559), .B0(n27564), .B1(n28093), .Y(
        n27303) );
  AOI211XL U22274 ( .A0(n28143), .A1(n27501), .B0(n7120), .C0(n27282), .Y(
        n27283) );
  OAI22XL U22275 ( .A0(n28125), .A1(n27499), .B0(n27379), .B1(n27498), .Y(
        n27282) );
  NOR2XL U22276 ( .A(n11991), .B(n11990), .Y(A5_WEN) );
  AOI211XL U22277 ( .A0(n28252), .A1(n27555), .B0(n28349), .C0(n27409), .Y(
        n27410) );
  OAI22XL U22278 ( .A0(n28186), .A1(n27553), .B0(n27557), .B1(n27431), .Y(
        n27409) );
  AOI211XL U22279 ( .A0(n28252), .A1(n27549), .B0(n28342), .C0(n27407), .Y(
        n27408) );
  OAI22XL U22280 ( .A0(n28186), .A1(n27547), .B0(n5916), .B1(n27546), .Y(
        n27407) );
  AOI211XL U22281 ( .A0(n28252), .A1(n27543), .B0(n28335), .C0(n27405), .Y(
        n27406) );
  OAI22XL U22282 ( .A0(n28186), .A1(n27541), .B0(n5825), .B1(n27545), .Y(
        n27405) );
  AOI211XL U22283 ( .A0(n28252), .A1(n27537), .B0(n28328), .C0(n27403), .Y(
        n27404) );
  OAI22XL U22284 ( .A0(n28186), .A1(n27535), .B0(n5916), .B1(n27534), .Y(
        n27403) );
  OAI22XL U22285 ( .A0(n28186), .A1(n27529), .B0(n27533), .B1(n27431), .Y(
        n27401) );
  AOI211XL U22286 ( .A0(n28252), .A1(n27811), .B0(n28625), .C0(n27494), .Y(
        n27495) );
  OAI22XL U22287 ( .A0(n28186), .A1(n27809), .B0(n27813), .B1(n28179), .Y(
        n27494) );
  AOI211XL U22288 ( .A0(n28252), .A1(n27805), .B0(n28625), .C0(n27492), .Y(
        n27493) );
  OAI22XL U22289 ( .A0(n28186), .A1(n27803), .B0(n5825), .B1(n27802), .Y(
        n27492) );
  OAI22XL U22290 ( .A0(n28186), .A1(n27523), .B0(n27522), .B1(n28179), .Y(
        n27399) );
  AOI211XL U22291 ( .A0(n28252), .A1(n27799), .B0(n28625), .C0(n27490), .Y(
        n27491) );
  OAI22XL U22292 ( .A0(n28186), .A1(n27797), .B0(n5916), .B1(n27796), .Y(
        n27490) );
  OAI22XL U22293 ( .A0(n28186), .A1(n27791), .B0(n5916), .B1(n27795), .Y(
        n27488) );
  AOI211XL U22294 ( .A0(n28252), .A1(n27787), .B0(n28625), .C0(n27486), .Y(
        n27487) );
  OAI22XL U22295 ( .A0(n28237), .A1(n27785), .B0(n5916), .B1(n27784), .Y(
        n27486) );
  AOI211XL U22296 ( .A0(n28252), .A1(n27781), .B0(n28625), .C0(n27484), .Y(
        n27485) );
  OAI22XL U22297 ( .A0(n28237), .A1(n27779), .B0(n5916), .B1(n27783), .Y(
        n27484) );
  AOI211XL U22298 ( .A0(n28252), .A1(n27775), .B0(n28625), .C0(n27482), .Y(
        n27483) );
  OAI22XL U22299 ( .A0(n28237), .A1(n27773), .B0(n27777), .B1(n28179), .Y(
        n27482) );
  AOI211XL U22300 ( .A0(n28252), .A1(n27768), .B0(n28625), .C0(n27480), .Y(
        n27481) );
  OAI22XL U22301 ( .A0(n28237), .A1(n27766), .B0(n5916), .B1(n7110), .Y(n27480) );
  AOI211XL U22302 ( .A0(n28252), .A1(n27762), .B0(n28625), .C0(n27478), .Y(
        n27479) );
  OAI22XL U22303 ( .A0(n28237), .A1(n27760), .B0(n5916), .B1(n27764), .Y(
        n27478) );
  AOI211XL U22304 ( .A0(n11929), .A1(n27756), .B0(n28625), .C0(n27476), .Y(
        n27477) );
  OAI22XL U22305 ( .A0(n28237), .A1(n27754), .B0(n5825), .B1(n27758), .Y(
        n27476) );
  AOI211XL U22306 ( .A0(n28252), .A1(n27750), .B0(n28625), .C0(n27474), .Y(
        n27475) );
  OAI22XL U22307 ( .A0(n28237), .A1(n27748), .B0(n27747), .B1(n28179), .Y(
        n27474) );
  AOI211XL U22308 ( .A0(n11929), .A1(n27744), .B0(n28557), .C0(n27472), .Y(
        n27473) );
  OAI22XL U22309 ( .A0(n28237), .A1(n27742), .B0(n28271), .B1(n27746), .Y(
        n27472) );
  AOI211XL U22310 ( .A0(n28252), .A1(n27519), .B0(n28306), .C0(n27397), .Y(
        n27398) );
  OAI22XL U22311 ( .A0(n28186), .A1(n27517), .B0(n27516), .B1(n28179), .Y(
        n27397) );
  AOI211XL U22312 ( .A0(n28252), .A1(n27738), .B0(n28550), .C0(n27470), .Y(
        n27471) );
  OAI22XL U22313 ( .A0(n28237), .A1(n27736), .B0(n7116), .B1(n28179), .Y(
        n27470) );
  AOI211XL U22314 ( .A0(n11929), .A1(n27732), .B0(n28543), .C0(n27468), .Y(
        n27469) );
  OAI22XL U22315 ( .A0(n28237), .A1(n27730), .B0(n27729), .B1(n28179), .Y(
        n27468) );
  AOI211XL U22316 ( .A0(n11929), .A1(n27726), .B0(n28536), .C0(n27466), .Y(
        n27467) );
  OAI22XL U22317 ( .A0(n28237), .A1(n27724), .B0(n5916), .B1(n27728), .Y(
        n27466) );
  AOI211XL U22318 ( .A0(n11929), .A1(n27720), .B0(n28529), .C0(n27464), .Y(
        n27465) );
  OAI22XL U22319 ( .A0(n28237), .A1(n27718), .B0(n5825), .B1(n27717), .Y(
        n27464) );
  OAI22XL U22320 ( .A0(n28237), .A1(n27712), .B0(n27711), .B1(n28179), .Y(
        n27462) );
  AOI211XL U22321 ( .A0(n11929), .A1(n27708), .B0(n28515), .C0(n27460), .Y(
        n27461) );
  OAI22XL U22322 ( .A0(n28237), .A1(n27706), .B0(n5825), .B1(n27710), .Y(
        n27460) );
  OAI22XL U22323 ( .A0(n28237), .A1(n27700), .B0(n27704), .B1(n28179), .Y(
        n27458) );
  OAI22XL U22324 ( .A0(n28237), .A1(n27694), .B0(n5825), .B1(n27698), .Y(
        n27456) );
  AOI211XL U22325 ( .A0(n28252), .A1(n27690), .B0(n28494), .C0(n27454), .Y(
        n27455) );
  OAI22XL U22326 ( .A0(n28237), .A1(n27688), .B0(n5916), .B1(n27692), .Y(
        n27454) );
  AOI211XL U22327 ( .A0(n28252), .A1(n27683), .B0(n28487), .C0(n27452), .Y(
        n27453) );
  OAI22XL U22328 ( .A0(n28237), .A1(n27681), .B0(n27685), .B1(n28179), .Y(
        n27452) );
  OAI22XL U22329 ( .A0(n28186), .A1(n27511), .B0(n27510), .B1(n27431), .Y(
        n27395) );
  AOI211XL U22330 ( .A0(n28252), .A1(n27677), .B0(n28480), .C0(n27450), .Y(
        n27451) );
  OAI22XL U22331 ( .A0(n28237), .A1(n27675), .B0(n5916), .B1(n27674), .Y(
        n27450) );
  AOI211XL U22332 ( .A0(n28252), .A1(n27671), .B0(n28473), .C0(n27448), .Y(
        n27449) );
  OAI22XL U22333 ( .A0(n28237), .A1(n27669), .B0(n27668), .B1(n28179), .Y(
        n27448) );
  OAI22XL U22334 ( .A0(n28237), .A1(n27663), .B0(n27662), .B1(n28179), .Y(
        n27446) );
  OAI22XL U22335 ( .A0(n28237), .A1(n27657), .B0(n5825), .B1(n27656), .Y(
        n27444) );
  AOI211XL U22336 ( .A0(n28252), .A1(n27653), .B0(n28452), .C0(n27442), .Y(
        n27443) );
  OAI22XL U22337 ( .A0(n28237), .A1(n27651), .B0(n27650), .B1(n28179), .Y(
        n27442) );
  AOI211XL U22338 ( .A0(n28252), .A1(n27647), .B0(n28452), .C0(n27440), .Y(
        n27441) );
  OAI22XL U22339 ( .A0(n28237), .A1(n27645), .B0(n5825), .B1(n27644), .Y(
        n27440) );
  AOI211XL U22340 ( .A0(n28252), .A1(n27641), .B0(n28452), .C0(n27438), .Y(
        n27439) );
  OAI22XL U22341 ( .A0(n28237), .A1(n27639), .B0(n5825), .B1(n27643), .Y(
        n27438) );
  AOI211XL U22342 ( .A0(n28252), .A1(n27635), .B0(n28452), .C0(n27436), .Y(
        n27437) );
  OAI22XL U22343 ( .A0(n28237), .A1(n27633), .B0(n27637), .B1(n28179), .Y(
        n27436) );
  AOI211XL U22344 ( .A0(n28252), .A1(n27628), .B0(n28452), .C0(n27434), .Y(
        n27435) );
  OAI22XL U22345 ( .A0(n28237), .A1(n27626), .B0(n27630), .B1(n28179), .Y(
        n27434) );
  AOI211XL U22346 ( .A0(n28252), .A1(n27622), .B0(n28452), .C0(n27432), .Y(
        n27433) );
  OAI22XL U22347 ( .A0(n28237), .A1(n27620), .B0(n5825), .B1(n7108), .Y(n27432) );
  OAI22XL U22348 ( .A0(n28186), .A1(n27505), .B0(n27504), .B1(n28179), .Y(
        n27393) );
  AOI211XL U22349 ( .A0(n28252), .A1(n27616), .B0(n28452), .C0(n27429), .Y(
        n27430) );
  OAI22XL U22350 ( .A0(n28237), .A1(n27614), .B0(n5825), .B1(n27613), .Y(
        n27429) );
  AOI211XL U22351 ( .A0(n28252), .A1(n27610), .B0(n28452), .C0(n27427), .Y(
        n27428) );
  OAI22XL U22352 ( .A0(n28237), .A1(n27608), .B0(n27607), .B1(n28179), .Y(
        n27427) );
  AOI211XL U22353 ( .A0(n28252), .A1(n27604), .B0(n28452), .C0(n27425), .Y(
        n27426) );
  OAI22XL U22354 ( .A0(n28237), .A1(n27602), .B0(n5825), .B1(n27601), .Y(
        n27425) );
  AOI211XL U22355 ( .A0(n28252), .A1(n27598), .B0(n28452), .C0(n27423), .Y(
        n27424) );
  OAI22XL U22356 ( .A0(n28237), .A1(n27596), .B0(n27595), .B1(n28179), .Y(
        n27423) );
  AOI211XL U22357 ( .A0(n28252), .A1(n27592), .B0(n28452), .C0(n27421), .Y(
        n27422) );
  OAI22XL U22358 ( .A0(n28237), .A1(n27590), .B0(n27589), .B1(n28179), .Y(
        n27421) );
  OAI22XL U22359 ( .A0(n28237), .A1(n27584), .B0(n5825), .B1(n27583), .Y(
        n27419) );
  OAI22XL U22360 ( .A0(n28237), .A1(n27578), .B0(n5825), .B1(n27582), .Y(
        n27417) );
  OAI22XL U22361 ( .A0(n28237), .A1(n27572), .B0(n5825), .B1(n7106), .Y(n27415) );
  AOI211XL U22362 ( .A0(n28252), .A1(n27568), .B0(n28364), .C0(n27413), .Y(
        n27414) );
  OAI22XL U22363 ( .A0(n28186), .A1(n27566), .B0(n27565), .B1(n27431), .Y(
        n27413) );
  AOI211XL U22364 ( .A0(n28252), .A1(n27562), .B0(n28357), .C0(n27411), .Y(
        n27412) );
  OAI22XL U22365 ( .A0(n28186), .A1(n27559), .B0(n27564), .B1(n27431), .Y(
        n27411) );
  AOI211XL U22366 ( .A0(n28252), .A1(n27501), .B0(n7120), .C0(n27391), .Y(
        n27392) );
  OAI22XL U22367 ( .A0(n28186), .A1(n27499), .B0(n27503), .B1(n27431), .Y(
        n27391) );
  NOR2XL U22368 ( .A(n11991), .B(n11983), .Y(A4_WEN) );
  AOI211XL U22369 ( .A0(n27631), .A1(n27555), .B0(n28349), .C0(n27554), .Y(
        n27556) );
  OAI22XL U22370 ( .A0(n27560), .A1(n27553), .B0(n28295), .B1(n27552), .Y(
        n27554) );
  AOI211XL U22371 ( .A0(n27631), .A1(n27549), .B0(n28342), .C0(n27548), .Y(
        n27550) );
  OAI22XL U22372 ( .A0(n27560), .A1(n27547), .B0(n28295), .B1(n27546), .Y(
        n27548) );
  AOI211XL U22373 ( .A0(n5827), .A1(n27543), .B0(n28335), .C0(n27542), .Y(
        n27544) );
  OAI22XL U22374 ( .A0(n28579), .A1(n27541), .B0(n27540), .B1(n27686), .Y(
        n27542) );
  AOI211XL U22375 ( .A0(n27631), .A1(n27537), .B0(n28328), .C0(n27536), .Y(
        n27538) );
  OAI22XL U22376 ( .A0(n28579), .A1(n27529), .B0(n28295), .B1(n27528), .Y(
        n27530) );
  AOI211XL U22377 ( .A0(n27631), .A1(n27811), .B0(n28625), .C0(n27810), .Y(
        n27812) );
  AOI211XL U22378 ( .A0(n27631), .A1(n27805), .B0(n28625), .C0(n27804), .Y(
        n27806) );
  OAI22XL U22379 ( .A0(n28579), .A1(n27523), .B0(n27522), .B1(n28353), .Y(
        n27524) );
  AOI211XL U22380 ( .A0(n27631), .A1(n27799), .B0(n28625), .C0(n27798), .Y(
        n27800) );
  OAI22XL U22381 ( .A0(n28579), .A1(n27791), .B0(n27790), .B1(n28353), .Y(
        n27792) );
  AOI211XL U22382 ( .A0(n27631), .A1(n27787), .B0(n28625), .C0(n27786), .Y(
        n27788) );
  AOI211XL U22383 ( .A0(n27631), .A1(n27781), .B0(n28625), .C0(n27780), .Y(
        n27782) );
  OAI22XL U22384 ( .A0(n28579), .A1(n27779), .B0(n27778), .B1(n28353), .Y(
        n27780) );
  AOI211XL U22385 ( .A0(n27631), .A1(n27775), .B0(n28625), .C0(n27774), .Y(
        n27776) );
  AOI211XL U22386 ( .A0(n27631), .A1(n27768), .B0(n28625), .C0(n27767), .Y(
        n27769) );
  OAI22XL U22387 ( .A0(n28579), .A1(n27766), .B0(n27765), .B1(n28353), .Y(
        n27767) );
  AOI211XL U22388 ( .A0(n27631), .A1(n27762), .B0(n28625), .C0(n27761), .Y(
        n27763) );
  OAI22XL U22389 ( .A0(n28579), .A1(n27760), .B0(n27759), .B1(n28353), .Y(
        n27761) );
  AOI211XL U22390 ( .A0(n27631), .A1(n27756), .B0(n28625), .C0(n27755), .Y(
        n27757) );
  OAI22XL U22391 ( .A0(n28579), .A1(n27754), .B0(n27753), .B1(n28353), .Y(
        n27755) );
  AOI211XL U22392 ( .A0(n27631), .A1(n27750), .B0(n28625), .C0(n27749), .Y(
        n27751) );
  OAI22XL U22393 ( .A0(n28579), .A1(n27748), .B0(n27747), .B1(n28353), .Y(
        n27749) );
  OAI22XL U22394 ( .A0(n28579), .A1(n27742), .B0(n27741), .B1(n28353), .Y(
        n27743) );
  AOI211XL U22395 ( .A0(n27631), .A1(n27519), .B0(n28306), .C0(n27518), .Y(
        n27520) );
  OAI22XL U22396 ( .A0(n28579), .A1(n27517), .B0(n27516), .B1(n28353), .Y(
        n27518) );
  AOI211XL U22397 ( .A0(n27631), .A1(n27738), .B0(n28550), .C0(n27737), .Y(
        n27739) );
  OAI22XL U22398 ( .A0(n28579), .A1(n27730), .B0(n27729), .B1(n28353), .Y(
        n27731) );
  AOI211XL U22399 ( .A0(n27631), .A1(n27726), .B0(n28536), .C0(n27725), .Y(
        n27727) );
  OAI22XL U22400 ( .A0(n28579), .A1(n27724), .B0(n27723), .B1(n28353), .Y(
        n27725) );
  AOI211XL U22401 ( .A0(n27631), .A1(n27720), .B0(n28529), .C0(n27719), .Y(
        n27721) );
  OAI22XL U22402 ( .A0(n28579), .A1(n27712), .B0(n27711), .B1(n28353), .Y(
        n27713) );
  OAI22XL U22403 ( .A0(n28579), .A1(n27706), .B0(n27705), .B1(n28353), .Y(
        n27707) );
  OAI22XL U22404 ( .A0(n28579), .A1(n27694), .B0(n27693), .B1(n28353), .Y(
        n27695) );
  AOI211XL U22405 ( .A0(n5798), .A1(n27690), .B0(n28494), .C0(n27689), .Y(
        n27691) );
  OAI22XL U22406 ( .A0(n28579), .A1(n27688), .B0(n27687), .B1(n27686), .Y(
        n27689) );
  AOI211XL U22407 ( .A0(n5827), .A1(n27683), .B0(n28487), .C0(n27682), .Y(
        n27684) );
  OAI22XL U22408 ( .A0(n27560), .A1(n27511), .B0(n27510), .B1(n28353), .Y(
        n27512) );
  AOI211XL U22409 ( .A0(n5798), .A1(n27677), .B0(n28480), .C0(n27676), .Y(
        n27678) );
  AOI211XL U22410 ( .A0(n27631), .A1(n27671), .B0(n28473), .C0(n27670), .Y(
        n27672) );
  OAI22XL U22411 ( .A0(n28579), .A1(n27669), .B0(n27668), .B1(n28353), .Y(
        n27670) );
  OAI22XL U22412 ( .A0(n28579), .A1(n27663), .B0(n27662), .B1(n28353), .Y(
        n27664) );
  AOI211XL U22413 ( .A0(n27631), .A1(n27653), .B0(n28452), .C0(n27652), .Y(
        n27654) );
  OAI22XL U22414 ( .A0(n28579), .A1(n27651), .B0(n27650), .B1(n28353), .Y(
        n27652) );
  AOI211XL U22415 ( .A0(n27631), .A1(n27647), .B0(n28452), .C0(n27646), .Y(
        n27648) );
  AOI211XL U22416 ( .A0(n5827), .A1(n27641), .B0(n28452), .C0(n27640), .Y(
        n27642) );
  OAI22XL U22417 ( .A0(n28579), .A1(n27639), .B0(n27638), .B1(n27686), .Y(
        n27640) );
  AOI211XL U22418 ( .A0(n27631), .A1(n27635), .B0(n28452), .C0(n27634), .Y(
        n27636) );
  AOI211XL U22419 ( .A0(n27631), .A1(n27628), .B0(n28452), .C0(n27627), .Y(
        n27629) );
  AOI211XL U22420 ( .A0(n5827), .A1(n27622), .B0(n28452), .C0(n27621), .Y(
        n27623) );
  OAI22XL U22421 ( .A0(n28579), .A1(n27620), .B0(n27619), .B1(n28353), .Y(
        n27621) );
  OAI22XL U22422 ( .A0(n28579), .A1(n27505), .B0(n27504), .B1(n28353), .Y(
        n27506) );
  AOI211XL U22423 ( .A0(n5918), .A1(n27616), .B0(n28452), .C0(n27615), .Y(
        n27617) );
  AOI211XL U22424 ( .A0(n27631), .A1(n27610), .B0(n28452), .C0(n27609), .Y(
        n27611) );
  OAI22XL U22425 ( .A0(n28579), .A1(n27608), .B0(n27607), .B1(n27686), .Y(
        n27609) );
  AOI211XL U22426 ( .A0(n5918), .A1(n27604), .B0(n28452), .C0(n27603), .Y(
        n27605) );
  AOI211XL U22427 ( .A0(n5918), .A1(n27598), .B0(n28452), .C0(n27597), .Y(
        n27599) );
  OAI22XL U22428 ( .A0(n28579), .A1(n27596), .B0(n27595), .B1(n27686), .Y(
        n27597) );
  AOI211XL U22429 ( .A0(n5918), .A1(n27592), .B0(n28452), .C0(n27591), .Y(
        n27593) );
  OAI22XL U22430 ( .A0(n28579), .A1(n27590), .B0(n27589), .B1(n28353), .Y(
        n27591) );
  OAI22XL U22431 ( .A0(n28579), .A1(n27584), .B0(n28295), .B1(n27583), .Y(
        n27585) );
  OAI22XL U22432 ( .A0(n28579), .A1(n27578), .B0(n27577), .B1(n28353), .Y(
        n27579) );
  OAI22XL U22433 ( .A0(n28579), .A1(n27572), .B0(n27571), .B1(n28353), .Y(
        n27573) );
  AOI211XL U22434 ( .A0(n27631), .A1(n27568), .B0(n28364), .C0(n27567), .Y(
        n27569) );
  OAI22XL U22435 ( .A0(n28579), .A1(n27566), .B0(n27565), .B1(n28353), .Y(
        n27567) );
  AOI211XL U22436 ( .A0(n27631), .A1(n27562), .B0(n28357), .C0(n27561), .Y(
        n27563) );
  OAI22XL U22437 ( .A0(n27560), .A1(n27559), .B0(n28295), .B1(n27558), .Y(
        n27561) );
  NOR2XL U22438 ( .A(n11989), .B(n11987), .Y(A3_WEN) );
  AOI211XL U22439 ( .A0(n27162), .A1(n28350), .B0(n28349), .C0(n27853), .Y(
        n27854) );
  OAI22XL U22440 ( .A0(n27959), .A1(n28347), .B0(n28352), .B1(n7140), .Y(
        n27853) );
  AOI211XL U22441 ( .A0(n27162), .A1(n28343), .B0(n28342), .C0(n27849), .Y(
        n27850) );
  OAI22XL U22442 ( .A0(n27959), .A1(n28340), .B0(n28345), .B1(n28050), .Y(
        n27849) );
  AOI211XL U22443 ( .A0(n27162), .A1(n28336), .B0(n28335), .C0(n27845), .Y(
        n27846) );
  OAI22XL U22444 ( .A0(n27959), .A1(n28333), .B0(n28338), .B1(n5823), .Y(
        n27845) );
  AOI211XL U22445 ( .A0(n27162), .A1(n28329), .B0(n28328), .C0(n27841), .Y(
        n27842) );
  OAI22XL U22446 ( .A0(n27959), .A1(n28326), .B0(n28331), .B1(n7140), .Y(
        n27841) );
  OAI22XL U22447 ( .A0(n27959), .A1(n28318), .B0(n28324), .B1(n28050), .Y(
        n27837) );
  AOI211XL U22448 ( .A0(n27162), .A1(n28626), .B0(n28625), .C0(n28056), .Y(
        n28057) );
  OAI22XL U22449 ( .A0(n28055), .A1(n28623), .B0(n28622), .B1(n28054), .Y(
        n28056) );
  AOI211XL U22450 ( .A0(n27162), .A1(n28619), .B0(n28625), .C0(n28048), .Y(
        n28049) );
  OAI22XL U22451 ( .A0(n28055), .A1(n28617), .B0(n28621), .B1(n5823), .Y(
        n28048) );
  OAI22XL U22452 ( .A0(n27959), .A1(n28311), .B0(n28316), .B1(n28050), .Y(
        n27833) );
  OAI22XL U22453 ( .A0(n28055), .A1(n28611), .B0(n28615), .B1(n5823), .Y(
        n28043) );
  AOI211XL U22454 ( .A0(n27162), .A1(n28607), .B0(n28625), .C0(n28038), .Y(
        n28039) );
  OAI22XL U22455 ( .A0(n28055), .A1(n28605), .B0(n28604), .B1(n7140), .Y(
        n28038) );
  AOI211XL U22456 ( .A0(n27162), .A1(n28601), .B0(n28625), .C0(n28033), .Y(
        n28034) );
  OAI22XL U22457 ( .A0(n27959), .A1(n28599), .B0(n28598), .B1(n7140), .Y(
        n28033) );
  AOI211XL U22458 ( .A0(n27162), .A1(n28595), .B0(n28625), .C0(n28028), .Y(
        n28029) );
  OAI22XL U22459 ( .A0(n28055), .A1(n28593), .B0(n28592), .B1(n7140), .Y(
        n28028) );
  AOI211XL U22460 ( .A0(n5826), .A1(n28589), .B0(n28625), .C0(n28023), .Y(
        n28024) );
  OAI22XL U22461 ( .A0(n28055), .A1(n28587), .B0(n28591), .B1(n7140), .Y(
        n28023) );
  AOI211XL U22462 ( .A0(n5826), .A1(n28583), .B0(n28625), .C0(n28018), .Y(
        n28019) );
  OAI22XL U22463 ( .A0(n28055), .A1(n28581), .B0(n28580), .B1(n5823), .Y(
        n28018) );
  AOI211XL U22464 ( .A0(n27162), .A1(n28576), .B0(n28625), .C0(n28013), .Y(
        n28014) );
  OAI22XL U22465 ( .A0(n27959), .A1(n28574), .B0(n28573), .B1(n7140), .Y(
        n28013) );
  AOI211XL U22466 ( .A0(n27162), .A1(n28570), .B0(n28625), .C0(n28008), .Y(
        n28009) );
  OAI22XL U22467 ( .A0(n27959), .A1(n28568), .B0(n28567), .B1(n7140), .Y(
        n28008) );
  AOI211XL U22468 ( .A0(n27162), .A1(n28564), .B0(n28625), .C0(n28003), .Y(
        n28004) );
  OAI22XL U22469 ( .A0(n27959), .A1(n28562), .B0(n28566), .B1(n5823), .Y(
        n28003) );
  AOI211XL U22470 ( .A0(n27162), .A1(n28558), .B0(n28557), .C0(n27998), .Y(
        n27999) );
  OAI22XL U22471 ( .A0(n27959), .A1(n28555), .B0(n28560), .B1(n5823), .Y(
        n27998) );
  AOI211XL U22472 ( .A0(n27162), .A1(n28307), .B0(n28306), .C0(n27829), .Y(
        n27830) );
  OAI22XL U22473 ( .A0(n27959), .A1(n28304), .B0(n28303), .B1(n5823), .Y(
        n27829) );
  AOI211XL U22474 ( .A0(n27162), .A1(n28551), .B0(n28550), .C0(n27993), .Y(
        n27994) );
  OAI22XL U22475 ( .A0(n27959), .A1(n28548), .B0(n28547), .B1(n7140), .Y(
        n27993) );
  AOI211XL U22476 ( .A0(n5826), .A1(n28544), .B0(n28543), .C0(n27988), .Y(
        n27989) );
  OAI22XL U22477 ( .A0(n27959), .A1(n28541), .B0(n28546), .B1(n7140), .Y(
        n27988) );
  AOI211XL U22478 ( .A0(n5826), .A1(n28537), .B0(n28536), .C0(n27983), .Y(
        n27984) );
  OAI22XL U22479 ( .A0(n27959), .A1(n28534), .B0(n28533), .B1(n5823), .Y(
        n27983) );
  AOI211XL U22480 ( .A0(n5826), .A1(n28530), .B0(n28529), .C0(n27978), .Y(
        n27979) );
  OAI22XL U22481 ( .A0(n27959), .A1(n28527), .B0(n28526), .B1(n5823), .Y(
        n27978) );
  OAI22XL U22482 ( .A0(n27959), .A1(n28520), .B0(n28519), .B1(n5823), .Y(
        n27973) );
  AOI211XL U22483 ( .A0(n5826), .A1(n28516), .B0(n28515), .C0(n27969), .Y(
        n27970) );
  OAI22XL U22484 ( .A0(n27959), .A1(n28513), .B0(n28512), .B1(n7140), .Y(
        n27969) );
  OAI22XL U22485 ( .A0(n27959), .A1(n28506), .B0(n28505), .B1(n5823), .Y(
        n27965) );
  OAI22XL U22486 ( .A0(n27959), .A1(n28499), .B0(n28504), .B1(n28050), .Y(
        n27961) );
  OAI22XL U22487 ( .A0(n27959), .A1(n28492), .B0(n28497), .B1(n7140), .Y(
        n27956) );
  AOI211XL U22488 ( .A0(n27162), .A1(n28488), .B0(n28487), .C0(n27952), .Y(
        n27953) );
  OAI22XL U22489 ( .A0(n27959), .A1(n28485), .B0(n28484), .B1(n5823), .Y(
        n27952) );
  OAI22XL U22490 ( .A0(n27959), .A1(n28297), .B0(n28296), .B1(n5823), .Y(
        n27825) );
  AOI211XL U22491 ( .A0(n27162), .A1(n28481), .B0(n28480), .C0(n27948), .Y(
        n27949) );
  OAI22XL U22492 ( .A0(n27959), .A1(n28478), .B0(n28477), .B1(n5823), .Y(
        n27948) );
  AOI211XL U22493 ( .A0(n27162), .A1(n28474), .B0(n28473), .C0(n27944), .Y(
        n27945) );
  OAI22XL U22494 ( .A0(n27959), .A1(n28471), .B0(n28470), .B1(n5823), .Y(
        n27944) );
  OAI22XL U22495 ( .A0(n27959), .A1(n28464), .B0(n28469), .B1(n7140), .Y(
        n27940) );
  OAI22XL U22496 ( .A0(n27959), .A1(n28457), .B0(n28462), .B1(n7140), .Y(
        n27936) );
  AOI211XL U22497 ( .A0(n27162), .A1(n28453), .B0(n28452), .C0(n27932), .Y(
        n27933) );
  OAI22XL U22498 ( .A0(n27959), .A1(n28450), .B0(n28449), .B1(n5823), .Y(
        n27932) );
  AOI211XL U22499 ( .A0(n27162), .A1(n28446), .B0(n28452), .C0(n27927), .Y(
        n27928) );
  OAI22XL U22500 ( .A0(n27959), .A1(n28444), .B0(n28443), .B1(n7140), .Y(
        n27927) );
  AOI211XL U22501 ( .A0(n27162), .A1(n28440), .B0(n28452), .C0(n27922), .Y(
        n27923) );
  OAI22XL U22502 ( .A0(n27959), .A1(n28438), .B0(n28437), .B1(n7140), .Y(
        n27922) );
  AOI211XL U22503 ( .A0(n5826), .A1(n28434), .B0(n28452), .C0(n27917), .Y(
        n27918) );
  OAI22XL U22504 ( .A0(n27959), .A1(n28432), .B0(n28436), .B1(n5823), .Y(
        n27917) );
  AOI211XL U22505 ( .A0(n5826), .A1(n28428), .B0(n28452), .C0(n27912), .Y(
        n27913) );
  OAI22XL U22506 ( .A0(n27959), .A1(n28426), .B0(n28425), .B1(n5823), .Y(
        n27912) );
  OAI22XL U22507 ( .A0(n27959), .A1(n28420), .B0(n28419), .B1(n5823), .Y(
        n27907) );
  OAI22XL U22508 ( .A0(n27959), .A1(n28289), .B0(n28294), .B1(n5823), .Y(
        n27821) );
  OAI22XL U22509 ( .A0(n27959), .A1(n28414), .B0(n28418), .B1(n7140), .Y(
        n27902) );
  AOI211XL U22510 ( .A0(n27162), .A1(n28410), .B0(n28452), .C0(n27897), .Y(
        n27898) );
  OAI22XL U22511 ( .A0(n27959), .A1(n28408), .B0(n28412), .B1(n5823), .Y(
        n27897) );
  AOI211XL U22512 ( .A0(n5826), .A1(n28404), .B0(n28452), .C0(n27892), .Y(
        n27893) );
  OAI22XL U22513 ( .A0(n27959), .A1(n28402), .B0(n28401), .B1(n7140), .Y(
        n27892) );
  AOI211XL U22514 ( .A0(n27162), .A1(n28398), .B0(n28452), .C0(n27887), .Y(
        n27888) );
  OAI22XL U22515 ( .A0(n27959), .A1(n28396), .B0(n28400), .B1(n5823), .Y(
        n27887) );
  AOI211XL U22516 ( .A0(n27162), .A1(n28392), .B0(n28452), .C0(n27882), .Y(
        n27883) );
  OAI22XL U22517 ( .A0(n27959), .A1(n28390), .B0(n28389), .B1(n5823), .Y(
        n27882) );
  OAI22XL U22518 ( .A0(n27959), .A1(n28383), .B0(n28388), .B1(n7140), .Y(
        n27877) );
  OAI22XL U22519 ( .A0(n27959), .A1(n28376), .B0(n28381), .B1(n7140), .Y(
        n27872) );
  OAI22XL U22520 ( .A0(n27959), .A1(n28369), .B0(n28368), .B1(n5823), .Y(
        n27867) );
  AOI211XL U22521 ( .A0(n27162), .A1(n28365), .B0(n28364), .C0(n27862), .Y(
        n27863) );
  OAI22XL U22522 ( .A0(n27959), .A1(n28362), .B0(n28367), .B1(n7140), .Y(
        n27862) );
  AOI211XL U22523 ( .A0(n5826), .A1(n28358), .B0(n28357), .C0(n27857), .Y(
        n27858) );
  OAI22XL U22524 ( .A0(n27959), .A1(n28355), .B0(n28354), .B1(n5823), .Y(
        n27857) );
  AOI211XL U22525 ( .A0(n5826), .A1(n28285), .B0(n7120), .C0(n27817), .Y(
        n27818) );
  OAI22XL U22526 ( .A0(n27959), .A1(n28282), .B0(n28281), .B1(n7140), .Y(
        n27817) );
  AOI22XL U22527 ( .A0(Q2_addr[7]), .A1(n27205), .B0(Q3_addr[7]), .B1(n27088), 
        .Y(n15039) );
  AOI22XL U22528 ( .A0(Q2_addr[6]), .A1(n27205), .B0(Q3_addr[6]), .B1(n27088), 
        .Y(n15032) );
  AOI21XL U22529 ( .A0(n27162), .A1(Q0_addr[6]), .B0(n15031), .Y(n15033) );
  AOI22XL U22530 ( .A0(Q2_addr[5]), .A1(n27205), .B0(Q3_addr[5]), .B1(n27088), 
        .Y(n15029) );
  AOI22XL U22531 ( .A0(Q2_addr[4]), .A1(n27205), .B0(Q3_addr[4]), .B1(n27088), 
        .Y(n15004) );
  AOI22XL U22532 ( .A0(Q2_addr[3]), .A1(n27205), .B0(Q3_addr[3]), .B1(n27088), 
        .Y(n14989) );
  AOI22XL U22533 ( .A0(Q2_addr[2]), .A1(n27205), .B0(Q3_addr[2]), .B1(n27088), 
        .Y(n14986) );
  AOI22XL U22534 ( .A0(Q2_addr[1]), .A1(n27205), .B0(Q3_addr[1]), .B1(n27088), 
        .Y(n14984) );
  AOI22XL U22535 ( .A0(Q3_addr[0]), .A1(n27088), .B0(Q2_addr[0]), .B1(n27205), 
        .Y(n14982) );
  NOR2XL U22536 ( .A(n11989), .B(n11981), .Y(A2_WEN) );
  AOI211XL U22537 ( .A0(n28143), .A1(n28350), .B0(n28349), .C0(n28077), .Y(
        n28078) );
  OAI22XL U22538 ( .A0(n28125), .A1(n28347), .B0(n28346), .B1(n28118), .Y(
        n28077) );
  AOI211XL U22539 ( .A0(n28143), .A1(n28343), .B0(n28342), .C0(n28075), .Y(
        n28076) );
  OAI22XL U22540 ( .A0(n28125), .A1(n28340), .B0(n28339), .B1(n28118), .Y(
        n28075) );
  AOI211XL U22541 ( .A0(n28143), .A1(n28336), .B0(n28335), .C0(n28073), .Y(
        n28074) );
  OAI22XL U22542 ( .A0(n28125), .A1(n28333), .B0(n28332), .B1(n28068), .Y(
        n28073) );
  AOI211XL U22543 ( .A0(n28143), .A1(n28329), .B0(n28328), .C0(n28071), .Y(
        n28072) );
  OAI22XL U22544 ( .A0(n28125), .A1(n28326), .B0(n28325), .B1(n28118), .Y(
        n28071) );
  OAI22XL U22545 ( .A0(n28125), .A1(n28318), .B0(n28324), .B1(n28068), .Y(
        n28069) );
  AOI211XL U22546 ( .A0(n28143), .A1(n28626), .B0(n28625), .C0(n28169), .Y(
        n28170) );
  OAI22XL U22547 ( .A0(n28168), .A1(n28623), .B0(n28622), .B1(n28093), .Y(
        n28169) );
  AOI211XL U22548 ( .A0(n28143), .A1(n28619), .B0(n28625), .C0(n28166), .Y(
        n28167) );
  OAI22XL U22549 ( .A0(n28168), .A1(n28617), .B0(n28621), .B1(n28158), .Y(
        n28166) );
  OAI22XL U22550 ( .A0(n28125), .A1(n28311), .B0(n28316), .B1(n28068), .Y(
        n28066) );
  AOI211XL U22551 ( .A0(n28143), .A1(n28613), .B0(n28625), .C0(n28163), .Y(
        n28164) );
  OAI22XL U22552 ( .A0(n28125), .A1(n28611), .B0(n28610), .B1(n28068), .Y(
        n28163) );
  AOI211XL U22553 ( .A0(n28143), .A1(n28607), .B0(n28625), .C0(n28161), .Y(
        n28162) );
  OAI22XL U22554 ( .A0(n28168), .A1(n28605), .B0(n28609), .B1(n28118), .Y(
        n28161) );
  AOI211XL U22555 ( .A0(n28143), .A1(n28601), .B0(n28625), .C0(n28159), .Y(
        n28160) );
  OAI22XL U22556 ( .A0(n28168), .A1(n28599), .B0(n28603), .B1(n28093), .Y(
        n28159) );
  AOI211XL U22557 ( .A0(n28143), .A1(n28595), .B0(n28625), .C0(n28156), .Y(
        n28157) );
  OAI22XL U22558 ( .A0(n28168), .A1(n28593), .B0(n28592), .B1(n28068), .Y(
        n28156) );
  AOI211XL U22559 ( .A0(n28143), .A1(n28589), .B0(n28625), .C0(n28154), .Y(
        n28155) );
  OAI22XL U22560 ( .A0(n28125), .A1(n28587), .B0(n28586), .B1(n28138), .Y(
        n28154) );
  AOI211XL U22561 ( .A0(n28143), .A1(n28583), .B0(n28625), .C0(n28152), .Y(
        n28153) );
  OAI22XL U22562 ( .A0(n28168), .A1(n28581), .B0(n28585), .B1(n28068), .Y(
        n28152) );
  AOI211XL U22563 ( .A0(n28143), .A1(n28576), .B0(n28625), .C0(n28150), .Y(
        n28151) );
  OAI22XL U22564 ( .A0(n28125), .A1(n28574), .B0(n28578), .B1(n28165), .Y(
        n28150) );
  AOI211XL U22565 ( .A0(n28143), .A1(n28570), .B0(n28625), .C0(n28148), .Y(
        n28149) );
  OAI22XL U22566 ( .A0(n28125), .A1(n28568), .B0(n28567), .B1(n28068), .Y(
        n28148) );
  AOI211XL U22567 ( .A0(n28143), .A1(n28564), .B0(n28625), .C0(n28146), .Y(
        n28147) );
  OAI22XL U22568 ( .A0(n28125), .A1(n28562), .B0(n28561), .B1(n28068), .Y(
        n28146) );
  AOI211XL U22569 ( .A0(n28143), .A1(n28558), .B0(n28557), .C0(n28144), .Y(
        n28145) );
  OAI22XL U22570 ( .A0(n28125), .A1(n28555), .B0(n28560), .B1(n28118), .Y(
        n28144) );
  AOI211XL U22571 ( .A0(n28143), .A1(n28307), .B0(n28306), .C0(n28064), .Y(
        n28065) );
  OAI22XL U22572 ( .A0(n28125), .A1(n28304), .B0(n28309), .B1(n28068), .Y(
        n28064) );
  AOI211XL U22573 ( .A0(n28143), .A1(n28551), .B0(n28550), .C0(n28141), .Y(
        n28142) );
  OAI22XL U22574 ( .A0(n28125), .A1(n28548), .B0(n28553), .B1(n28138), .Y(
        n28141) );
  AOI211XL U22575 ( .A0(n28143), .A1(n28544), .B0(n28543), .C0(n28139), .Y(
        n28140) );
  OAI22XL U22576 ( .A0(n28125), .A1(n28541), .B0(n28540), .B1(n28138), .Y(
        n28139) );
  AOI211XL U22577 ( .A0(n28143), .A1(n28537), .B0(n28536), .C0(n28136), .Y(
        n28137) );
  OAI22XL U22578 ( .A0(n28168), .A1(n28534), .B0(n28539), .B1(n28068), .Y(
        n28136) );
  AOI211XL U22579 ( .A0(n28143), .A1(n28530), .B0(n28529), .C0(n28134), .Y(
        n28135) );
  OAI22XL U22580 ( .A0(n28125), .A1(n28527), .B0(n28532), .B1(n28068), .Y(
        n28134) );
  OAI22XL U22581 ( .A0(n28125), .A1(n28520), .B0(n28519), .B1(n28118), .Y(
        n28132) );
  AOI211XL U22582 ( .A0(n28143), .A1(n28516), .B0(n28515), .C0(n28130), .Y(
        n28131) );
  OAI22XL U22583 ( .A0(n28125), .A1(n28513), .B0(n28518), .B1(n28165), .Y(
        n28130) );
  OAI22XL U22584 ( .A0(n28125), .A1(n28506), .B0(n28511), .B1(n28068), .Y(
        n28128) );
  OAI22XL U22585 ( .A0(n28125), .A1(n28499), .B0(n28498), .B1(n28158), .Y(
        n28126) );
  AOI211XL U22586 ( .A0(n28143), .A1(n28495), .B0(n28494), .C0(n28123), .Y(
        n28124) );
  OAI22XL U22587 ( .A0(n28125), .A1(n28492), .B0(n28497), .B1(n28068), .Y(
        n28123) );
  AOI211XL U22588 ( .A0(n28143), .A1(n28488), .B0(n28487), .C0(n28121), .Y(
        n28122) );
  OAI22XL U22589 ( .A0(n28125), .A1(n28485), .B0(n28484), .B1(n28138), .Y(
        n28121) );
  OAI22XL U22590 ( .A0(n28125), .A1(n28297), .B0(n28296), .B1(n28165), .Y(
        n28062) );
  AOI211XL U22591 ( .A0(n28143), .A1(n28481), .B0(n28480), .C0(n28119), .Y(
        n28120) );
  OAI22XL U22592 ( .A0(n28125), .A1(n28478), .B0(n28477), .B1(n28118), .Y(
        n28119) );
  AOI211XL U22593 ( .A0(n28143), .A1(n28474), .B0(n28473), .C0(n28116), .Y(
        n28117) );
  OAI22XL U22594 ( .A0(n28125), .A1(n28471), .B0(n28470), .B1(n28118), .Y(
        n28116) );
  OAI22XL U22595 ( .A0(n28168), .A1(n28464), .B0(n28463), .B1(n28118), .Y(
        n28114) );
  OAI22XL U22596 ( .A0(n28125), .A1(n28457), .B0(n28462), .B1(n28068), .Y(
        n28112) );
  AOI211XL U22597 ( .A0(n28143), .A1(n28453), .B0(n28452), .C0(n28110), .Y(
        n28111) );
  OAI22XL U22598 ( .A0(n28168), .A1(n28450), .B0(n28455), .B1(n28068), .Y(
        n28110) );
  AOI211XL U22599 ( .A0(n28143), .A1(n28446), .B0(n28452), .C0(n28108), .Y(
        n28109) );
  OAI22XL U22600 ( .A0(n28168), .A1(n28444), .B0(n28443), .B1(n28068), .Y(
        n28108) );
  AOI211XL U22601 ( .A0(n28143), .A1(n28440), .B0(n28452), .C0(n28106), .Y(
        n28107) );
  OAI22XL U22602 ( .A0(n28168), .A1(n28438), .B0(n28442), .B1(n28118), .Y(
        n28106) );
  AOI211XL U22603 ( .A0(n28143), .A1(n28434), .B0(n28452), .C0(n28104), .Y(
        n28105) );
  OAI22XL U22604 ( .A0(n28168), .A1(n28432), .B0(n28431), .B1(n28068), .Y(
        n28104) );
  AOI211XL U22605 ( .A0(n28143), .A1(n28428), .B0(n28452), .C0(n28102), .Y(
        n28103) );
  OAI22XL U22606 ( .A0(n28168), .A1(n28426), .B0(n28430), .B1(n28068), .Y(
        n28102) );
  AOI211XL U22607 ( .A0(n28143), .A1(n28422), .B0(n28452), .C0(n28100), .Y(
        n28101) );
  OAI22XL U22608 ( .A0(n28168), .A1(n28420), .B0(n28419), .B1(n28118), .Y(
        n28100) );
  OAI22XL U22609 ( .A0(n28125), .A1(n28289), .B0(n28288), .B1(n28068), .Y(
        n28060) );
  AOI211XL U22610 ( .A0(n28143), .A1(n28416), .B0(n28452), .C0(n28098), .Y(
        n28099) );
  OAI22XL U22611 ( .A0(n28125), .A1(n28414), .B0(n28418), .B1(n28068), .Y(
        n28098) );
  AOI211XL U22612 ( .A0(n28143), .A1(n28410), .B0(n28452), .C0(n28096), .Y(
        n28097) );
  OAI22XL U22613 ( .A0(n28125), .A1(n28408), .B0(n28412), .B1(n28118), .Y(
        n28096) );
  AOI211XL U22614 ( .A0(n28143), .A1(n28404), .B0(n28452), .C0(n28094), .Y(
        n28095) );
  OAI22XL U22615 ( .A0(n28125), .A1(n28402), .B0(n28406), .B1(n28118), .Y(
        n28094) );
  AOI211XL U22616 ( .A0(n28143), .A1(n28398), .B0(n28452), .C0(n28091), .Y(
        n28092) );
  OAI22XL U22617 ( .A0(n28125), .A1(n28396), .B0(n28395), .B1(n28068), .Y(
        n28091) );
  AOI211XL U22618 ( .A0(n28143), .A1(n28392), .B0(n28452), .C0(n28089), .Y(
        n28090) );
  OAI22XL U22619 ( .A0(n28125), .A1(n28390), .B0(n28389), .B1(n28118), .Y(
        n28089) );
  OAI22XL U22620 ( .A0(n28125), .A1(n28383), .B0(n28388), .B1(n28068), .Y(
        n28087) );
  OAI22XL U22621 ( .A0(n28125), .A1(n28376), .B0(n28381), .B1(n28068), .Y(
        n28085) );
  OAI22XL U22622 ( .A0(n28125), .A1(n28369), .B0(n28374), .B1(n28068), .Y(
        n28083) );
  AOI211XL U22623 ( .A0(n28143), .A1(n28365), .B0(n28364), .C0(n28081), .Y(
        n28082) );
  OAI22XL U22624 ( .A0(n28125), .A1(n28362), .B0(n28367), .B1(n28068), .Y(
        n28081) );
  AOI211XL U22625 ( .A0(n28143), .A1(n28358), .B0(n28357), .C0(n28079), .Y(
        n28080) );
  OAI22XL U22626 ( .A0(n28125), .A1(n28355), .B0(n28354), .B1(n28118), .Y(
        n28079) );
  AOI211XL U22627 ( .A0(n28143), .A1(n28285), .B0(n7120), .C0(n28058), .Y(
        n28059) );
  OAI22XL U22628 ( .A0(n28125), .A1(n28282), .B0(n28287), .B1(n28158), .Y(
        n28058) );
  AOI22XL U22629 ( .A0(n15027), .A1(n28679), .B0(n11614), .B1(n15025), .Y(
        n11615) );
  AOI21XL U22630 ( .A0(n15023), .A1(n11999), .B0(n11874), .Y(n11614) );
  OAI21XL U22631 ( .A0(n11999), .A1(n11911), .B0(n11910), .Y(n11912) );
  AOI22XL U22632 ( .A0(Q2_addr[7]), .A1(n5904), .B0(Q3_addr[7]), .B1(n27281), 
        .Y(n11921) );
  AOI22XL U22633 ( .A0(Q2_addr[6]), .A1(n5904), .B0(Q3_addr[6]), .B1(n27281), 
        .Y(n11925) );
  AOI22XL U22634 ( .A0(Q2_addr[5]), .A1(n5904), .B0(Q3_addr[5]), .B1(n27281), 
        .Y(n11923) );
  AOI21XL U22635 ( .A0(n5921), .A1(Q0_addr[4]), .B0(n27078), .Y(n27080) );
  AOI22XL U22636 ( .A0(Q3_addr[4]), .A1(n27281), .B0(Q2_addr[4]), .B1(n5904), 
        .Y(n27079) );
  AOI22XL U22637 ( .A0(Q3_addr[3]), .A1(n27281), .B0(Q2_addr[3]), .B1(n5904), 
        .Y(n11927) );
  AOI22XL U22638 ( .A0(Q3_addr[2]), .A1(n27281), .B0(Q2_addr[2]), .B1(n5904), 
        .Y(n27076) );
  AOI22XL U22639 ( .A0(Q3_addr[1]), .A1(n27281), .B0(Q2_addr[1]), .B1(n5904), 
        .Y(n27074) );
  AOI22XL U22640 ( .A0(Q3_addr[0]), .A1(n27281), .B0(Q2_addr[0]), .B1(n5904), 
        .Y(n27071) );
  NOR2XL U22641 ( .A(n11989), .B(n11990), .Y(A1_WEN) );
  AOI211XL U22642 ( .A0(n28252), .A1(n28350), .B0(n28349), .C0(n28191), .Y(
        n28192) );
  OAI22XL U22643 ( .A0(n28237), .A1(n28347), .B0(n28346), .B1(n28179), .Y(
        n28191) );
  AOI211XL U22644 ( .A0(n28252), .A1(n28343), .B0(n28342), .C0(n28189), .Y(
        n28190) );
  OAI22XL U22645 ( .A0(n28237), .A1(n28340), .B0(n28345), .B1(n5825), .Y(
        n28189) );
  AOI211XL U22646 ( .A0(n28252), .A1(n28336), .B0(n28335), .C0(n28187), .Y(
        n28188) );
  OAI22XL U22647 ( .A0(n28186), .A1(n28333), .B0(n28338), .B1(n28179), .Y(
        n28187) );
  AOI211XL U22648 ( .A0(n28252), .A1(n28329), .B0(n28328), .C0(n28184), .Y(
        n28185) );
  OAI22XL U22649 ( .A0(n28237), .A1(n28326), .B0(n28331), .B1(n5825), .Y(
        n28184) );
  OAI22XL U22650 ( .A0(n28237), .A1(n28318), .B0(n28324), .B1(n5825), .Y(
        n28182) );
  AOI211XL U22651 ( .A0(n11929), .A1(n28626), .B0(n28625), .C0(n28279), .Y(
        n28280) );
  OAI22XL U22652 ( .A0(n28237), .A1(n28623), .B0(n28628), .B1(n5825), .Y(
        n28279) );
  AOI211XL U22653 ( .A0(n28252), .A1(n28619), .B0(n28625), .C0(n28276), .Y(
        n28277) );
  OAI22XL U22654 ( .A0(n28237), .A1(n28617), .B0(n28621), .B1(n27431), .Y(
        n28276) );
  OAI22XL U22655 ( .A0(n28186), .A1(n28311), .B0(n28310), .B1(n27431), .Y(
        n28180) );
  AOI211XL U22656 ( .A0(n28252), .A1(n28613), .B0(n28625), .C0(n28274), .Y(
        n28275) );
  OAI22XL U22657 ( .A0(n28237), .A1(n28611), .B0(n28610), .B1(n5916), .Y(
        n28274) );
  AOI211XL U22658 ( .A0(n28252), .A1(n28607), .B0(n28625), .C0(n28272), .Y(
        n28273) );
  OAI22XL U22659 ( .A0(n28237), .A1(n28605), .B0(n28604), .B1(n5916), .Y(
        n28272) );
  AOI211XL U22660 ( .A0(n28252), .A1(n28601), .B0(n28625), .C0(n28269), .Y(
        n28270) );
  OAI22XL U22661 ( .A0(n28237), .A1(n28599), .B0(n28603), .B1(n27431), .Y(
        n28269) );
  AOI211XL U22662 ( .A0(n28252), .A1(n28595), .B0(n28625), .C0(n28267), .Y(
        n28268) );
  OAI22XL U22663 ( .A0(n28237), .A1(n28593), .B0(n28597), .B1(n28179), .Y(
        n28267) );
  AOI211XL U22664 ( .A0(n28252), .A1(n28589), .B0(n28625), .C0(n28265), .Y(
        n28266) );
  OAI22XL U22665 ( .A0(n28237), .A1(n28587), .B0(n28586), .B1(n28179), .Y(
        n28265) );
  AOI211XL U22666 ( .A0(n28252), .A1(n28583), .B0(n28625), .C0(n28263), .Y(
        n28264) );
  OAI22XL U22667 ( .A0(n28237), .A1(n28581), .B0(n28580), .B1(n28179), .Y(
        n28263) );
  AOI211XL U22668 ( .A0(n28252), .A1(n28576), .B0(n28625), .C0(n28261), .Y(
        n28262) );
  OAI22XL U22669 ( .A0(n28237), .A1(n28574), .B0(n28573), .B1(n5916), .Y(
        n28261) );
  AOI211XL U22670 ( .A0(n28252), .A1(n28570), .B0(n28625), .C0(n28259), .Y(
        n28260) );
  OAI22XL U22671 ( .A0(n28237), .A1(n28568), .B0(n28572), .B1(n28179), .Y(
        n28259) );
  AOI211XL U22672 ( .A0(n28252), .A1(n28564), .B0(n28625), .C0(n28257), .Y(
        n28258) );
  OAI22XL U22673 ( .A0(n28237), .A1(n28562), .B0(n28561), .B1(n5916), .Y(
        n28257) );
  AOI211XL U22674 ( .A0(n28252), .A1(n28558), .B0(n28557), .C0(n28255), .Y(
        n28256) );
  OAI22XL U22675 ( .A0(n28237), .A1(n28555), .B0(n28560), .B1(n28179), .Y(
        n28255) );
  AOI211XL U22676 ( .A0(n28252), .A1(n28307), .B0(n28306), .C0(n28177), .Y(
        n28178) );
  OAI22XL U22677 ( .A0(n28237), .A1(n28304), .B0(n28309), .B1(n5825), .Y(
        n28177) );
  AOI211XL U22678 ( .A0(n28252), .A1(n28551), .B0(n28550), .C0(n28253), .Y(
        n28254) );
  OAI22XL U22679 ( .A0(n28237), .A1(n28548), .B0(n28553), .B1(n28179), .Y(
        n28253) );
  AOI211XL U22680 ( .A0(n28252), .A1(n28544), .B0(n28543), .C0(n28250), .Y(
        n28251) );
  OAI22XL U22681 ( .A0(n28237), .A1(n28541), .B0(n28546), .B1(n5916), .Y(
        n28250) );
  AOI211XL U22682 ( .A0(n28252), .A1(n28537), .B0(n28536), .C0(n28248), .Y(
        n28249) );
  OAI22XL U22683 ( .A0(n28237), .A1(n28534), .B0(n28533), .B1(n28179), .Y(
        n28248) );
  AOI211XL U22684 ( .A0(n28252), .A1(n28530), .B0(n28529), .C0(n28246), .Y(
        n28247) );
  OAI22XL U22685 ( .A0(n28237), .A1(n28527), .B0(n28532), .B1(n5916), .Y(
        n28246) );
  OAI22XL U22686 ( .A0(n28186), .A1(n28520), .B0(n28519), .B1(n28179), .Y(
        n28244) );
  AOI211XL U22687 ( .A0(n28252), .A1(n28516), .B0(n28515), .C0(n28242), .Y(
        n28243) );
  OAI22XL U22688 ( .A0(n28186), .A1(n28513), .B0(n28518), .B1(n28179), .Y(
        n28242) );
  OAI22XL U22689 ( .A0(n28186), .A1(n28506), .B0(n28511), .B1(n5916), .Y(
        n28240) );
  OAI22XL U22690 ( .A0(n28186), .A1(n28499), .B0(n28504), .B1(n5916), .Y(
        n28238) );
  AOI211XL U22691 ( .A0(n28252), .A1(n28495), .B0(n28494), .C0(n28235), .Y(
        n28236) );
  OAI22XL U22692 ( .A0(n28237), .A1(n28492), .B0(n28497), .B1(n5916), .Y(
        n28235) );
  AOI211XL U22693 ( .A0(n28252), .A1(n28488), .B0(n28487), .C0(n28233), .Y(
        n28234) );
  OAI22XL U22694 ( .A0(n28237), .A1(n28485), .B0(n28484), .B1(n28179), .Y(
        n28233) );
  OAI22XL U22695 ( .A0(n28186), .A1(n28297), .B0(n28296), .B1(n28179), .Y(
        n28175) );
  AOI211XL U22696 ( .A0(n28252), .A1(n28481), .B0(n28480), .C0(n28231), .Y(
        n28232) );
  OAI22XL U22697 ( .A0(n28237), .A1(n28478), .B0(n28477), .B1(n28179), .Y(
        n28231) );
  AOI211XL U22698 ( .A0(n28252), .A1(n28474), .B0(n28473), .C0(n28229), .Y(
        n28230) );
  OAI22XL U22699 ( .A0(n28237), .A1(n28471), .B0(n28470), .B1(n28179), .Y(
        n28229) );
  OAI22XL U22700 ( .A0(n28237), .A1(n28464), .B0(n28469), .B1(n5916), .Y(
        n28227) );
  OAI22XL U22701 ( .A0(n28237), .A1(n28457), .B0(n28456), .B1(n28179), .Y(
        n28225) );
  AOI211XL U22702 ( .A0(n28252), .A1(n28453), .B0(n28452), .C0(n28223), .Y(
        n28224) );
  OAI22XL U22703 ( .A0(n28237), .A1(n28450), .B0(n28449), .B1(n28179), .Y(
        n28223) );
  AOI211XL U22704 ( .A0(n28252), .A1(n28446), .B0(n28452), .C0(n28221), .Y(
        n28222) );
  OAI22XL U22705 ( .A0(n28237), .A1(n28444), .B0(n28448), .B1(n28179), .Y(
        n28221) );
  AOI211XL U22706 ( .A0(n28252), .A1(n28440), .B0(n28452), .C0(n28219), .Y(
        n28220) );
  OAI22XL U22707 ( .A0(n28237), .A1(n28438), .B0(n28437), .B1(n5916), .Y(
        n28219) );
  AOI211XL U22708 ( .A0(n28252), .A1(n28434), .B0(n28452), .C0(n28217), .Y(
        n28218) );
  OAI22XL U22709 ( .A0(n28237), .A1(n28432), .B0(n28431), .B1(n5916), .Y(
        n28217) );
  AOI211XL U22710 ( .A0(n28252), .A1(n28428), .B0(n28452), .C0(n28215), .Y(
        n28216) );
  OAI22XL U22711 ( .A0(n28237), .A1(n28426), .B0(n28430), .B1(n5916), .Y(
        n28215) );
  AOI211XL U22712 ( .A0(n28252), .A1(n28422), .B0(n28452), .C0(n28213), .Y(
        n28214) );
  OAI22XL U22713 ( .A0(n28237), .A1(n28420), .B0(n28424), .B1(n5825), .Y(
        n28213) );
  OAI22XL U22714 ( .A0(n28186), .A1(n28289), .B0(n28294), .B1(n28179), .Y(
        n28173) );
  AOI211XL U22715 ( .A0(n28252), .A1(n28416), .B0(n28452), .C0(n28211), .Y(
        n28212) );
  OAI22XL U22716 ( .A0(n28237), .A1(n28414), .B0(n28413), .B1(n28179), .Y(
        n28211) );
  AOI211XL U22717 ( .A0(n28252), .A1(n28410), .B0(n28452), .C0(n28209), .Y(
        n28210) );
  OAI22XL U22718 ( .A0(n28237), .A1(n28408), .B0(n28407), .B1(n5825), .Y(
        n28209) );
  AOI211XL U22719 ( .A0(n28252), .A1(n28404), .B0(n28452), .C0(n28207), .Y(
        n28208) );
  OAI22XL U22720 ( .A0(n28237), .A1(n28402), .B0(n28401), .B1(n5916), .Y(
        n28207) );
  AOI211XL U22721 ( .A0(n28252), .A1(n28398), .B0(n28452), .C0(n28205), .Y(
        n28206) );
  OAI22XL U22722 ( .A0(n28237), .A1(n28396), .B0(n28400), .B1(n28179), .Y(
        n28205) );
  AOI211XL U22723 ( .A0(n28252), .A1(n28392), .B0(n28452), .C0(n28203), .Y(
        n28204) );
  OAI22XL U22724 ( .A0(n28237), .A1(n28390), .B0(n28389), .B1(n27431), .Y(
        n28203) );
  OAI22XL U22725 ( .A0(n28237), .A1(n28383), .B0(n28382), .B1(n27431), .Y(
        n28201) );
  OAI22XL U22726 ( .A0(n28237), .A1(n28376), .B0(n28381), .B1(n5916), .Y(
        n28199) );
  OAI22XL U22727 ( .A0(n28237), .A1(n28369), .B0(n28368), .B1(n27431), .Y(
        n28197) );
  AOI211XL U22728 ( .A0(n28252), .A1(n28365), .B0(n28364), .C0(n28195), .Y(
        n28196) );
  OAI22XL U22729 ( .A0(n28237), .A1(n28362), .B0(n28367), .B1(n5916), .Y(
        n28195) );
  AOI211XL U22730 ( .A0(n28252), .A1(n28358), .B0(n28357), .C0(n28193), .Y(
        n28194) );
  OAI22XL U22731 ( .A0(n28237), .A1(n28355), .B0(n28360), .B1(n5916), .Y(
        n28193) );
  AOI211XL U22732 ( .A0(n11929), .A1(n28285), .B0(n7120), .C0(n28171), .Y(
        n28172) );
  OAI22XL U22733 ( .A0(n28237), .A1(n28282), .B0(n28281), .B1(n5825), .Y(
        n28171) );
  INVXL U22734 ( .A(n11897), .Y(n11898) );
  INVXL U22735 ( .A(n28657), .Y(n11899) );
  AOI22XL U22736 ( .A0(n15027), .A1(n28674), .B0(n11626), .B1(n15025), .Y(
        n11627) );
  AOI22XL U22737 ( .A0(Q2_addr[7]), .A1(n27390), .B0(Q3_addr[7]), .B1(n27389), 
        .Y(n11916) );
  AOI22XL U22738 ( .A0(Q2_addr[6]), .A1(n27390), .B0(Q3_addr[6]), .B1(n27389), 
        .Y(n11918) );
  AOI22XL U22739 ( .A0(Q2_addr[5]), .A1(n27390), .B0(Q3_addr[5]), .B1(n27389), 
        .Y(n11901) );
  AOI22XL U22740 ( .A0(Q3_addr[4]), .A1(n27389), .B0(Q2_addr[4]), .B1(n27390), 
        .Y(n11905) );
  AOI22XL U22741 ( .A0(Q3_addr[3]), .A1(n27389), .B0(Q2_addr[3]), .B1(n27390), 
        .Y(n11903) );
  AOI22XL U22742 ( .A0(Q3_addr[2]), .A1(n27389), .B0(Q2_addr[2]), .B1(n27390), 
        .Y(n11914) );
  AOI22XL U22743 ( .A0(Q3_addr[1]), .A1(n27389), .B0(Q2_addr[1]), .B1(n27390), 
        .Y(n11892) );
  AOI22XL U22744 ( .A0(Q3_addr[0]), .A1(n27389), .B0(Q2_addr[0]), .B1(n27390), 
        .Y(n11894) );
  NOR2XL U22745 ( .A(n11989), .B(n11983), .Y(A0_WEN) );
  OAI22XL U22746 ( .A0(n28579), .A1(n28347), .B0(n28346), .B1(n28353), .Y(
        n28348) );
  OAI22XL U22747 ( .A0(n28579), .A1(n28340), .B0(n28339), .B1(n28353), .Y(
        n28341) );
  AOI211XL U22748 ( .A0(n27631), .A1(n28336), .B0(n28335), .C0(n28334), .Y(
        n28337) );
  OAI22XL U22749 ( .A0(n28579), .A1(n28333), .B0(n28332), .B1(n28295), .Y(
        n28334) );
  OAI22XL U22750 ( .A0(n28579), .A1(n28326), .B0(n28325), .B1(n28353), .Y(
        n28327) );
  OAI22XL U22751 ( .A0(n28579), .A1(n28318), .B0(n28317), .B1(n28353), .Y(
        n28319) );
  AOI211XL U22752 ( .A0(n5918), .A1(n28626), .B0(n28625), .C0(n28624), .Y(
        n28627) );
  OAI22XL U22753 ( .A0(n28579), .A1(n28623), .B0(n28622), .B1(n28353), .Y(
        n28624) );
  AOI211XL U22754 ( .A0(n5827), .A1(n28619), .B0(n28625), .C0(n28618), .Y(
        n28620) );
  OAI22XL U22755 ( .A0(n28579), .A1(n28617), .B0(n28616), .B1(n28295), .Y(
        n28618) );
  OAI22XL U22756 ( .A0(n28579), .A1(n28311), .B0(n28310), .B1(n28353), .Y(
        n28312) );
  AOI211XL U22757 ( .A0(n5798), .A1(n28613), .B0(n28625), .C0(n28612), .Y(
        n28614) );
  OAI22XL U22758 ( .A0(n28579), .A1(n28611), .B0(n28610), .B1(n28295), .Y(
        n28612) );
  AOI211XL U22759 ( .A0(n5798), .A1(n28607), .B0(n28625), .C0(n28606), .Y(
        n28608) );
  OAI22XL U22760 ( .A0(n28579), .A1(n28605), .B0(n28604), .B1(n28295), .Y(
        n28606) );
  AOI211XL U22761 ( .A0(n5798), .A1(n28601), .B0(n28625), .C0(n28600), .Y(
        n28602) );
  OAI22XL U22762 ( .A0(n28579), .A1(n28599), .B0(n28598), .B1(n28295), .Y(
        n28600) );
  AOI211XL U22763 ( .A0(n5827), .A1(n28595), .B0(n28625), .C0(n28594), .Y(
        n28596) );
  OAI22XL U22764 ( .A0(n28579), .A1(n28593), .B0(n28592), .B1(n28295), .Y(
        n28594) );
  AOI211XL U22765 ( .A0(n5827), .A1(n28589), .B0(n28625), .C0(n28588), .Y(
        n28590) );
  OAI22XL U22766 ( .A0(n27560), .A1(n28587), .B0(n28586), .B1(n28353), .Y(
        n28588) );
  AOI211XL U22767 ( .A0(n5918), .A1(n28583), .B0(n28625), .C0(n28582), .Y(
        n28584) );
  OAI22XL U22768 ( .A0(n28579), .A1(n28581), .B0(n28580), .B1(n28353), .Y(
        n28582) );
  AOI211XL U22769 ( .A0(n5827), .A1(n28576), .B0(n28625), .C0(n28575), .Y(
        n28577) );
  OAI22XL U22770 ( .A0(n28579), .A1(n28574), .B0(n28573), .B1(n28295), .Y(
        n28575) );
  AOI211XL U22771 ( .A0(n27631), .A1(n28570), .B0(n28625), .C0(n28569), .Y(
        n28571) );
  OAI22XL U22772 ( .A0(n28579), .A1(n28568), .B0(n28567), .B1(n28295), .Y(
        n28569) );
  AOI211XL U22773 ( .A0(n27631), .A1(n28564), .B0(n28625), .C0(n28563), .Y(
        n28565) );
  OAI22XL U22774 ( .A0(n28579), .A1(n28562), .B0(n28561), .B1(n28295), .Y(
        n28563) );
  OAI22XL U22775 ( .A0(n28579), .A1(n28555), .B0(n28554), .B1(n28295), .Y(
        n28556) );
  AOI211XL U22776 ( .A0(n5827), .A1(n28307), .B0(n28306), .C0(n28305), .Y(
        n28308) );
  OAI22XL U22777 ( .A0(n28579), .A1(n28304), .B0(n28303), .B1(n28353), .Y(
        n28305) );
  AOI211XL U22778 ( .A0(n27631), .A1(n28551), .B0(n28550), .C0(n28549), .Y(
        n28552) );
  OAI22XL U22779 ( .A0(n28579), .A1(n28548), .B0(n28547), .B1(n28295), .Y(
        n28549) );
  OAI22XL U22780 ( .A0(n28579), .A1(n28541), .B0(n28540), .B1(n28353), .Y(
        n28542) );
  OAI22XL U22781 ( .A0(n28579), .A1(n28534), .B0(n28533), .B1(n28353), .Y(
        n28535) );
  AOI211XL U22782 ( .A0(n5798), .A1(n28530), .B0(n28529), .C0(n28528), .Y(
        n28531) );
  OAI22XL U22783 ( .A0(n28579), .A1(n28527), .B0(n28526), .B1(n28353), .Y(
        n28528) );
  OAI22XL U22784 ( .A0(n28579), .A1(n28520), .B0(n28519), .B1(n28353), .Y(
        n28521) );
  AOI211XL U22785 ( .A0(n27631), .A1(n28516), .B0(n28515), .C0(n28514), .Y(
        n28517) );
  OAI22XL U22786 ( .A0(n28579), .A1(n28513), .B0(n28512), .B1(n28295), .Y(
        n28514) );
  OAI22XL U22787 ( .A0(n28579), .A1(n28506), .B0(n28505), .B1(n28353), .Y(
        n28507) );
  OAI22XL U22788 ( .A0(n28579), .A1(n28499), .B0(n28498), .B1(n28353), .Y(
        n28500) );
  AOI211XL U22789 ( .A0(n5918), .A1(n28495), .B0(n28494), .C0(n28493), .Y(
        n28496) );
  OAI22XL U22790 ( .A0(n28579), .A1(n28492), .B0(n28491), .B1(n28353), .Y(
        n28493) );
  OAI22XL U22791 ( .A0(n28579), .A1(n28485), .B0(n28484), .B1(n28353), .Y(
        n28486) );
  OAI22XL U22792 ( .A0(n28579), .A1(n28297), .B0(n28296), .B1(n28353), .Y(
        n28298) );
  OAI22XL U22793 ( .A0(n28579), .A1(n28478), .B0(n28477), .B1(n28353), .Y(
        n28479) );
  AOI211XL U22794 ( .A0(n5827), .A1(n28474), .B0(n28473), .C0(n28472), .Y(
        n28475) );
  OAI22XL U22795 ( .A0(n28579), .A1(n28471), .B0(n28470), .B1(n28353), .Y(
        n28472) );
  OAI22XL U22796 ( .A0(n28579), .A1(n28464), .B0(n28463), .B1(n28353), .Y(
        n28465) );
  OAI22XL U22797 ( .A0(n28579), .A1(n28457), .B0(n28456), .B1(n28353), .Y(
        n28458) );
  AOI211XL U22798 ( .A0(n27631), .A1(n28453), .B0(n28452), .C0(n28451), .Y(
        n28454) );
  OAI22XL U22799 ( .A0(n28579), .A1(n28450), .B0(n28449), .B1(n28353), .Y(
        n28451) );
  AOI211XL U22800 ( .A0(n27631), .A1(n28446), .B0(n28452), .C0(n28445), .Y(
        n28447) );
  OAI22XL U22801 ( .A0(n28579), .A1(n28444), .B0(n28443), .B1(n28295), .Y(
        n28445) );
  AOI211XL U22802 ( .A0(n27631), .A1(n28440), .B0(n28452), .C0(n28439), .Y(
        n28441) );
  OAI22XL U22803 ( .A0(n28579), .A1(n28438), .B0(n28437), .B1(n28295), .Y(
        n28439) );
  AOI211XL U22804 ( .A0(n5827), .A1(n28434), .B0(n28452), .C0(n28433), .Y(
        n28435) );
  OAI22XL U22805 ( .A0(n28579), .A1(n28432), .B0(n28431), .B1(n28295), .Y(
        n28433) );
  AOI211XL U22806 ( .A0(n27631), .A1(n28428), .B0(n28452), .C0(n28427), .Y(
        n28429) );
  OAI22XL U22807 ( .A0(n28579), .A1(n28426), .B0(n28425), .B1(n28353), .Y(
        n28427) );
  AOI211XL U22808 ( .A0(n27631), .A1(n28422), .B0(n28452), .C0(n28421), .Y(
        n28423) );
  OAI22XL U22809 ( .A0(n28579), .A1(n28420), .B0(n28419), .B1(n28353), .Y(
        n28421) );
  OAI22XL U22810 ( .A0(n28579), .A1(n28289), .B0(n28288), .B1(n28295), .Y(
        n28290) );
  AOI211XL U22811 ( .A0(n5918), .A1(n28416), .B0(n28452), .C0(n28415), .Y(
        n28417) );
  OAI22XL U22812 ( .A0(n28579), .A1(n28414), .B0(n28413), .B1(n28353), .Y(
        n28415) );
  AOI211XL U22813 ( .A0(n27631), .A1(n28410), .B0(n28452), .C0(n28409), .Y(
        n28411) );
  OAI22XL U22814 ( .A0(n28579), .A1(n28408), .B0(n28407), .B1(n28295), .Y(
        n28409) );
  AOI211XL U22815 ( .A0(n27631), .A1(n28404), .B0(n28452), .C0(n28403), .Y(
        n28405) );
  OAI22XL U22816 ( .A0(n28579), .A1(n28402), .B0(n28401), .B1(n28295), .Y(
        n28403) );
  AOI211XL U22817 ( .A0(n5827), .A1(n28398), .B0(n28452), .C0(n28397), .Y(
        n28399) );
  OAI22XL U22818 ( .A0(n28579), .A1(n28396), .B0(n28395), .B1(n28295), .Y(
        n28397) );
  AOI211XL U22819 ( .A0(n5827), .A1(n28392), .B0(n28452), .C0(n28391), .Y(
        n28393) );
  OAI22XL U22820 ( .A0(n28579), .A1(n28390), .B0(n28389), .B1(n28353), .Y(
        n28391) );
  OAI22XL U22821 ( .A0(n28579), .A1(n28383), .B0(n28382), .B1(n28353), .Y(
        n28384) );
  OAI22XL U22822 ( .A0(n28579), .A1(n28376), .B0(n28375), .B1(n28353), .Y(
        n28377) );
  OAI22XL U22823 ( .A0(n28579), .A1(n28369), .B0(n28368), .B1(n28353), .Y(
        n28370) );
  OAI22XL U22824 ( .A0(n28579), .A1(n28362), .B0(n28361), .B1(n28353), .Y(
        n28363) );
  AOI211XL U22825 ( .A0(n27631), .A1(n28358), .B0(n28357), .C0(n28356), .Y(
        n28359) );
  OAI22XL U22826 ( .A0(n28579), .A1(n28355), .B0(n28354), .B1(n28353), .Y(
        n28356) );
  AOI211XL U22827 ( .A0(n27631), .A1(n28285), .B0(n7120), .C0(n28283), .Y(
        n28286) );
  OAI22XL U22828 ( .A0(n28579), .A1(n28282), .B0(n28281), .B1(n28295), .Y(
        n28283) );
  NOR2BXL U22829 ( .AN(n29242), .B(n15027), .Y(n5750) );
  AOI22XL U22830 ( .A0(n15027), .A1(n28709), .B0(n11616), .B1(n15025), .Y(
        n11617) );
  AOI21XL U22831 ( .A0(n28666), .A1(n28665), .B0(n11897), .Y(n11616) );
  NAND2XL U22832 ( .A(n15027), .B(n28674), .Y(n7138) );
  NAND2XL U22833 ( .A(n15026), .B(n15025), .Y(n7139) );
  AOI21XL U22834 ( .A0(n15024), .A1(n15023), .B0(n28642), .Y(n15026) );
  AOI22XL U22835 ( .A0(n15027), .A1(n28680), .B0(n11634), .B1(n15025), .Y(
        n11635) );
  NAND2XL U22836 ( .A(n15027), .B(n28704), .Y(n7136) );
  NAND2XL U22837 ( .A(n8267), .B(n15025), .Y(n7137) );
  AOI22XL U22838 ( .A0(Q2_addr[7]), .A1(n27496), .B0(Q3_addr[7]), .B1(n27497), 
        .Y(n11932) );
  AOI22XL U22839 ( .A0(Q2_addr[6]), .A1(n27496), .B0(Q3_addr[6]), .B1(n27497), 
        .Y(n11934) );
  AOI22XL U22840 ( .A0(Q2_addr[5]), .A1(n27496), .B0(Q3_addr[5]), .B1(n27497), 
        .Y(n11936) );
  AOI22XL U22841 ( .A0(Q3_addr[4]), .A1(n27497), .B0(Q2_addr[4]), .B1(n27496), 
        .Y(n11938) );
  AOI22XL U22842 ( .A0(Q3_addr[3]), .A1(n27497), .B0(Q2_addr[3]), .B1(n27496), 
        .Y(n11941) );
  AOI22XL U22843 ( .A0(Q3_addr[1]), .A1(n27497), .B0(Q2_addr[1]), .B1(n27496), 
        .Y(n11943) );
  XOR2X2 U22844 ( .A(n11533), .B(n11532), .Y(n6889) );
  CLKINVX3 U22845 ( .A(n14976), .Y(n7863) );
  XOR2X4 U22846 ( .A(n11578), .B(n11577), .Y(n6890) );
  AND2X2 U22847 ( .A(n9899), .B(n9898), .Y(n6891) );
  NAND2X1 U22848 ( .A(n5853), .B(n14948), .Y(n6900) );
  AND2X1 U22849 ( .A(n7843), .B(n14956), .Y(n6901) );
  XOR2X4 U22850 ( .A(n7408), .B(n7407), .Y(n6902) );
  AND2X1 U22851 ( .A(n7388), .B(n10777), .Y(n6903) );
  OR2X2 U22852 ( .A(n24662), .B(n22932), .Y(n6904) );
  NAND2X1 U22853 ( .A(n8675), .B(n7081), .Y(n6906) );
  OR2X2 U22854 ( .A(n7543), .B(U1_A_i_d0[18]), .Y(n6907) );
  INVX1 U22855 ( .A(n14776), .Y(n7884) );
  NAND3XL U22856 ( .A(n7795), .B(n14706), .C(n7034), .Y(n14691) );
  AOI21X2 U22857 ( .A0(n7151), .A1(n8273), .B0(n8272), .Y(n10616) );
  AND2X2 U22858 ( .A(U0_U0_y1[24]), .B(U0_U0_y0[24]), .Y(n6911) );
  OR2X2 U22859 ( .A(BOPB[7]), .B(n7045), .Y(n6912) );
  NAND2X1 U22860 ( .A(n8591), .B(n8590), .Y(n6913) );
  AND2X2 U22861 ( .A(n20014), .B(n20013), .Y(n6915) );
  AND2X4 U22862 ( .A(n7138), .B(n7139), .Y(n6928) );
  AND2X4 U22863 ( .A(n7136), .B(n7137), .Y(n6929) );
  OR2X2 U22864 ( .A(n7434), .B(n20003), .Y(n6938) );
  OR2X2 U22865 ( .A(n19993), .B(n14954), .Y(n6941) );
  AND2X1 U22866 ( .A(n14560), .B(n24643), .Y(n6942) );
  XNOR2X2 U22867 ( .A(n13475), .B(n13476), .Y(n22449) );
  XOR2X4 U22868 ( .A(n7766), .B(n7361), .Y(n6945) );
  AND2X1 U22869 ( .A(n9435), .B(n9434), .Y(n6946) );
  OR2X2 U22870 ( .A(n19259), .B(n20015), .Y(n6947) );
  XOR2X1 U22871 ( .A(n13498), .B(n13497), .Y(n22454) );
  XOR2X1 U22872 ( .A(n14407), .B(n14406), .Y(n25193) );
  OR2X2 U22873 ( .A(n25162), .B(U2_A_r_d[20]), .Y(n6948) );
  XOR2X1 U22874 ( .A(n9546), .B(n9545), .Y(n13717) );
  XNOR2X1 U22875 ( .A(n5875), .B(n12147), .Y(n14530) );
  OR2X2 U22876 ( .A(n20023), .B(n20029), .Y(n6949) );
  INVX1 U22877 ( .A(n14956), .Y(n19999) );
  OR2X2 U22878 ( .A(n25162), .B(U2_A_i_d[20]), .Y(n6951) );
  OR2X2 U22879 ( .A(n9681), .B(U1_A_r_d0[12]), .Y(n6953) );
  AND2X1 U22880 ( .A(n11106), .B(n11105), .Y(n6955) );
  AND2X1 U22881 ( .A(n10626), .B(n10625), .Y(n6959) );
  AND2X1 U22882 ( .A(n12604), .B(n12603), .Y(n6963) );
  AND2X1 U22883 ( .A(n9117), .B(n9116), .Y(n6969) );
  AND2X1 U22884 ( .A(n13407), .B(n13406), .Y(n6970) );
  AND2X1 U22885 ( .A(n12599), .B(n12621), .Y(n6971) );
  AND2X2 U22886 ( .A(n13071), .B(n13073), .Y(n6972) );
  AND2X1 U22887 ( .A(n11082), .B(n11081), .Y(n6976) );
  AND2X1 U22888 ( .A(n13008), .B(n13042), .Y(n6977) );
  AND2X1 U22889 ( .A(n11286), .B(n11285), .Y(n6979) );
  OR2X2 U22890 ( .A(n25212), .B(U2_A_r_d[12]), .Y(n6980) );
  OR2X2 U22891 ( .A(n7837), .B(n13918), .Y(n6982) );
  NAND2X1 U22892 ( .A(n14819), .B(n14818), .Y(n6983) );
  OR2X2 U22893 ( .A(n5820), .B(n7410), .Y(n6984) );
  OR2X2 U22894 ( .A(n19259), .B(n5857), .Y(n6985) );
  OR2X2 U22895 ( .A(n24043), .B(n24042), .Y(n6986) );
  INVX1 U22896 ( .A(n14713), .Y(n7359) );
  OAI21XL U22897 ( .A0(n12841), .A1(n12754), .B0(n12753), .Y(n12906) );
  OR2X2 U22898 ( .A(n22958), .B(n13167), .Y(n6987) );
  OR2X2 U22899 ( .A(n13125), .B(n7346), .Y(n6988) );
  NOR2X1 U22900 ( .A(n25665), .B(n25302), .Y(n6990) );
  OR2X2 U22901 ( .A(n12378), .B(n24620), .Y(n6992) );
  INVX1 U22902 ( .A(n13446), .Y(n7289) );
  OR2X2 U22903 ( .A(n14053), .B(U2_A_r_d[20]), .Y(n6995) );
  OR2X2 U22904 ( .A(n13692), .B(U1_A_i_d0[14]), .Y(n6996) );
  OR2X2 U22905 ( .A(n22917), .B(n24633), .Y(n6997) );
  NOR2X1 U22906 ( .A(n9694), .B(n7070), .Y(n7688) );
  OR2X2 U22907 ( .A(n13699), .B(U1_A_i_d0[18]), .Y(n7001) );
  NAND2X1 U22908 ( .A(n9301), .B(n9300), .Y(n7681) );
  OR2X2 U22909 ( .A(n9681), .B(U1_A_i_d0[12]), .Y(n7007) );
  INVX1 U22910 ( .A(n19563), .Y(n7906) );
  XNOR2X1 U22911 ( .A(n8542), .B(n8532), .Y(n19732) );
  INVX1 U22912 ( .A(n14804), .Y(n7898) );
  INVX1 U22913 ( .A(n19994), .Y(n7434) );
  INVX1 U22914 ( .A(n9476), .Y(n7699) );
  OR2X2 U22915 ( .A(n13387), .B(n13388), .Y(n7015) );
  INVX1 U22916 ( .A(n22917), .Y(n22926) );
  INVX1 U22917 ( .A(n24675), .Y(n24681) );
  AND2X2 U22918 ( .A(n21568), .B(n5765), .Y(n7023) );
  NAND2X2 U22919 ( .A(n7930), .B(n12890), .Y(n7826) );
  OR2X2 U22920 ( .A(n13692), .B(U1_A_r_d0[14]), .Y(n7024) );
  INVX1 U22921 ( .A(n17454), .Y(n7631) );
  NOR2X1 U22922 ( .A(n19237), .B(n14968), .Y(n17299) );
  INVX1 U22923 ( .A(n9485), .Y(n7748) );
  NOR2X2 U22924 ( .A(n9321), .B(n9320), .Y(n9468) );
  AND3X2 U22925 ( .A(n29105), .B(n6910), .C(n8354), .Y(n7031) );
  OR2X2 U22926 ( .A(n14639), .B(n14638), .Y(n7034) );
  NAND2X1 U22927 ( .A(n21996), .B(n21992), .Y(n22319) );
  NOR2X2 U22928 ( .A(n14252), .B(n14253), .Y(n14429) );
  OR2X2 U22929 ( .A(n14952), .B(n7466), .Y(n7035) );
  AND2X2 U22930 ( .A(n8930), .B(n8936), .Y(n7036) );
  NOR2X1 U22931 ( .A(n9068), .B(n9067), .Y(n9162) );
  NOR2X1 U22932 ( .A(n14856), .B(n19237), .Y(n7038) );
  XNOR2X2 U22933 ( .A(n13991), .B(n6957), .Y(n20028) );
  OR2X2 U22934 ( .A(n14837), .B(n19257), .Y(n7040) );
  NAND2X2 U22935 ( .A(n7358), .B(n7452), .Y(n7795) );
  INVX1 U22936 ( .A(n7278), .Y(n13601) );
  NAND2BX1 U22937 ( .AN(n13574), .B(n7279), .Y(n7278) );
  INVX1 U22938 ( .A(n19745), .Y(n19734) );
  INVX1 U22939 ( .A(n13852), .Y(n7869) );
  OR2X2 U22940 ( .A(n7777), .B(BOPA[40]), .Y(n7043) );
  INVX1 U22941 ( .A(n7894), .Y(n7443) );
  NOR2X1 U22942 ( .A(n13925), .B(n13924), .Y(n13938) );
  NOR2X1 U22943 ( .A(n7872), .B(n5837), .Y(n7489) );
  NAND2X1 U22944 ( .A(n8273), .B(n10627), .Y(n10617) );
  CLKINVX3 U22945 ( .A(n7223), .Y(n10647) );
  NAND2X2 U22946 ( .A(n7045), .B(BOPB[7]), .Y(n7223) );
  NAND2X1 U22947 ( .A(n10979), .B(n8320), .Y(n10966) );
  INVX1 U22948 ( .A(n7880), .Y(n13565) );
  OAI21X2 U22949 ( .A0(n7595), .A1(n14393), .B0(n14247), .Y(n14422) );
  INVX1 U22950 ( .A(n7560), .Y(n26606) );
  NAND2X1 U22951 ( .A(U2_U0_y0[28]), .B(U2_U0_y1[28]), .Y(n7560) );
  OR2X2 U22952 ( .A(n18909), .B(n18908), .Y(n7050) );
  INVX1 U22953 ( .A(n9700), .Y(n13698) );
  NOR2X2 U22954 ( .A(n12940), .B(n12941), .Y(n12974) );
  OR2X2 U22955 ( .A(n7133), .B(n7134), .Y(n7078) );
  INVX4 U22956 ( .A(n28998), .Y(n27040) );
  INVX4 U22957 ( .A(n28998), .Y(n21700) );
  CLKINVX3 U22958 ( .A(U2_B_i[9]), .Y(n9629) );
  OAI21X2 U22959 ( .A0(n8359), .A1(n11427), .B0(n8358), .Y(U2_B_i[9]) );
  XNOR2X2 U22960 ( .A(n9644), .B(n9643), .Y(U2_U0_z0[13]) );
  AND2X2 U22961 ( .A(n29105), .B(n29104), .Y(n7422) );
  INVX1 U22962 ( .A(n13687), .Y(n9680) );
  AOI21X1 U22963 ( .A0(n9924), .A1(n9923), .B0(n9922), .Y(n9925) );
  NOR2X1 U22964 ( .A(n23798), .B(n23797), .Y(n23922) );
  NAND2X1 U22965 ( .A(n13857), .B(n13856), .Y(n13870) );
  XOR2X2 U22966 ( .A(n7858), .B(n14772), .Y(n19976) );
  AOI2BB1X1 U22967 ( .A0N(n14768), .A1N(n14767), .B0(n7859), .Y(n7858) );
  OAI21X1 U22968 ( .A0(n29007), .A1(n14974), .B0(n7676), .Y(n7674) );
  AND2X1 U22969 ( .A(n19272), .B(n14833), .Y(n8003) );
  AOI21X1 U22970 ( .A0(n14090), .A1(n22797), .B0(n14089), .Y(n22784) );
  OAI21XL U22971 ( .A0(n17527), .A1(n9458), .B0(n9457), .Y(n9459) );
  CLKINVX3 U22972 ( .A(n11436), .Y(n11555) );
  ADDHX2 U22973 ( .A(U1_U0_y1[26]), .B(U1_U0_y0[26]), .CO(n9317), .S(n9314) );
  AOI21X1 U22974 ( .A0(n21881), .A1(n21770), .B0(n21769), .Y(n21839) );
  NAND2X1 U22975 ( .A(n19637), .B(n19595), .Y(n7177) );
  NAND2BX1 U22976 ( .AN(n19544), .B(n20005), .Y(n19287) );
  XNOR2X2 U22977 ( .A(n10535), .B(n10534), .Y(U1_U0_z0[25]) );
  NAND2X1 U22978 ( .A(n11580), .B(n11579), .Y(n11581) );
  XOR2X2 U22979 ( .A(n8946), .B(n8945), .Y(n24615) );
  AOI21X1 U22980 ( .A0(n25345), .A1(n25337), .B0(n6942), .Y(n25341) );
  XOR2X2 U22981 ( .A(n7216), .B(n6939), .Y(n14922) );
  NOR2X1 U22982 ( .A(n12885), .B(n19519), .Y(n17708) );
  OAI21X1 U22983 ( .A0(n12773), .A1(n12777), .B0(n12779), .Y(n7216) );
  CMPR22X1 U22984 ( .A(U1_U0_y2[19]), .B(U1_U0_y0[19]), .CO(n8416), .S(n8413)
         );
  XOR2X1 U22985 ( .A(n20339), .B(n7799), .Y(n20340) );
  CMPR22X1 U22986 ( .A(U1_U2_y1[22]), .B(U1_U2_y0[22]), .CO(n12908), .S(n12902) );
  CMPR22X1 U22987 ( .A(U1_U2_y2[22]), .B(U1_U2_y0[22]), .CO(n13854), .S(n13849) );
  NAND2X1 U22988 ( .A(n7949), .B(W1[21]), .Y(n10195) );
  OAI21X1 U22989 ( .A0(n10327), .A1(n10326), .B0(n10325), .Y(n10328) );
  INVX1 U22990 ( .A(n25567), .Y(n25572) );
  AOI21X2 U22991 ( .A0(n25594), .A1(n25486), .B0(n25485), .Y(n25550) );
  AOI21X1 U22992 ( .A0(n19234), .A1(n7904), .B0(n7903), .Y(n7811) );
  INVX1 U22993 ( .A(n19234), .Y(n19254) );
  NAND3X1 U22994 ( .A(n19234), .B(n7904), .C(n7254), .Y(n7856) );
  AND2X2 U22995 ( .A(n14789), .B(n14790), .Y(n7847) );
  NOR2X1 U22996 ( .A(n19979), .B(n19321), .Y(n19527) );
  AOI21X2 U22997 ( .A0(n20388), .A1(n14882), .B0(n14881), .Y(n20320) );
  ADDHX2 U22998 ( .A(U0_U0_y2[21]), .B(U0_U0_y0[21]), .CO(n14225), .S(n14222)
         );
  OAI21X1 U22999 ( .A0(n14407), .A1(n14403), .B0(n14404), .Y(n14401) );
  AOI21X4 U23000 ( .A0(n25536), .A1(n25521), .B0(n25520), .Y(n25534) );
  NAND2X1 U23001 ( .A(n9720), .B(U1_A_i_d0[25]), .Y(n9547) );
  NOR2X1 U23002 ( .A(n14212), .B(n14211), .Y(n14331) );
  CMPR22X1 U23003 ( .A(U0_U0_y2[15]), .B(U0_U0_y0[15]), .CO(n14212), .S(n14209) );
  INVXL U23004 ( .A(n27771), .Y(n7085) );
  OAI21X1 U23005 ( .A0(Q5[53]), .A1(OP_done1), .B0(n27278), .Y(n27808) );
  OAI21XL U23006 ( .A0(n17056), .A1(n16789), .B0(n16790), .Y(n17053) );
  INVXL U23007 ( .A(U2_B_r[5]), .Y(n7087) );
  CLKINVX3 U23008 ( .A(n14997), .Y(n16375) );
  INVXL U23009 ( .A(n27618), .Y(n7089) );
  INVXL U23010 ( .A(n27649), .Y(n7091) );
  INVXL U23011 ( .A(n27655), .Y(n7093) );
  CMPR22X1 U23012 ( .A(U1_U0_y2[15]), .B(U1_U0_y0[15]), .CO(n8408), .S(n8405)
         );
  CMPR22X1 U23013 ( .A(U1_U0_y1[39]), .B(U1_U0_y0[39]), .CO(n9347), .S(n9345)
         );
  CMPR22X1 U23014 ( .A(U0_U2_y1[39]), .B(U0_U2_y0[39]), .CO(n12351), .S(n9234)
         );
  CMPR22X1 U23015 ( .A(U0_U1_y2[39]), .B(U0_U1_y0[39]), .CO(n13189), .S(n13182) );
  CMPR22X1 U23016 ( .A(U1_U1_y2[39]), .B(U1_U1_y0[39]), .CO(n13655), .S(n13640) );
  CMPR22X1 U23017 ( .A(U1_U2_y1[39]), .B(U1_U2_y0[39]), .CO(n13661), .S(n13647) );
  CMPR22X1 U23018 ( .A(U0_U0_y2[39]), .B(U0_U0_y0[39]), .CO(n14272), .S(n14270) );
  CMPR22X1 U23019 ( .A(U0_U0_y1[36]), .B(U0_U0_y0[36]), .CO(n13290), .S(n13286) );
  INVXL U23020 ( .A(n27570), .Y(n7097) );
  INVXL U23021 ( .A(n27594), .Y(n7099) );
  INVXL U23022 ( .A(n27612), .Y(n7101) );
  INVXL U23023 ( .A(n27734), .Y(n7103) );
  INVXL U23024 ( .A(n27576), .Y(n7105) );
  INVXL U23025 ( .A(n27624), .Y(n7107) );
  INVXL U23026 ( .A(n27770), .Y(n7109) );
  INVXL U23027 ( .A(n27588), .Y(n7111) );
  INVXL U23028 ( .A(n27606), .Y(n7113) );
  OAI21X1 U23029 ( .A0(Q6[23]), .A1(OP_done1), .B0(n27172), .Y(n27638) );
  INVXL U23030 ( .A(n27740), .Y(n7115) );
  OAI21X1 U23031 ( .A0(Q6[50]), .A1(OP_done1), .B0(n27266), .Y(n27790) );
  CMPR22X1 U23032 ( .A(U2_U0_y1[15]), .B(U2_U0_y0[15]), .CO(n25887), .S(n25848) );
  OAI2BB2X2 U23033 ( .B0(n11876), .B1(n15027), .A0N(n15027), .A1N(n28679), .Y(
        n11877) );
  INVXL U23034 ( .A(U2_B_r[22]), .Y(n7117) );
  NAND2X1 U23035 ( .A(n9530), .B(n9529), .Y(n9531) );
  NAND2X1 U23036 ( .A(n11509), .B(n11508), .Y(n11510) );
  NAND2X1 U23037 ( .A(n11570), .B(n11569), .Y(n11571) );
  NAND2X1 U23038 ( .A(n7875), .B(n19565), .Y(n7269) );
  NAND2X1 U23039 ( .A(n12249), .B(n12248), .Y(n12254) );
  CMPR22X1 U23040 ( .A(U1_U2_y1[15]), .B(U1_U2_y0[15]), .CO(n12758), .S(n12755) );
  OAI21XL U23041 ( .A0(n11998), .A1(n11911), .B0(n11910), .Y(n11909) );
  NAND2X2 U23042 ( .A(n7758), .B(n8245), .Y(U2_B_i[11]) );
  AOI21XL U23043 ( .A0(B6_q[33]), .A1(n5926), .B0(n16564), .Y(n15645) );
  AOI21XL U23044 ( .A0(B2_q[1]), .A1(n16570), .B0(n16564), .Y(n16566) );
  AOI21XL U23045 ( .A0(B6_q[0]), .A1(n16570), .B0(n16564), .Y(n15385) );
  AOI21XL U23046 ( .A0(B4_q[34]), .A1(n15687), .B0(n16564), .Y(n15641) );
  AOI21XL U23047 ( .A0(B4_q[36]), .A1(n15687), .B0(n16564), .Y(n15634) );
  AOI21XL U23048 ( .A0(B4_q[30]), .A1(n15687), .B0(n16487), .Y(n15655) );
  AOI21XL U23049 ( .A0(B7_q[31]), .A1(n16325), .B0(n16487), .Y(n15652) );
  AOI21XL U23050 ( .A0(B7_q[32]), .A1(n16325), .B0(n16487), .Y(n15648) );
  AOI21XL U23051 ( .A0(B1_q[20]), .A1(n16559), .B0(n16487), .Y(n16489) );
  AOI21XL U23052 ( .A0(B5_q[49]), .A1(n16165), .B0(n16487), .Y(n15396) );
  NAND2X2 U23053 ( .A(A_sel_reg[0]), .B(n11920), .Y(n15003) );
  NOR2X4 U23054 ( .A(n28677), .B(C_sel_reg[9]), .Y(n15747) );
  XOR2X2 U23055 ( .A(n13646), .B(n7003), .Y(n19237) );
  NOR2X2 U23056 ( .A(n28678), .B(n28671), .Y(n16136) );
  NAND2X2 U23057 ( .A(C_sel_reg[8]), .B(C_sel_reg[9]), .Y(n16348) );
  AOI211XL U23058 ( .A0(n5918), .A1(n28460), .B0(n28459), .C0(n28458), .Y(
        n28461) );
  AOI211XL U23059 ( .A0(n28143), .A1(n28460), .B0(n28459), .C0(n28112), .Y(
        n28113) );
  AOI211XL U23060 ( .A0(n28252), .A1(n28460), .B0(n28459), .C0(n28225), .Y(
        n28226) );
  NOR2BX2 U23061 ( .AN(buffer[18]), .B(n5922), .Y(n28473) );
  NAND2X2 U23062 ( .A(n28678), .B(n28671), .Y(n16154) );
  AOI211XL U23063 ( .A0(n28143), .A1(n28300), .B0(n28299), .C0(n28062), .Y(
        n28063) );
  AOI211XL U23064 ( .A0(n28252), .A1(n28300), .B0(n28299), .C0(n28175), .Y(
        n28176) );
  AOI211XL U23065 ( .A0(n27162), .A1(n28314), .B0(n28313), .C0(n27833), .Y(
        n27834) );
  AOI211XL U23066 ( .A0(n28143), .A1(n28314), .B0(n28313), .C0(n28066), .Y(
        n28067) );
  AOI211XL U23067 ( .A0(n28252), .A1(n28314), .B0(n28313), .C0(n28180), .Y(
        n28181) );
  NOR2BX2 U23068 ( .AN(buffer[7]), .B(n27122), .Y(n28335) );
  NOR2BX2 U23069 ( .AN(buffer[10]), .B(n27122), .Y(n28357) );
  AOI211XL U23070 ( .A0(n5918), .A1(n28379), .B0(n28378), .C0(n28377), .Y(
        n28380) );
  AOI211XL U23071 ( .A0(n28252), .A1(n28379), .B0(n28378), .C0(n28199), .Y(
        n28200) );
  AOI211XL U23072 ( .A0(n28143), .A1(n28379), .B0(n28378), .C0(n28085), .Y(
        n28086) );
  NOR2BX2 U23073 ( .AN(buffer[21]), .B(n5922), .Y(n28494) );
  AOI211XL U23074 ( .A0(n28143), .A1(n28502), .B0(n28501), .C0(n28126), .Y(
        n28127) );
  AOI211XL U23075 ( .A0(n28252), .A1(n28502), .B0(n28501), .C0(n28238), .Y(
        n28239) );
  AOI211X4 U23076 ( .A0(n5918), .A1(n27696), .B0(n28501), .C0(n27695), .Y(
        n27697) );
  AOI211XL U23077 ( .A0(n28143), .A1(n28523), .B0(n28522), .C0(n28132), .Y(
        n28133) );
  AOI211XL U23078 ( .A0(n28252), .A1(n28523), .B0(n28522), .C0(n28244), .Y(
        n28245) );
  NOR2BX2 U23079 ( .AN(buffer[28]), .B(n5922), .Y(n28543) );
  NOR2BX2 U23080 ( .AN(buffer[29]), .B(n5922), .Y(n28550) );
  CLKINVX3 U23081 ( .A(n11953), .Y(n11957) );
  AOI211XL U23082 ( .A0(n27631), .A1(n28292), .B0(n28291), .C0(n28290), .Y(
        n28293) );
  AOI211XL U23083 ( .A0(n28143), .A1(n28292), .B0(n28291), .C0(n28060), .Y(
        n28061) );
  AOI211XL U23084 ( .A0(n28252), .A1(n28292), .B0(n28291), .C0(n28173), .Y(
        n28174) );
  NOR2BX2 U23085 ( .AN(buffer[3]), .B(n27122), .Y(n28306) );
  AOI211XL U23086 ( .A0(n27162), .A1(n28321), .B0(n28320), .C0(n27837), .Y(
        n27838) );
  AOI211XL U23087 ( .A0(n28143), .A1(n28321), .B0(n28320), .C0(n28069), .Y(
        n28070) );
  AOI211XL U23088 ( .A0(n28252), .A1(n28321), .B0(n28320), .C0(n28182), .Y(
        n28183) );
  NOR2BX2 U23089 ( .AN(buffer[6]), .B(n27122), .Y(n28328) );
  NOR2BX2 U23090 ( .AN(buffer[11]), .B(n27122), .Y(n28364) );
  AOI211XL U23091 ( .A0(n28143), .A1(n28372), .B0(n28371), .C0(n28083), .Y(
        n28084) );
  AOI211XL U23092 ( .A0(n5827), .A1(n28372), .B0(n28371), .C0(n28370), .Y(
        n28373) );
  AOI211XL U23093 ( .A0(n28252), .A1(n28372), .B0(n28371), .C0(n28197), .Y(
        n28198) );
  AOI211XL U23094 ( .A0(n28143), .A1(n28386), .B0(n28385), .C0(n28087), .Y(
        n28088) );
  AOI211XL U23095 ( .A0(n5827), .A1(n28386), .B0(n28385), .C0(n28384), .Y(
        n28387) );
  AOI211XL U23096 ( .A0(n28252), .A1(n28386), .B0(n28385), .C0(n28201), .Y(
        n28202) );
  AOI211XL U23097 ( .A0(n28143), .A1(n28467), .B0(n28466), .C0(n28114), .Y(
        n28115) );
  AOI211XL U23098 ( .A0(n5827), .A1(n28467), .B0(n28466), .C0(n28465), .Y(
        n28468) );
  AOI211XL U23099 ( .A0(n28252), .A1(n28467), .B0(n28466), .C0(n28227), .Y(
        n28228) );
  NOR2BX2 U23100 ( .AN(buffer[19]), .B(n5922), .Y(n28480) );
  AOI211XL U23101 ( .A0(n5798), .A1(n28488), .B0(n28487), .C0(n28486), .Y(
        n28489) );
  NOR2BX2 U23102 ( .AN(buffer[20]), .B(n5922), .Y(n28487) );
  AOI211XL U23103 ( .A0(n28252), .A1(n28509), .B0(n28508), .C0(n28240), .Y(
        n28241) );
  AOI211XL U23104 ( .A0(n28143), .A1(n28509), .B0(n28508), .C0(n28128), .Y(
        n28129) );
  AOI211XL U23105 ( .A0(n5826), .A1(n28509), .B0(n28508), .C0(n27965), .Y(
        n27966) );
  NOR2BX2 U23106 ( .AN(buffer[24]), .B(n5922), .Y(n28515) );
  AOI211XL U23107 ( .A0(n5798), .A1(n28537), .B0(n28536), .C0(n28535), .Y(
        n28538) );
  NOR2BX2 U23108 ( .AN(buffer[27]), .B(n5922), .Y(n28536) );
  NOR2BX2 U23109 ( .AN(buffer[30]), .B(n5922), .Y(n28557) );
  MXI2X1 U23110 ( .A(U1_pipe0[27]), .B(n19389), .S0(n19405), .Y(n5130) );
  OAI21XL U23111 ( .A0(n11913), .A1(n28673), .B0(n11909), .Y(B0_addr[3]) );
  INVX12 U23112 ( .A(n7125), .Y(n7126) );
  XNOR2X1 U23113 ( .A(n8013), .B(W0[16]), .Y(U0_U0_z1[0]) );
  CMPR22X1 U23114 ( .A(U0_U1_y1[15]), .B(U0_U1_y0[15]), .CO(n8803), .S(n8800)
         );
  CMPR22X1 U23115 ( .A(U0_U1_y1[16]), .B(U0_U1_y0[16]), .CO(n8805), .S(n8802)
         );
  CMPR22X1 U23116 ( .A(U0_U0_y2[16]), .B(U0_U0_y0[16]), .CO(n14214), .S(n14211) );
  OAI21X1 U23117 ( .A0(n28688), .A1(n11428), .B0(n11407), .Y(U2_B_r[17]) );
  AOI21X1 U23118 ( .A0(n10839), .A1(n10837), .B0(n10831), .Y(n7321) );
  CMPR22X1 U23119 ( .A(U1_U0_y2[16]), .B(U1_U0_y0[16]), .CO(n8410), .S(n8407)
         );
  CMPR22X1 U23120 ( .A(U0_U1_y2[16]), .B(U0_U1_y0[16]), .CO(n12459), .S(n12456) );
  CMPR22X1 U23121 ( .A(U0_U2_y1[35]), .B(U0_U2_y0[35]), .CO(n9192), .S(n9158)
         );
  NOR2X1 U23122 ( .A(n19394), .B(n19085), .Y(n13715) );
  NOR2X1 U23123 ( .A(n22305), .B(n21961), .Y(n13171) );
  NOR2X1 U23124 ( .A(n25538), .B(n25519), .Y(n25521) );
  NOR2X1 U23125 ( .A(n25291), .B(n12401), .Y(n12403) );
  CMPR22X1 U23126 ( .A(U0_U0_y2[14]), .B(U0_U0_y0[14]), .CO(n14210), .S(n14173) );
  CMPR22X1 U23127 ( .A(U0_U0_y2[17]), .B(U0_U0_y0[17]), .CO(n14216), .S(n14213) );
  NOR2X1 U23128 ( .A(n7847), .B(n14788), .Y(n19302) );
  AOI21X2 U23129 ( .A0(n25531), .A1(n5774), .B0(n25525), .Y(n7598) );
  CMPR22X1 U23130 ( .A(U1_U0_y2[39]), .B(U1_U0_y0[39]), .CO(n8459), .S(n8457)
         );
  CMPR22X1 U23131 ( .A(U0_U1_y1[39]), .B(U0_U1_y0[39]), .CO(n12345), .S(n9228)
         );
  CMPR22X1 U23132 ( .A(U1_U1_y1[39]), .B(U1_U1_y0[39]), .CO(n14687), .S(n14685) );
  NOR2X1 U23133 ( .A(n12865), .B(n12866), .Y(n12796) );
  NAND3BX1 U23134 ( .AN(n14716), .B(n14633), .C(n14718), .Y(n7852) );
  CMPR22X1 U23135 ( .A(U1_U2_y2[35]), .B(U1_U2_y0[35]), .CO(n13965), .S(n13956) );
  CMPR22X1 U23136 ( .A(U0_U2_y2[36]), .B(U0_U2_y0[36]), .CO(n12266), .S(n12260) );
  CMPR22X1 U23137 ( .A(U0_U0_y2[36]), .B(U0_U0_y0[36]), .CO(n14265), .S(n14261) );
  OAI21X1 U23138 ( .A0(Q5[45]), .A1(OP_done1), .B0(n27245), .Y(n27764) );
  XOR2X1 U23139 ( .A(n7435), .B(n20342), .Y(n20343) );
  NAND2X2 U23140 ( .A(n9858), .B(n9857), .Y(n10175) );
  NAND2X2 U23141 ( .A(W0[10]), .B(W0[26]), .Y(n9857) );
  NAND2X2 U23142 ( .A(n9894), .B(n9893), .Y(n10307) );
  NAND2X2 U23143 ( .A(n5932), .B(n9840), .Y(n10150) );
  OAI21X1 U23144 ( .A0(Q6[51]), .A1(OP_done1), .B0(n27270), .Y(n27801) );
  NAND2X1 U23145 ( .A(n9899), .B(n9898), .Y(n7129) );
  NAND2X2 U23146 ( .A(n8353), .B(n9811), .Y(n10137) );
  NAND2X2 U23147 ( .A(n9959), .B(n9958), .Y(n10220) );
  CMPR22X1 U23148 ( .A(U2_U0_y1[18]), .B(U2_U0_y0[18]), .CO(n26035), .S(n25986) );
  CMPR22X1 U23149 ( .A(U2_U0_y1[17]), .B(U2_U0_y0[17]), .CO(n25985), .S(n25944) );
  OAI21X1 U23150 ( .A0(n6932), .A1(n11428), .B0(n9614), .Y(U2_B_r[9]) );
  CLKINVX3 U23151 ( .A(n28700), .Y(n11945) );
  NAND2X1 U23152 ( .A(n24710), .B(n24686), .Y(n24703) );
  NOR2X1 U23153 ( .A(n24724), .B(n24683), .Y(n24710) );
  NAND2X1 U23154 ( .A(n19573), .B(n19572), .Y(n19574) );
  NAND2X1 U23155 ( .A(n11485), .B(n11484), .Y(n11486) );
  NAND2X1 U23156 ( .A(n11476), .B(n11475), .Y(n11477) );
  XOR2X2 U23157 ( .A(n11494), .B(n11493), .Y(U2_U0_z0[22]) );
  NAND2X1 U23158 ( .A(n11466), .B(n11463), .Y(n11460) );
  NAND2X1 U23159 ( .A(n14814), .B(n14813), .Y(n14815) );
  XOR2X1 U23160 ( .A(n12962), .B(n12961), .Y(n19311) );
  XOR2X1 U23161 ( .A(n12914), .B(n12913), .Y(n19321) );
  XOR2X1 U23162 ( .A(n14712), .B(n14711), .Y(n19962) );
  NAND2X1 U23163 ( .A(n9424), .B(n9423), .Y(n9425) );
  NAND2X1 U23164 ( .A(n9499), .B(n9498), .Y(n9500) );
  NAND2X1 U23165 ( .A(n13368), .B(n13367), .Y(n13369) );
  NAND2X1 U23166 ( .A(n8958), .B(n8991), .Y(n8959) );
  NAND2X1 U23167 ( .A(n9002), .B(n9015), .Y(n9003) );
  NAND2X1 U23168 ( .A(n5885), .B(n13137), .Y(n12643) );
  NAND2X1 U23169 ( .A(n12227), .B(n12226), .Y(n12228) );
  NAND2X1 U23170 ( .A(n7289), .B(n13447), .Y(n13448) );
  XOR2X2 U23171 ( .A(n7218), .B(n14354), .Y(n25226) );
  NAND2X1 U23172 ( .A(n14427), .B(n14426), .Y(n14428) );
  XOR2X2 U23173 ( .A(n11518), .B(n11517), .Y(U2_U0_z0[18]) );
  XOR2X2 U23174 ( .A(n10829), .B(n10828), .Y(U1_U2_z0[6]) );
  XOR2X1 U23175 ( .A(n7321), .B(n10835), .Y(U1_U2_z0[5]) );
  XNOR2X2 U23176 ( .A(n7498), .B(n13077), .Y(n19553) );
  XNOR2X1 U23177 ( .A(n12956), .B(n12955), .Y(n19532) );
  NAND2X1 U23178 ( .A(n9523), .B(n9522), .Y(n9524) );
  NAND2X1 U23179 ( .A(n9494), .B(n9493), .Y(n9495) );
  NAND2X1 U23180 ( .A(n9441), .B(n9440), .Y(n9442) );
  XNOR2X1 U23181 ( .A(n7221), .B(n8829), .Y(n24610) );
  NAND2X1 U23182 ( .A(n11258), .B(n11257), .Y(n11259) );
  NAND2X1 U23183 ( .A(n11588), .B(n11587), .Y(n11589) );
  NAND2X1 U23184 ( .A(n10401), .B(n10400), .Y(n10402) );
  XNOR2X1 U23185 ( .A(n11180), .B(n11179), .Y(U1_U1_z0[7]) );
  XNOR2X1 U23186 ( .A(n17467), .B(n17466), .Y(n17468) );
  CMPR22X1 U23187 ( .A(U2_U0_y1[36]), .B(U2_U0_y0[36]), .CO(n26990), .S(n26949) );
  CMPR22X1 U23188 ( .A(U2_U0_y2[15]), .B(U2_U0_y0[15]), .CO(n23224), .S(n23177) );
  NOR2X1 U23189 ( .A(n22452), .B(U2_A_r_d[23]), .Y(n24434) );
  XOR2X2 U23190 ( .A(n13481), .B(n13480), .Y(n22452) );
  INVX1 U23191 ( .A(n12946), .Y(n12917) );
  NOR2X2 U23192 ( .A(n12946), .B(n12949), .Y(n12993) );
  CMPR22X1 U23193 ( .A(U2_U0_y1[16]), .B(U2_U0_y0[16]), .CO(n25943), .S(n25888) );
  AOI21X1 U23194 ( .A0(n17462), .A1(n9539), .B0(n9538), .Y(n17456) );
  OAI211X4 U23195 ( .A0(n28755), .A1(n27772), .B0(n27086), .C0(n27085), .Y(
        A0_addr[2]) );
  NAND2X1 U23196 ( .A(n11608), .B(U2_B_r[3]), .Y(n11592) );
  INVX1 U23197 ( .A(n12255), .Y(n7244) );
  NAND2X1 U23198 ( .A(n20012), .B(n20070), .Y(n20058) );
  NOR2X1 U23199 ( .A(n25132), .B(U2_A_r_d[24]), .Y(n25523) );
  CMPR22X1 U23200 ( .A(U1_U1_y2[15]), .B(U1_U1_y0[15]), .CO(n12697), .S(n12694) );
  CMPR22X1 U23201 ( .A(U1_U2_y2[17]), .B(U1_U2_y0[17]), .CO(n13782), .S(n13779) );
  CMPR22X1 U23202 ( .A(U1_U1_y1[36]), .B(U1_U1_y0[36]), .CO(n14680), .S(n14677) );
  OAI21X1 U23203 ( .A0(n28686), .A1(n11428), .B0(n9725), .Y(U2_B_r[19]) );
  NOR2X1 U23204 ( .A(n24677), .B(n13178), .Y(n25292) );
  CMPR22X1 U23205 ( .A(U0_U1_y2[17]), .B(U0_U1_y0[17]), .CO(n12461), .S(n12458) );
  CMPR22X1 U23206 ( .A(U0_U0_y2[19]), .B(U0_U0_y0[19]), .CO(n14221), .S(n14218) );
  AOI21X2 U23207 ( .A0(n25372), .A1(n12384), .B0(n12383), .Y(n25320) );
  CMPR22X1 U23208 ( .A(U1_U2_y1[35]), .B(U1_U2_y0[35]), .CO(n13606), .S(n13574) );
  AOI21X1 U23209 ( .A0(n20420), .A1(n14865), .B0(n14870), .Y(n14871) );
  NAND2X1 U23210 ( .A(n14796), .B(n14795), .Y(n14797) );
  XOR2X2 U23211 ( .A(n13627), .B(n13613), .Y(n14966) );
  NAND2X2 U23212 ( .A(n9965), .B(n9964), .Y(n10227) );
  NOR2X1 U23213 ( .A(n17457), .B(n9541), .Y(n7412) );
  AOI211XL U23214 ( .A0(n28252), .A1(n27793), .B0(n28625), .C0(n27488), .Y(
        n27489) );
  AOI211XL U23215 ( .A0(n28143), .A1(n27793), .B0(n28625), .C0(n27380), .Y(
        n27381) );
  CMPR22X1 U23216 ( .A(U1_U2_y2[15]), .B(U1_U2_y0[15]), .CO(n13778), .S(n13775) );
  CMPR22X1 U23217 ( .A(U0_U2_y1[15]), .B(U0_U2_y0[15]), .CO(n8741), .S(n8738)
         );
  OAI21XL U23218 ( .A0(n12776), .A1(n12786), .B0(n12788), .Y(n12770) );
  CMPR22X1 U23219 ( .A(U1_U0_y1[15]), .B(U1_U0_y0[15]), .CO(n9293), .S(n9290)
         );
  CMPR22X1 U23220 ( .A(U1_U1_y2[16]), .B(U1_U1_y0[16]), .CO(n12699), .S(n12696) );
  NAND2X1 U23221 ( .A(n13247), .B(n13246), .Y(n13355) );
  NOR2X1 U23222 ( .A(n13246), .B(n13247), .Y(n13354) );
  CMPR22X1 U23223 ( .A(U0_U0_y1[15]), .B(U0_U0_y0[15]), .CO(n13247), .S(n13244) );
  NAND2BX1 U23224 ( .AN(n9694), .B(U1_A_i_d0[16]), .Y(n17216) );
  CMPR22X1 U23225 ( .A(U1_U1_y1[35]), .B(U1_U1_y0[35]), .CO(n14678), .S(n14675) );
  CMPR22X1 U23226 ( .A(U1_U0_y1[19]), .B(U1_U0_y0[19]), .CO(n9303), .S(n9300)
         );
  NOR2X1 U23227 ( .A(n13284), .B(n13283), .Y(n13470) );
  CMPR22X1 U23228 ( .A(U0_U0_y1[35]), .B(U0_U0_y0[35]), .CO(n13287), .S(n13283) );
  AOI22X2 U23229 ( .A0(cnt[9]), .A1(n11998), .B0(n11999), .B1(n28758), .Y(
        n11993) );
  CLKINVX3 U23230 ( .A(in_valid), .Y(n11971) );
  OAI21X2 U23231 ( .A0(n29100), .A1(n11428), .B0(n9611), .Y(U2_B_r[7]) );
  INVX12 U23232 ( .A(n11651), .Y(T1_rom_addr[3]) );
  NOR2X2 U23233 ( .A(n11445), .B(U2_B_r[18]), .Y(n11514) );
  BUFX3 U23234 ( .A(T1_rom_addr[6]), .Y(n7131) );
  BUFX3 U23235 ( .A(T1_rom_addr[7]), .Y(n7132) );
  NOR2BX2 U23236 ( .AN(buffer[26]), .B(n5922), .Y(n28529) );
  NOR2BX2 U23237 ( .AN(buffer[8]), .B(n5922), .Y(n28342) );
  NOR2BX2 U23238 ( .AN(buffer[9]), .B(n27122), .Y(n28349) );
  OAI21XL U23239 ( .A0(n12945), .A1(n7820), .B0(n7818), .Y(n7817) );
  OR2X2 U23240 ( .A(n13387), .B(n7609), .Y(n7608) );
  NOR2X4 U23241 ( .A(n11655), .B(n11653), .Y(n11864) );
  NOR2X1 U23242 ( .A(n14897), .B(n29008), .Y(n12338) );
  NOR2X2 U23243 ( .A(C_sel_reg[1]), .B(n27298), .Y(n27496) );
  NAND3X2 U23244 ( .A(n27122), .B(n28707), .C(A_sel_reg[0]), .Y(n27298) );
  OR2X2 U23245 ( .A(n7696), .B(U1_A_i_d0[20]), .Y(n13728) );
  INVX12 U23246 ( .A(n16348), .Y(n16325) );
  OAI21XL U23247 ( .A0(n11913), .A1(n28673), .B0(n11912), .Y(B2_addr[3]) );
  AOI211XL U23248 ( .A0(n5826), .A1(n28416), .B0(n28452), .C0(n27902), .Y(
        n27903) );
  AOI211XL U23249 ( .A0(n5826), .A1(n28422), .B0(n28452), .C0(n27907), .Y(
        n27908) );
  AOI211XL U23250 ( .A0(n5826), .A1(n27653), .B0(n28452), .C0(n27181), .Y(
        n27182) );
  AOI211XL U23251 ( .A0(n5826), .A1(n27647), .B0(n28452), .C0(n27177), .Y(
        n27178) );
  AOI211XL U23252 ( .A0(n5826), .A1(n28300), .B0(n28299), .C0(n27825), .Y(
        n27826) );
  AOI211XL U23253 ( .A0(n5826), .A1(n28502), .B0(n28501), .C0(n27961), .Y(
        n27962) );
  AOI211XL U23254 ( .A0(n5826), .A1(n28495), .B0(n28494), .C0(n27956), .Y(
        n27957) );
  AOI211XL U23255 ( .A0(n5826), .A1(n28523), .B0(n28522), .C0(n27973), .Y(
        n27974) );
  CLKINVX3 U23256 ( .A(n16293), .Y(n15633) );
  NOR2X4 U23257 ( .A(C_sel_reg[8]), .B(n28671), .Y(n16293) );
  INVX12 U23258 ( .A(n15948), .Y(n15958) );
  OAI21XL U23259 ( .A0(n7768), .A1(n11427), .B0(n11426), .Y(U2_B_i[25]) );
  OAI21X2 U23260 ( .A0(n9551), .A1(n11427), .B0(n9550), .Y(U2_B_i[6]) );
  AOI21X1 U23261 ( .A0(n7024), .A1(n19443), .B0(n13693), .Y(n19432) );
  AOI21XL U23262 ( .A0(n20067), .A1(n20059), .B0(n6915), .Y(n20063) );
  AOI21X1 U23263 ( .A0(n20957), .A1(n20956), .B0(n20955), .Y(n21186) );
  NAND2XL U23264 ( .A(n20815), .B(n20814), .Y(n20849) );
  NAND2X2 U23265 ( .A(n21528), .B(n7023), .Y(n7343) );
  NAND3X4 U23266 ( .A(n7657), .B(n7655), .C(n7660), .Y(n7628) );
  OAI21X1 U23267 ( .A0(n10119), .A1(n10130), .B0(n10118), .Y(n10120) );
  CMPR22X1 U23268 ( .A(U1_U0_y1[16]), .B(U1_U0_y0[16]), .CO(n9295), .S(n9292)
         );
  OAI21XL U23269 ( .A0(n7141), .A1(n8053), .B0(n7347), .Y(n4951) );
  XOR2X1 U23270 ( .A(n7676), .B(n7675), .Y(n14975) );
  NAND2X1 U23271 ( .A(n7619), .B(n8617), .Y(n16944) );
  AOI21X1 U23272 ( .A0(n8402), .A1(n8494), .B0(n8401), .Y(n8403) );
  NAND2X1 U23273 ( .A(n13694), .B(U1_A_r_d0[15]), .Y(n19435) );
  NOR2X2 U23274 ( .A(W0[28]), .B(W0[12]), .Y(n9859) );
  OAI21X1 U23275 ( .A0(n10202), .A1(n10218), .B0(n10201), .Y(n10203) );
  NAND2X1 U23276 ( .A(n5774), .B(n25524), .Y(n25530) );
  INVX1 U23277 ( .A(n10212), .Y(n7583) );
  AOI21X1 U23278 ( .A0(n14472), .A1(n14260), .B0(n14263), .Y(n14477) );
  AOI21X1 U23279 ( .A0(n23049), .A1(n23029), .B0(n23028), .Y(n23039) );
  NOR2X1 U23280 ( .A(n12457), .B(n12456), .Y(n12482) );
  NOR2X1 U23281 ( .A(n22908), .B(n24608), .Y(n23093) );
  AOI21X2 U23282 ( .A0(n10121), .A1(n10128), .B0(n10120), .Y(n10185) );
  INVX1 U23283 ( .A(n9864), .Y(n9815) );
  CLKINVX3 U23284 ( .A(n7627), .Y(n13692) );
  INVX4 U23285 ( .A(n8585), .Y(n7398) );
  BUFX3 U23286 ( .A(n7197), .Y(n7142) );
  OAI21X1 U23287 ( .A0(n11134), .A1(n11142), .B0(n11135), .Y(n11119) );
  NOR2X4 U23288 ( .A(n8123), .B(BOPB[32]), .Y(n10650) );
  NOR2X4 U23289 ( .A(W0[9]), .B(W0[25]), .Y(n9812) );
  CLKINVX3 U23290 ( .A(n7144), .Y(n7205) );
  XNOR2X2 U23291 ( .A(n9819), .B(n10126), .Y(U0_U0_z2[14]) );
  XOR2X2 U23292 ( .A(n7147), .B(n6892), .Y(n22917) );
  OAI21X1 U23293 ( .A0(n12571), .A1(n12581), .B0(n12584), .Y(n7147) );
  AOI2BB1X2 U23294 ( .A0N(n13154), .A1N(n12563), .B0(n12587), .Y(n12571) );
  XOR2X4 U23295 ( .A(n7149), .B(n6924), .Y(U1_U0_z0[22]) );
  AOI21X1 U23296 ( .A0(n10556), .A1(n10548), .B0(n10547), .Y(n7150) );
  OAI21X4 U23297 ( .A0(n10634), .A1(n10640), .B0(n10635), .Y(n7151) );
  AOI21XL U23298 ( .A0(n7151), .A1(n10631), .B0(n10622), .Y(n10623) );
  NAND2XL U23299 ( .A(n7493), .B(n7153), .Y(n7492) );
  NAND2X1 U23300 ( .A(n12064), .B(n12065), .Y(n12095) );
  AOI21X2 U23301 ( .A0(n7156), .A1(n13923), .B0(n7155), .Y(n7154) );
  NOR2X2 U23302 ( .A(n13902), .B(n13903), .Y(n13922) );
  AOI21X1 U23303 ( .A0(n7157), .A1(n7864), .B0(n7436), .Y(n7435) );
  NAND2X2 U23304 ( .A(n8441), .B(n8440), .Y(n8597) );
  NOR2X2 U23305 ( .A(n8444), .B(n8445), .Y(n8589) );
  XOR2XL U23306 ( .A(n19790), .B(n29008), .Y(n7165) );
  XOR2X4 U23307 ( .A(n11389), .B(n11291), .Y(U0_U1_z0[16]) );
  XOR2X4 U23308 ( .A(n11249), .B(n6960), .Y(U0_U1_z0[23]) );
  NAND2X2 U23309 ( .A(n7169), .B(n7168), .Y(n13476) );
  NAND2X2 U23310 ( .A(n13278), .B(n13277), .Y(n13438) );
  NAND2X1 U23311 ( .A(n8196), .B(AOPD[41]), .Y(n10941) );
  NAND2X1 U23312 ( .A(n7170), .B(n10217), .Y(n10211) );
  NAND2X2 U23313 ( .A(n8103), .B(AOPD[27]), .Y(n11033) );
  NOR2X2 U23314 ( .A(n8103), .B(AOPD[27]), .Y(n11032) );
  NAND2X4 U23315 ( .A(n7201), .B(n7447), .Y(n13048) );
  NAND2X1 U23316 ( .A(n12756), .B(n12755), .Y(n12871) );
  NAND2X1 U23317 ( .A(n13570), .B(n13569), .Y(n7176) );
  OAI21X2 U23318 ( .A0(n13073), .A1(n13074), .B0(n13072), .Y(n13569) );
  OAI21XL U23319 ( .A0(n19607), .A1(n19600), .B0(n19604), .Y(n19602) );
  XOR2X1 U23320 ( .A(n8052), .B(n7178), .Y(n17298) );
  XOR2X4 U23321 ( .A(n11478), .B(n11477), .Y(U2_U0_z0[24]) );
  NOR2X1 U23322 ( .A(n8954), .B(n8955), .Y(n8990) );
  NAND2X1 U23323 ( .A(n8951), .B(n7740), .Y(n7181) );
  NAND2X1 U23324 ( .A(n8947), .B(n7740), .Y(n7182) );
  NAND2X1 U23325 ( .A(n13906), .B(n7184), .Y(n13907) );
  OAI21X1 U23326 ( .A0(n9135), .A1(n9131), .B0(n9132), .Y(n7186) );
  AND2X2 U23327 ( .A(n7063), .B(n19724), .Y(n19917) );
  NOR2X4 U23328 ( .A(n10313), .B(n10269), .Y(n7193) );
  OAI21X4 U23329 ( .A0(n7342), .A1(n14991), .B0(n7195), .Y(n10339) );
  BUFX12 U23330 ( .A(n11030), .Y(n7197) );
  XOR2X4 U23331 ( .A(n7198), .B(n6975), .Y(U0_U2_z0[18]) );
  OAI21X2 U23332 ( .A0(n7197), .A1(n10923), .B0(n10922), .Y(n7198) );
  AOI21X4 U23333 ( .A0(n10988), .A1(n8326), .B0(n8325), .Y(n11030) );
  OAI21X4 U23334 ( .A0(n11163), .A1(n11169), .B0(n11164), .Y(n11156) );
  NOR2X2 U23335 ( .A(n8117), .B(BOPC[35]), .Y(n11163) );
  NAND2X2 U23336 ( .A(n12999), .B(n12993), .Y(n13041) );
  NOR2X2 U23337 ( .A(n12992), .B(n12996), .Y(n12999) );
  NOR2X1 U23338 ( .A(W1[29]), .B(W1[13]), .Y(n9948) );
  NAND2X1 U23339 ( .A(n8179), .B(BOPB[41]), .Y(n9554) );
  OAI21X1 U23340 ( .A0(n19277), .A1(n14832), .B0(n14831), .Y(n7203) );
  NAND2X2 U23341 ( .A(n7844), .B(n7848), .Y(n19299) );
  NAND2X2 U23342 ( .A(n11014), .B(n7207), .Y(n7206) );
  NAND2X1 U23343 ( .A(n13584), .B(n13578), .Y(n13588) );
  NOR2X1 U23344 ( .A(n13081), .B(n13078), .Y(n13578) );
  XOR2X2 U23345 ( .A(n7211), .B(n13657), .Y(n14976) );
  OAI21XL U23346 ( .A0(n13654), .A1(n13653), .B0(n13652), .Y(n7211) );
  XOR2X2 U23347 ( .A(n10151), .B(n10152), .Y(U0_U0_z1[5]) );
  OAI21X4 U23348 ( .A0(n9839), .A1(n9842), .B0(n9840), .Y(n9830) );
  NAND2X2 U23349 ( .A(W0[21]), .B(W0[5]), .Y(n9840) );
  NOR2X4 U23350 ( .A(W0[5]), .B(W0[21]), .Y(n9839) );
  XOR2X1 U23351 ( .A(n17632), .B(n17640), .Y(n17642) );
  XNOR2X2 U23352 ( .A(n11607), .B(n11606), .Y(U2_U0_z0[20]) );
  NOR2X4 U23353 ( .A(W1[26]), .B(W1[10]), .Y(n9986) );
  NAND2BX2 U23354 ( .AN(BOPA[41]), .B(n28683), .Y(n7331) );
  AOI21XL U23355 ( .A0(n8661), .A1(n7217), .B0(n8660), .Y(n16703) );
  AOI21X2 U23356 ( .A0(n14369), .A1(n14356), .B0(n14350), .Y(n7218) );
  CLKINVX3 U23357 ( .A(n7934), .Y(n10643) );
  NAND2XL U23358 ( .A(n7934), .B(n7048), .Y(n7935) );
  OAI21X2 U23359 ( .A0(n10651), .A1(n10647), .B0(n6912), .Y(n7567) );
  NOR2X1 U23360 ( .A(n8076), .B(AOPB[30]), .Y(n10490) );
  XOR2X2 U23361 ( .A(n7224), .B(n6983), .Y(n14826) );
  NOR2X2 U23362 ( .A(W3[6]), .B(W3[22]), .Y(n9799) );
  NOR2X2 U23363 ( .A(W3[23]), .B(W3[7]), .Y(n9748) );
  NAND2BX1 U23364 ( .AN(n24666), .B(n24665), .Y(n8035) );
  AND2X2 U23365 ( .A(n14775), .B(n14657), .Y(n7815) );
  NOR2X1 U23366 ( .A(n14779), .B(n14776), .Y(n14657) );
  NOR2X1 U23367 ( .A(n14654), .B(n14655), .Y(n14779) );
  XOR2X1 U23368 ( .A(n24862), .B(n13532), .Y(n13533) );
  NAND2X1 U23369 ( .A(n24662), .B(n7229), .Y(n23016) );
  NAND2X1 U23370 ( .A(n13355), .B(n7610), .Y(n13318) );
  AND2X2 U23371 ( .A(n7606), .B(n7608), .Y(n7232) );
  XOR2X4 U23372 ( .A(n7236), .B(n7235), .Y(U1_U2_z2[15]) );
  XOR2X1 U23373 ( .A(n7978), .B(n8001), .Y(n7235) );
  OAI2BB1X2 U23374 ( .A0N(n9930), .A1N(n9934), .B0(n9929), .Y(n7236) );
  NOR2X2 U23375 ( .A(n14229), .B(n14230), .Y(n14351) );
  AOI21X2 U23376 ( .A0(n7238), .A1(n7704), .B0(n7702), .Y(n7706) );
  OAI21XL U23377 ( .A0(n10820), .A1(n10826), .B0(n10821), .Y(n7239) );
  NAND2X1 U23378 ( .A(n8122), .B(BOPD[33]), .Y(n10821) );
  NOR2X2 U23379 ( .A(n10825), .B(n10820), .Y(n8251) );
  NOR2X2 U23380 ( .A(n8122), .B(BOPD[33]), .Y(n10820) );
  NAND2X1 U23381 ( .A(n8128), .B(BOPD[31]), .Y(n10833) );
  CLKINVX3 U23382 ( .A(n7247), .Y(n7240) );
  NOR2XL U23383 ( .A(n7250), .B(n7240), .Y(n7249) );
  INVX2 U23384 ( .A(n12217), .Y(n7242) );
  NAND2X1 U23385 ( .A(n12224), .B(n7249), .Y(n7248) );
  XOR2X2 U23386 ( .A(n7251), .B(n14274), .Y(n25123) );
  NOR2X1 U23387 ( .A(n14425), .B(n14429), .Y(n14256) );
  NAND2X4 U23388 ( .A(n11636), .B(cs[0]), .Y(n27122) );
  OR2X2 U23389 ( .A(n24666), .B(n22930), .Y(n14117) );
  NOR2X1 U23390 ( .A(n11114), .B(n11123), .Y(n8286) );
  NOR2X1 U23391 ( .A(n8180), .B(BOPC[41]), .Y(n11114) );
  XOR2X2 U23392 ( .A(n10321), .B(n10320), .Y(U1_U2_z1[5]) );
  NOR2BX1 U23393 ( .AN(n9180), .B(n9195), .Y(n7253) );
  INVXL U23394 ( .A(n19233), .Y(n7255) );
  AOI2BB1X2 U23395 ( .A0N(n14839), .A1N(n14841), .B0(n7805), .Y(n7370) );
  NOR2X1 U23396 ( .A(n14675), .B(n14676), .Y(n14841) );
  NAND2X1 U23397 ( .A(n14678), .B(n14677), .Y(n14844) );
  OAI21X2 U23398 ( .A0(n9846), .A1(n9851), .B0(n9847), .Y(n7260) );
  NOR2X2 U23399 ( .A(n9846), .B(n9850), .Y(n7261) );
  NOR2X4 U23400 ( .A(n6876), .B(W0[18]), .Y(n9850) );
  NOR2X4 U23401 ( .A(W0[19]), .B(W0[3]), .Y(n9846) );
  OAI21X4 U23402 ( .A0(n10159), .A1(n12001), .B0(n10160), .Y(n9845) );
  NAND2X2 U23403 ( .A(W0[16]), .B(W0[0]), .Y(n12001) );
  NOR2X4 U23404 ( .A(W0[17]), .B(W0[1]), .Y(n10159) );
  XOR2X4 U23405 ( .A(n11538), .B(n11537), .Y(U2_U0_z0[15]) );
  INVX1 U23406 ( .A(n9824), .Y(n7264) );
  XOR2X4 U23407 ( .A(n7267), .B(n5763), .Y(U0_U0_z2[11]) );
  MXI2X1 U23408 ( .A(n7268), .B(U1_pipe1[26]), .S0(n5928), .Y(n5010) );
  NOR2X4 U23409 ( .A(W0[10]), .B(W0[26]), .Y(n9856) );
  OR2X4 U23410 ( .A(n13603), .B(n7912), .Y(n13573) );
  AOI21X4 U23411 ( .A0(n12999), .A1(n12998), .B0(n12997), .Y(n13047) );
  NAND2X2 U23412 ( .A(n8116), .B(BOPB[35]), .Y(n10635) );
  NOR2X4 U23413 ( .A(n8116), .B(BOPB[35]), .Y(n10634) );
  NOR2X4 U23414 ( .A(n13269), .B(n13270), .Y(n13409) );
  CLKINVX8 U23415 ( .A(n9873), .Y(U0_U0_z2[16]) );
  OAI21X1 U23416 ( .A0(n7273), .A1(n10125), .B0(n10124), .Y(n7578) );
  XOR2X1 U23417 ( .A(n7273), .B(n10167), .Y(U0_U0_z1[12]) );
  NAND2X1 U23418 ( .A(n7274), .B(n14853), .Y(n19240) );
  CLKINVX3 U23419 ( .A(n14146), .Y(n22448) );
  NAND2X1 U23420 ( .A(n12761), .B(n12762), .Y(n12814) );
  INVX2 U23421 ( .A(n7306), .Y(n13469) );
  NAND2BX4 U23422 ( .AN(n13429), .B(n13428), .Y(n7306) );
  AOI21X2 U23423 ( .A0(n13403), .A1(n7571), .B0(n7570), .Y(n7282) );
  NAND2X4 U23424 ( .A(n7571), .B(n13404), .Y(n7283) );
  AOI21X2 U23425 ( .A0(n13048), .A1(n12993), .B0(n12998), .Y(n12962) );
  XOR2X1 U23426 ( .A(n7284), .B(n24990), .Y(n24991) );
  NOR2X1 U23427 ( .A(n8940), .B(n8939), .Y(n8979) );
  NOR2X1 U23428 ( .A(n22475), .B(n22476), .Y(n7285) );
  XOR2X4 U23429 ( .A(n7287), .B(n6922), .Y(n14100) );
  AOI21X4 U23430 ( .A0(n7306), .A1(n7289), .B0(n7288), .Y(n7287) );
  NOR2XL U23431 ( .A(n25010), .B(n25007), .Y(n7291) );
  XOR2X2 U23432 ( .A(n7294), .B(n11184), .Y(U1_U1_z0[6]) );
  AOI21X2 U23433 ( .A0(n11195), .A1(n11175), .B0(n11174), .Y(n7294) );
  OAI2BB2X4 U23434 ( .B0(n10162), .B1(n7295), .A0N(n8029), .A1N(W0[17]), .Y(
        n10153) );
  NOR2X4 U23435 ( .A(n8029), .B(W0[17]), .Y(n7295) );
  NOR2X4 U23436 ( .A(n8013), .B(W0[16]), .Y(n10162) );
  OAI21X1 U23437 ( .A0(n7296), .A1(n14138), .B0(n14137), .Y(n14139) );
  NAND3BX4 U23438 ( .AN(n8312), .B(n7762), .C(n7761), .Y(n7297) );
  AOI21X4 U23439 ( .A0(n7297), .A1(n9625), .B0(n9624), .Y(n11557) );
  NOR2X2 U23440 ( .A(n8425), .B(n8426), .Y(n8548) );
  AOI21XL U23441 ( .A0(n20194), .A1(n12331), .B0(n12330), .Y(n7304) );
  NAND4X2 U23442 ( .A(n7451), .B(n7797), .C(n14703), .D(n14690), .Y(n7307) );
  AOI21X1 U23443 ( .A0(n7359), .A1(n7795), .B0(n7794), .Y(n7309) );
  NAND2X1 U23444 ( .A(n14644), .B(n14645), .Y(n14693) );
  NAND2X1 U23445 ( .A(n17180), .B(n7314), .Y(n7313) );
  NAND3X1 U23446 ( .A(n7317), .B(n17177), .C(n7316), .Y(n7638) );
  NAND2XL U23447 ( .A(n9603), .B(n17178), .Y(n7316) );
  NAND2X1 U23448 ( .A(n17180), .B(n7318), .Y(n7317) );
  NOR2X2 U23449 ( .A(n7319), .B(n7749), .Y(n12339) );
  NAND2X1 U23450 ( .A(n7325), .B(n13504), .Y(n24919) );
  OR2X2 U23451 ( .A(n13505), .B(n24943), .Y(n7325) );
  NAND2X2 U23452 ( .A(n7330), .B(n7329), .Y(n9323) );
  CLKINVX3 U23453 ( .A(n7693), .Y(n7329) );
  NOR2X4 U23454 ( .A(n9464), .B(n9468), .Y(n7330) );
  INVX1 U23455 ( .A(n7332), .Y(n8246) );
  NAND2X2 U23456 ( .A(n7334), .B(n7333), .Y(n7332) );
  NOR2X2 U23457 ( .A(BOPA[37]), .B(BOPA[36]), .Y(n7333) );
  NOR2X4 U23458 ( .A(BOPA[35]), .B(BOPA[34]), .Y(n7334) );
  XOR2X4 U23459 ( .A(n10778), .B(n6903), .Y(U1_U2_z0[14]) );
  NAND2X2 U23460 ( .A(n10773), .B(n8254), .Y(n8256) );
  OAI21X4 U23461 ( .A0(n7339), .A1(n11427), .B0(n8269), .Y(U2_B_i[10]) );
  NAND2X2 U23462 ( .A(n7576), .B(n7334), .Y(n8268) );
  NAND3X1 U23463 ( .A(n9485), .B(n7640), .C(n7341), .Y(n7683) );
  OAI21X1 U23464 ( .A0(n6878), .A1(n10740), .B0(n10739), .Y(n10745) );
  OAI21X1 U23465 ( .A0(n6878), .A1(n10732), .B0(n10731), .Y(n10736) );
  OAI21XL U23466 ( .A0(n6878), .A1(n10714), .B0(n10713), .Y(n10719) );
  XNOR2X2 U23467 ( .A(n6878), .B(n7002), .Y(U1_U2_z0[16]) );
  OAI21XL U23468 ( .A0(n6878), .A1(n10855), .B0(n10854), .Y(n10856) );
  OAI21XL U23469 ( .A0(n6878), .A1(n10700), .B0(n10699), .Y(n10703) );
  NOR2X4 U23470 ( .A(n8028), .B(W2[17]), .Y(n7342) );
  NAND2X1 U23471 ( .A(n21188), .B(n21189), .Y(n7344) );
  NAND2X1 U23472 ( .A(n7345), .B(n12582), .Y(n12620) );
  AOI21X2 U23473 ( .A0(n7345), .A1(n12587), .B0(n12586), .Y(n12627) );
  NOR2X1 U23474 ( .A(n12581), .B(n12585), .Y(n7345) );
  NOR2XL U23475 ( .A(n7346), .B(n24654), .Y(n12600) );
  NAND2XL U23476 ( .A(n7346), .B(n24654), .Y(n22637) );
  NAND2XL U23477 ( .A(n13125), .B(n7346), .Y(n22342) );
  NAND2XL U23478 ( .A(n14555), .B(n7346), .Y(n22005) );
  AOI21X1 U23479 ( .A0(n23012), .A1(n23010), .B0(n23004), .Y(n7348) );
  OAI21X1 U23480 ( .A0(n23014), .A1(n23003), .B0(n23002), .Y(n23012) );
  NAND2XL U23481 ( .A(n7678), .B(n19072), .Y(n7353) );
  NAND3BX2 U23482 ( .AN(n9722), .B(n19072), .C(n7678), .Y(n7349) );
  NAND2X1 U23483 ( .A(n7677), .B(n7351), .Y(n7350) );
  NAND2BXL U23484 ( .AN(n7677), .B(n7353), .Y(n7352) );
  XNOR2X1 U23485 ( .A(n19070), .B(n7352), .Y(n19071) );
  NAND2X1 U23486 ( .A(n9480), .B(n7628), .Y(n7356) );
  NOR2X1 U23487 ( .A(n10185), .B(n10184), .Y(n7363) );
  NOR2X2 U23488 ( .A(n8139), .B(BOPD[28]), .Y(n10861) );
  NOR2X2 U23489 ( .A(n8137), .B(BOPD[29]), .Y(n10841) );
  OAI21X4 U23490 ( .A0(n11349), .A1(n7366), .B0(n7364), .Y(n9645) );
  AOI21X2 U23491 ( .A0(n11350), .A1(n7367), .B0(n7365), .Y(n7364) );
  OAI21X1 U23492 ( .A0(n11352), .A1(n11358), .B0(n11353), .Y(n7365) );
  NAND2X1 U23493 ( .A(n11351), .B(n7367), .Y(n7366) );
  NOR2X2 U23494 ( .A(n11352), .B(n11357), .Y(n7367) );
  NOR2X2 U23495 ( .A(n11362), .B(n11364), .Y(n11351) );
  AOI21X4 U23496 ( .A0(n11373), .A1(n7369), .B0(n7368), .Y(n11349) );
  OAI21X2 U23497 ( .A0(n11374), .A1(n11392), .B0(n11375), .Y(n7368) );
  NOR2X2 U23498 ( .A(n11391), .B(n11374), .Y(n7369) );
  NOR2X2 U23499 ( .A(n8079), .B(AOPC[29]), .Y(n11374) );
  OAI21X2 U23500 ( .A0(n9831), .A1(n9834), .B0(n9832), .Y(n7372) );
  NOR2X2 U23501 ( .A(n9831), .B(n9833), .Y(n7373) );
  NOR2BX2 U23502 ( .AN(U2_B_i[8]), .B(n7130), .Y(n11568) );
  OAI21X4 U23503 ( .A0(n7375), .A1(n11427), .B0(n9610), .Y(U2_B_i[8]) );
  XOR2X2 U23504 ( .A(n7576), .B(BOPA[34]), .Y(n7375) );
  NOR2X1 U23505 ( .A(n18549), .B(n18548), .Y(n18594) );
  AOI21X1 U23506 ( .A0(n18904), .A1(n7050), .B0(n7378), .Y(n7377) );
  NAND3X1 U23507 ( .A(n18905), .B(n18865), .C(n7050), .Y(n7379) );
  NAND2BX1 U23508 ( .AN(n14957), .B(n19998), .Y(n14958) );
  XOR2X4 U23509 ( .A(n7381), .B(n6894), .Y(n14957) );
  AOI21XL U23510 ( .A0(n24247), .A1(n24246), .B0(n24245), .Y(n24288) );
  NAND2BX1 U23511 ( .AN(n14562), .B(n24642), .Y(n25338) );
  NOR2X4 U23512 ( .A(n7946), .B(W2[22]), .Y(n10313) );
  NOR2X4 U23513 ( .A(n8039), .B(W0[22]), .Y(n10143) );
  AOI21X2 U23514 ( .A0(n10772), .A1(n8254), .B0(n7385), .Y(n8255) );
  OAI2BB1X2 U23515 ( .A0N(n7387), .A1N(n7386), .B0(n10769), .Y(n7385) );
  AOI21X2 U23516 ( .A0(n9913), .A1(n9896), .B0(n7391), .Y(n9904) );
  XOR2X4 U23517 ( .A(n9889), .B(n5769), .Y(U1_U2_z2[11]) );
  NOR2X4 U23518 ( .A(W1[23]), .B(W1[7]), .Y(n9968) );
  NOR2X4 U23519 ( .A(W1[22]), .B(W1[6]), .Y(n9982) );
  XOR2X4 U23520 ( .A(n9951), .B(n10215), .Y(U1_U1_z2[13]) );
  OAI21X4 U23521 ( .A0(n7403), .A1(n9986), .B0(n9987), .Y(n9960) );
  AOI21X2 U23522 ( .A0(n7397), .A1(n5772), .B0(n9727), .Y(n9955) );
  XOR2X1 U23523 ( .A(n7397), .B(n7008), .Y(U1_U1_z2[8]) );
  NAND2X2 U23524 ( .A(n8586), .B(n8542), .Y(n7399) );
  NAND2BX1 U23525 ( .AN(n16634), .B(n16633), .Y(n7401) );
  NAND2XL U23526 ( .A(n7410), .B(n22935), .Y(n22648) );
  NAND2XL U23527 ( .A(n7410), .B(n24646), .Y(n25039) );
  INVXL U23528 ( .A(n7410), .Y(n7409) );
  NAND2XL U23529 ( .A(n22939), .B(n7410), .Y(n23042) );
  NAND2XL U23530 ( .A(n5820), .B(n7410), .Y(n24767) );
  NAND3BX2 U23531 ( .AN(n9516), .B(n7413), .C(n7626), .Y(n17455) );
  NAND2X1 U23532 ( .A(n17477), .B(n9517), .Y(n7413) );
  AND2X2 U23533 ( .A(n7801), .B(n7034), .Y(n7796) );
  INVX1 U23534 ( .A(n9462), .Y(n7421) );
  OAI2BB1X4 U23535 ( .A0N(n7628), .A1N(n7421), .B0(n9461), .Y(n9472) );
  NAND2X2 U23536 ( .A(n9615), .B(n7422), .Y(n9552) );
  NOR2X4 U23537 ( .A(n8042), .B(W2[23]), .Y(n10269) );
  INVXL U23538 ( .A(n7423), .Y(n11576) );
  NOR2X2 U23539 ( .A(n11573), .B(n7423), .Y(n11567) );
  NOR2X4 U23540 ( .A(n9627), .B(U2_B_r[7]), .Y(n7423) );
  NAND2X1 U23541 ( .A(n13121), .B(n22361), .Y(n7424) );
  OAI21X1 U23542 ( .A0(n22362), .A1(n13120), .B0(n13119), .Y(n7425) );
  AOI21X1 U23543 ( .A0(n13133), .A1(n6934), .B0(n13132), .Y(n7427) );
  NAND2BX1 U23544 ( .AN(n22323), .B(n6934), .Y(n7428) );
  OAI21X1 U23545 ( .A0(n12134), .A1(n12122), .B0(n7429), .Y(n12082) );
  AOI21X2 U23546 ( .A0(n12067), .A1(n12089), .B0(n12066), .Y(n7429) );
  NAND2BX2 U23547 ( .AN(n9459), .B(n7629), .Y(n17524) );
  XOR2X1 U23548 ( .A(n16784), .B(n16785), .Y(n16786) );
  INVX2 U23549 ( .A(n14640), .Y(n7452) );
  NOR2X1 U23550 ( .A(n19967), .B(n14900), .Y(n20428) );
  XOR2X2 U23551 ( .A(n13788), .B(n6993), .Y(n14900) );
  XOR2X2 U23552 ( .A(n14695), .B(n6930), .Y(n19967) );
  OAI21XL U23553 ( .A0(n7446), .A1(n19571), .B0(n19572), .Y(n19569) );
  XOR2X4 U23554 ( .A(n10929), .B(n6895), .Y(U0_U2_z0[17]) );
  NAND2X1 U23555 ( .A(n7450), .B(n7449), .Y(n14702) );
  NOR2X1 U23556 ( .A(n12757), .B(n12758), .Y(n12874) );
  AOI21X1 U23557 ( .A0(n16812), .A1(n6900), .B0(n7956), .Y(n7456) );
  AND2X2 U23558 ( .A(n20014), .B(n14959), .Y(n16812) );
  NAND2X1 U23559 ( .A(n12695), .B(n12694), .Y(n12864) );
  OAI21XL U23560 ( .A0(n13934), .A1(n13939), .B0(n13935), .Y(n13954) );
  NAND2X1 U23561 ( .A(n7489), .B(n7491), .Y(n7488) );
  NOR2X1 U23562 ( .A(n7495), .B(n13621), .Y(n17305) );
  NAND2X1 U23563 ( .A(n13563), .B(n17322), .Y(n7496) );
  OAI21X1 U23564 ( .A0(n12978), .A1(n12977), .B0(n12976), .Y(n12979) );
  OAI21X1 U23565 ( .A0(n13585), .A1(n13588), .B0(n13592), .Y(n7512) );
  XOR2X4 U23566 ( .A(n7513), .B(n6896), .Y(n14951) );
  OAI21X2 U23567 ( .A0(n13030), .A1(n13026), .B0(n13027), .Y(n7513) );
  OAI21X1 U23568 ( .A0(n17350), .A1(n13557), .B0(n7516), .Y(n17322) );
  NAND2X1 U23569 ( .A(n14953), .B(n19544), .Y(n17358) );
  NAND2X1 U23570 ( .A(n17355), .B(n17359), .Y(n13557) );
  AND2X2 U23571 ( .A(U1_U0_y0[21]), .B(U1_U0_y2[21]), .Y(n8420) );
  NOR2X4 U23572 ( .A(n8419), .B(n8420), .Y(n8536) );
  AOI21X1 U23573 ( .A0(n7528), .A1(n19827), .B0(n19826), .Y(n19831) );
  XOR2X2 U23574 ( .A(U1_U0_y2[29]), .B(U1_U0_y0[29]), .Y(n8434) );
  AOI21XL U23575 ( .A0(n16944), .A1(n8631), .B0(n8630), .Y(n16942) );
  INVXL U23576 ( .A(n16635), .Y(n7537) );
  NAND2X1 U23577 ( .A(n7539), .B(n26905), .Y(n7538) );
  NAND2X1 U23578 ( .A(n7543), .B(n8173), .Y(n8174) );
  XOR2X4 U23579 ( .A(n8600), .B(n8599), .Y(n7543) );
  OAI2BB1X2 U23580 ( .A0N(n7548), .A1N(n26756), .B0(n7545), .Y(n26862) );
  NOR2X1 U23581 ( .A(n7547), .B(n7546), .Y(n7545) );
  OAI2BB1XL U23582 ( .A0N(n26755), .A1N(n26756), .B0(n26754), .Y(n26757) );
  NAND2BX1 U23583 ( .AN(n22459), .B(n22460), .Y(n7555) );
  OAI21X4 U23584 ( .A0(n13442), .A1(n13447), .B0(n13443), .Y(n13430) );
  NOR2X4 U23585 ( .A(n13276), .B(n13275), .Y(n13442) );
  OAI21X2 U23586 ( .A0(n13481), .A1(n13477), .B0(n13478), .Y(n13485) );
  NAND2X1 U23587 ( .A(n7558), .B(n25303), .Y(n7557) );
  OR2X2 U23588 ( .A(n25664), .B(n25302), .Y(n7558) );
  NOR2X2 U23589 ( .A(n8181), .B(BOPC[40]), .Y(n11123) );
  AOI21X4 U23590 ( .A0(n7564), .A1(n11107), .B0(n7563), .Y(n8289) );
  OAI21X2 U23591 ( .A0(n8288), .A1(n11139), .B0(n8287), .Y(n7563) );
  NAND2XL U23592 ( .A(n7565), .B(n22913), .Y(n22673) );
  NOR2X1 U23593 ( .A(n7565), .B(n24615), .Y(n24796) );
  NAND2XL U23594 ( .A(n24625), .B(n7565), .Y(n24626) );
  NOR2XL U23595 ( .A(n24625), .B(n7565), .Y(n24627) );
  NAND2XL U23596 ( .A(n22922), .B(n7565), .Y(n23069) );
  XOR2X4 U23597 ( .A(n8960), .B(n8959), .Y(n7565) );
  AOI21X4 U23598 ( .A0(n10645), .A1(n8270), .B0(n7567), .Y(n7566) );
  NAND2X4 U23599 ( .A(n10646), .B(n8270), .Y(n7568) );
  NAND2X1 U23600 ( .A(n13398), .B(n7080), .Y(n22526) );
  OAI21X1 U23601 ( .A0(n13405), .A1(n13410), .B0(n13406), .Y(n7570) );
  NOR2X4 U23602 ( .A(n13405), .B(n13409), .Y(n7571) );
  OAI21X1 U23603 ( .A0(n13384), .A1(n13389), .B0(n13385), .Y(n7572) );
  OAI21X1 U23604 ( .A0(n13469), .A1(n13468), .B0(n13467), .Y(n7573) );
  OAI2BB1X2 U23605 ( .A0N(n22434), .A1N(n5854), .B0(n7575), .Y(n22498) );
  INVX1 U23606 ( .A(n22442), .Y(n7575) );
  NAND3XL U23607 ( .A(n9607), .B(n7576), .C(n28712), .Y(n8247) );
  OAI2BB1X2 U23608 ( .A0N(n24784), .A1N(n24415), .B0(n7577), .Y(n4376) );
  XOR2X4 U23609 ( .A(n7578), .B(n10127), .Y(U0_U0_z1[14]) );
  XOR2X4 U23610 ( .A(n7582), .B(n7581), .Y(U1_U1_z1[13]) );
  INVX1 U23611 ( .A(n14056), .Y(n13359) );
  NAND2X2 U23612 ( .A(n7587), .B(n7585), .Y(n24501) );
  AOI21X2 U23613 ( .A0(n7602), .A1(n7601), .B0(n7599), .Y(n7585) );
  INVX1 U23614 ( .A(U0_U0_y0[19]), .Y(n7605) );
  OR2X2 U23615 ( .A(n13354), .B(n13352), .Y(n7610) );
  AOI21X1 U23616 ( .A0(n22494), .A1(n14050), .B0(n14049), .Y(n22439) );
  NOR2XL U23617 ( .A(n14047), .B(U2_A_i_d[17]), .Y(n22492) );
  OAI21X2 U23618 ( .A0(n13416), .A1(n13422), .B0(n13417), .Y(n13403) );
  NOR2BX2 U23619 ( .AN(n13426), .B(n13402), .Y(n7724) );
  OAI21XL U23620 ( .A0(n24888), .A1(n14002), .B0(n24460), .Y(n14004) );
  NAND2X2 U23621 ( .A(n6875), .B(W0[18]), .Y(n10154) );
  OAI21XL U23622 ( .A0(n24992), .A1(n24714), .B0(n24715), .Y(n9210) );
  INVX1 U23623 ( .A(n9194), .Y(n24721) );
  XNOR2X2 U23624 ( .A(n9203), .B(n9193), .Y(n24680) );
  INVX1 U23625 ( .A(n14129), .Y(n14136) );
  NAND2X1 U23626 ( .A(n12546), .B(n12545), .Y(n12560) );
  MXI2X1 U23627 ( .A(n7736), .B(U0_pipe15[26]), .S0(n8053), .Y(n4610) );
  NOR2X2 U23628 ( .A(n22952), .B(n23003), .Y(n22954) );
  NOR2X4 U23629 ( .A(n10650), .B(n10647), .Y(n8270) );
  OAI21X2 U23630 ( .A0(n10624), .A1(n10630), .B0(n10625), .Y(n8272) );
  XNOR2X1 U23631 ( .A(n9844), .B(n10188), .Y(U0_U0_z2[4]) );
  NOR2X1 U23632 ( .A(n26698), .B(n26701), .Y(n26753) );
  NAND2X1 U23633 ( .A(n21518), .B(n21524), .Y(n21526) );
  CLKINVX3 U23634 ( .A(n26820), .Y(n21480) );
  NAND2X1 U23635 ( .A(n8072), .B(AOPB[31]), .Y(n10493) );
  OAI21X2 U23636 ( .A0(n10522), .A1(n10409), .B0(n10410), .Y(n10408) );
  OAI21X2 U23637 ( .A0(n11389), .A1(n11245), .B0(n11244), .Y(n11249) );
  NAND2X1 U23638 ( .A(n13455), .B(n13414), .Y(n13457) );
  NOR2XL U23639 ( .A(n13452), .B(U2_A_r_d[16]), .Y(n13408) );
  AOI21X1 U23640 ( .A0(n24450), .A1(n13464), .B0(n13463), .Y(n13465) );
  XOR2X2 U23641 ( .A(n13441), .B(n13440), .Y(n14102) );
  NOR2X2 U23642 ( .A(n11433), .B(n11543), .Y(n11435) );
  OAI21X2 U23643 ( .A0(n13441), .A1(n13437), .B0(n13438), .Y(n13436) );
  XNOR2X1 U23644 ( .A(n22763), .B(n22762), .Y(n22764) );
  XNOR2X1 U23645 ( .A(n22749), .B(n22748), .Y(n22750) );
  XNOR2X1 U23646 ( .A(n22757), .B(n22756), .Y(n22758) );
  OAI21X1 U23647 ( .A0(n21830), .A1(n21797), .B0(n21796), .Y(n21823) );
  AOI21X1 U23648 ( .A0(n25048), .A1(n9012), .B0(n9011), .Y(n25006) );
  NOR2X1 U23649 ( .A(n24796), .B(n24802), .Y(n9007) );
  INVX2 U23650 ( .A(n17230), .Y(n13719) );
  NAND2XL U23651 ( .A(n25216), .B(U2_A_r_d[11]), .Y(n25480) );
  NOR2X2 U23652 ( .A(n11444), .B(n11526), .Y(n11513) );
  AOI2BB1X2 U23653 ( .A0N(n9430), .A1N(n9433), .B0(n7656), .Y(n7655) );
  CLKINVX3 U23654 ( .A(n14421), .Y(n14369) );
  AOI21X1 U23655 ( .A0(n6980), .A1(n25597), .B0(n25482), .Y(n25483) );
  NAND2X1 U23656 ( .A(n9585), .B(n17232), .Y(n7621) );
  AOI21X1 U23657 ( .A0(n12536), .A1(n12535), .B0(n12534), .Y(n12537) );
  NOR2X1 U23658 ( .A(n9864), .B(n9868), .Y(n9871) );
  ADDHX2 U23659 ( .A(U2_U0_y2[29]), .B(U2_U0_y0[29]), .CO(n23981), .S(n23937)
         );
  NAND2X1 U23660 ( .A(n23939), .B(n23938), .Y(n24038) );
  OAI21X2 U23661 ( .A0(n10336), .A1(n10296), .B0(n10295), .Y(n10297) );
  NOR2X2 U23662 ( .A(n9812), .B(n9810), .Y(n9825) );
  NAND2X1 U23663 ( .A(n7835), .B(n7833), .Y(n7917) );
  OAI21X2 U23664 ( .A0(n10114), .A1(n10142), .B0(n10113), .Y(n10115) );
  NOR2X2 U23665 ( .A(n8167), .B(BOPC[27]), .Y(n11218) );
  AOI21X2 U23666 ( .A0(n22954), .A1(n23000), .B0(n22953), .Y(n22955) );
  NAND2X1 U23667 ( .A(n12565), .B(n12564), .Y(n12584) );
  XNOR2X4 U23668 ( .A(n10403), .B(n10402), .Y(U0_U0_z0[18]) );
  NAND2X1 U23669 ( .A(n7990), .B(AOPB[40]), .Y(n10431) );
  NAND2X2 U23670 ( .A(n8138), .B(BOPC[28]), .Y(n11203) );
  OAI21X4 U23671 ( .A0(n7197), .A1(n8331), .B0(n8330), .Y(n8334) );
  NAND2X1 U23672 ( .A(n8062), .B(AOPC[34]), .Y(n11345) );
  XNOR2X4 U23673 ( .A(n10883), .B(n10882), .Y(U0_U2_z0[24]) );
  XNOR2X2 U23674 ( .A(n11234), .B(n11233), .Y(U0_U1_z0[25]) );
  XOR2X2 U23675 ( .A(n11501), .B(n11500), .Y(U2_U0_z0[21]) );
  NOR2X4 U23676 ( .A(n10112), .B(n10146), .Y(n10141) );
  AOI21X2 U23677 ( .A0(n11582), .A1(n11580), .B0(n11574), .Y(n11578) );
  XNOR2X2 U23678 ( .A(n8309), .B(BOPA[28]), .Y(n8305) );
  INVX1 U23679 ( .A(n24863), .Y(n24864) );
  OR2X2 U23680 ( .A(n14048), .B(U2_A_r_d[18]), .Y(n24469) );
  AOI21X1 U23681 ( .A0(n8078), .A1(n24454), .B0(n13460), .Y(n13461) );
  NOR2X2 U23682 ( .A(n8443), .B(n8442), .Y(n8592) );
  OAI21XL U23683 ( .A0(n8614), .A1(n16960), .B0(n8613), .Y(n8615) );
  OAI21X1 U23684 ( .A0(n11562), .A1(n11569), .B0(n11563), .Y(n9630) );
  OAI21X2 U23685 ( .A0(n11555), .A1(n11543), .B0(n11542), .Y(n11547) );
  OAI21X1 U23686 ( .A0(n11472), .A1(n11462), .B0(n11475), .Y(n11457) );
  OAI21X1 U23687 ( .A0(n19523), .A1(n19664), .B0(n19522), .Y(n19639) );
  INVX1 U23688 ( .A(n19578), .Y(n19591) );
  AOI21X2 U23689 ( .A0(n10190), .A1(n10149), .B0(n10148), .Y(n10152) );
  OAI21XL U23690 ( .A0(n25689), .A1(n25684), .B0(n25683), .Y(n25686) );
  OAI21X1 U23691 ( .A0(n9140), .A1(n25028), .B0(n9139), .Y(n25007) );
  OR2X4 U23692 ( .A(n24619), .B(n14532), .Y(n25728) );
  OAI21X1 U23693 ( .A0(n25724), .A1(n12173), .B0(n12172), .Y(n12174) );
  INVX4 U23694 ( .A(n11349), .Y(n11372) );
  AOI21X1 U23695 ( .A0(n25722), .A1(n25679), .B0(n25678), .Y(n25693) );
  OAI21X1 U23696 ( .A0(n11361), .A1(n11357), .B0(n11358), .Y(n11356) );
  NOR2X1 U23697 ( .A(n13698), .B(U1_A_r_d0[17]), .Y(n19423) );
  AND2X2 U23698 ( .A(n24644), .B(n24654), .Y(n8086) );
  AOI21XL U23699 ( .A0(n21849), .A1(n21845), .B0(n21844), .Y(n21846) );
  AOI21XL U23700 ( .A0(n25168), .A1(n25161), .B0(n25160), .Y(n25164) );
  NAND2X1 U23701 ( .A(n14225), .B(n14224), .Y(n14362) );
  CLKINVX2 U23702 ( .A(n25155), .Y(n25205) );
  CLKINVX2 U23703 ( .A(n21839), .Y(n21879) );
  OAI21X2 U23704 ( .A0(n10469), .A1(n10475), .B0(n10470), .Y(n10462) );
  XNOR2X1 U23705 ( .A(n10771), .B(n10770), .Y(U1_U2_z0[15]) );
  OAI21X1 U23706 ( .A0(n26456), .A1(n26455), .B0(n26454), .Y(n26598) );
  XNOR2X4 U23707 ( .A(n11283), .B(n11282), .Y(U0_U1_z0[18]) );
  BUFX8 U23708 ( .A(n8343), .Y(n11389) );
  AOI21X1 U23709 ( .A0(n14034), .A1(n14033), .B0(n14032), .Y(n22522) );
  NAND2X1 U23710 ( .A(n9305), .B(n9304), .Y(n9430) );
  NOR2X1 U23711 ( .A(n9504), .B(U1_A_i_d0[15]), .Y(n17507) );
  CMPR22X1 U23712 ( .A(U1_U0_y2[35]), .B(U1_U0_y0[35]), .CO(n8451), .S(n8447)
         );
  AOI21X4 U23713 ( .A0(n10260), .A1(n10259), .B0(n10258), .Y(n10263) );
  NAND2X1 U23714 ( .A(n22931), .B(n14550), .Y(n22322) );
  AOI21X1 U23715 ( .A0(n14141), .A1(n14140), .B0(n14139), .Y(n14142) );
  OAI21XL U23716 ( .A0(n18252), .A1(n18483), .B0(n18492), .Y(n18301) );
  NOR2X1 U23717 ( .A(n18040), .B(n18044), .Y(n18047) );
  CLKINVX3 U23718 ( .A(n24040), .Y(n18650) );
  XNOR2X1 U23719 ( .A(n27039), .B(n27038), .Y(n27041) );
  OAI21X2 U23720 ( .A0(n11542), .A1(n11433), .B0(n11432), .Y(n11434) );
  NAND2X2 U23721 ( .A(W2[5]), .B(W2[21]), .Y(n9908) );
  NAND2X1 U23722 ( .A(n8433), .B(n8432), .Y(n8577) );
  OR2X2 U23723 ( .A(n7627), .B(U1_A_r_d0[14]), .Y(n9692) );
  OAI21X1 U23724 ( .A0(n9432), .A1(n9431), .B0(n9430), .Y(n7620) );
  NAND2X2 U23725 ( .A(n7622), .B(n7665), .Y(n9532) );
  NAND2X1 U23726 ( .A(n7622), .B(n7666), .Y(n7662) );
  INVX1 U23727 ( .A(n9717), .Y(n13716) );
  INVX2 U23728 ( .A(n13710), .Y(n9712) );
  XOR2X4 U23729 ( .A(n7634), .B(n6961), .Y(n13710) );
  NAND2X2 U23730 ( .A(n7668), .B(n7725), .Y(n7634) );
  OAI21X2 U23731 ( .A0(n9518), .A1(n9521), .B0(n9522), .Y(n9335) );
  AOI21X2 U23732 ( .A0(n9332), .A1(n9481), .B0(n7635), .Y(n9518) );
  OAI21X1 U23733 ( .A0(n7636), .A1(n9487), .B0(n9483), .Y(n7635) );
  XOR2X1 U23734 ( .A(n7638), .B(n7012), .Y(n7637) );
  INVXL U23735 ( .A(n7652), .Y(n7644) );
  INVXL U23736 ( .A(n9547), .Y(n7647) );
  XNOR2XL U23737 ( .A(n14974), .B(U1_A_i_d0[25]), .Y(n7654) );
  NAND2X2 U23738 ( .A(n9360), .B(n7741), .Y(n7660) );
  NAND2X1 U23739 ( .A(n7662), .B(n9529), .Y(n9534) );
  CLKINVX3 U23740 ( .A(n9335), .Y(n7668) );
  INVXL U23741 ( .A(n7671), .Y(n17469) );
  NAND2XL U23742 ( .A(n9491), .B(n7673), .Y(n7672) );
  XOR2X1 U23743 ( .A(n14974), .B(n29007), .Y(n7675) );
  NAND2X1 U23744 ( .A(n7679), .B(n9689), .Y(n19105) );
  NAND3X1 U23745 ( .A(n9490), .B(n7748), .C(n9487), .Y(n7682) );
  NAND2X1 U23746 ( .A(n7691), .B(n7689), .Y(n7694) );
  NOR2X4 U23747 ( .A(n9322), .B(n7029), .Y(n9464) );
  NOR2X2 U23748 ( .A(n9306), .B(n9307), .Y(n9433) );
  NAND2BX1 U23749 ( .AN(n13694), .B(n7077), .Y(n17221) );
  AOI21X1 U23750 ( .A0(n17209), .A1(n13725), .B0(n13724), .Y(n17200) );
  CLKINVX2 U23751 ( .A(n13720), .Y(n7700) );
  XOR2X1 U23752 ( .A(n25528), .B(n29009), .Y(n7710) );
  NAND2X1 U23753 ( .A(n21193), .B(n21192), .Y(n21306) );
  NAND2X1 U23754 ( .A(n7696), .B(n7082), .Y(n9705) );
  NOR2X2 U23755 ( .A(n11316), .B(n11310), .Y(n11302) );
  NOR2X2 U23756 ( .A(n7954), .B(AOPC[39]), .Y(n11316) );
  NOR2X2 U23757 ( .A(n10507), .B(n10502), .Y(n8212) );
  NAND2X2 U23758 ( .A(n13275), .B(n13276), .Y(n13443) );
  OAI21X1 U23759 ( .A0(n7720), .A1(n24439), .B0(n13487), .Y(n24431) );
  NOR2X1 U23760 ( .A(n5846), .B(n24693), .Y(n7728) );
  NOR2X1 U23761 ( .A(n12225), .B(n12229), .Y(n12242) );
  XOR2X1 U23762 ( .A(n5815), .B(n25286), .Y(n7732) );
  AOI2BB1X2 U23763 ( .A0N(n12339), .A1N(n12338), .B0(n7752), .Y(n12340) );
  OAI2BB1X2 U23764 ( .A0N(n24784), .A1N(n22971), .B0(n7754), .Y(n4522) );
  NAND2X1 U23765 ( .A(n11593), .B(n11591), .Y(n7761) );
  NAND2X1 U23766 ( .A(n8180), .B(BOPC[41]), .Y(n11115) );
  NOR2X2 U23767 ( .A(n7767), .B(BOPA[45]), .Y(n11415) );
  XOR2X2 U23768 ( .A(n7770), .B(n10969), .Y(U0_U2_z0[12]) );
  AOI21X1 U23769 ( .A0(n10988), .A1(n10955), .B0(n10957), .Y(n7770) );
  OAI21X1 U23770 ( .A0(n8289), .A1(n11086), .B0(n11085), .Y(n11091) );
  OAI21XL U23771 ( .A0(n8289), .A1(n11095), .B0(n11094), .Y(n11099) );
  OAI21X1 U23772 ( .A0(n8289), .A1(n11074), .B0(n11073), .Y(n11079) );
  OAI21XL U23773 ( .A0(n8289), .A1(n11054), .B0(n11053), .Y(n11059) );
  OAI21X1 U23774 ( .A0(n8296), .A1(n8289), .B0(n8295), .Y(n8298) );
  OAI21XL U23775 ( .A0(n8289), .A1(n11216), .B0(n11215), .Y(n11217) );
  NOR2X2 U23776 ( .A(n7056), .B(AOPC[33]), .Y(n11352) );
  NAND2X1 U23777 ( .A(n9068), .B(n9067), .Y(n9165) );
  NOR2X1 U23778 ( .A(n5815), .B(n5814), .Y(n24987) );
  XOR2X4 U23779 ( .A(n7771), .B(n10144), .Y(U0_U0_z2[7]) );
  OAI21X2 U23780 ( .A0(n9836), .A1(n9833), .B0(n9834), .Y(n7771) );
  OAI21XL U23781 ( .A0(n9075), .A1(n7774), .B0(n9072), .Y(n7773) );
  AOI21X4 U23782 ( .A0(n11512), .A1(n11447), .B0(n7778), .Y(n11448) );
  NOR2X2 U23783 ( .A(n11507), .B(n11514), .Y(n11447) );
  NOR2X2 U23784 ( .A(n11446), .B(U2_B_r[19]), .Y(n11507) );
  OAI21X4 U23785 ( .A0(n11527), .A1(n11444), .B0(n7779), .Y(n11512) );
  AOI2BB1X4 U23786 ( .A0N(n11437), .A1N(n11539), .B0(n11440), .Y(n11527) );
  XOR2X2 U23787 ( .A(n7785), .B(n13663), .Y(n7861) );
  OAI21X1 U23788 ( .A0(n13660), .A1(n13659), .B0(n13658), .Y(n7785) );
  AOI21X4 U23789 ( .A0(n13646), .A1(n13634), .B0(n13645), .Y(n13660) );
  OAI21X4 U23790 ( .A0(n13063), .A1(n7788), .B0(n7787), .Y(n13593) );
  AOI21X4 U23791 ( .A0(n13062), .A1(n7927), .B0(n7926), .Y(n7787) );
  NOR2X4 U23792 ( .A(n7928), .B(n12979), .Y(n13063) );
  XOR2X1 U23793 ( .A(n7789), .B(n19249), .Y(n19250) );
  AOI21X1 U23794 ( .A0(n19234), .A1(n7790), .B0(n7275), .Y(n7789) );
  INVXL U23795 ( .A(n7793), .Y(n14742) );
  NAND2X1 U23796 ( .A(n14741), .B(n7793), .Y(n7801) );
  NOR2X1 U23797 ( .A(n14739), .B(n7793), .Y(n14706) );
  NOR2X2 U23798 ( .A(n14636), .B(n14637), .Y(n7793) );
  NAND2X1 U23799 ( .A(n14738), .B(n14741), .Y(n7800) );
  NOR2X1 U23800 ( .A(n14634), .B(n14635), .Y(n14739) );
  INVXL U23801 ( .A(n19620), .Y(n19625) );
  OR2X2 U23802 ( .A(n19281), .B(n19620), .Y(n19549) );
  NAND2BX1 U23803 ( .AN(n19539), .B(n19540), .Y(n19616) );
  NAND2X2 U23804 ( .A(n14637), .B(n14636), .Y(n14741) );
  XOR2X1 U23805 ( .A(n7811), .B(n7810), .Y(n7809) );
  CLKINVX3 U23806 ( .A(n14785), .Y(n19979) );
  XOR2X2 U23807 ( .A(n7812), .B(n6921), .Y(n14785) );
  XNOR2X1 U23808 ( .A(n20333), .B(n7814), .Y(n7813) );
  INVXL U23809 ( .A(n7825), .Y(n7824) );
  AOI21X4 U23810 ( .A0(n7930), .A1(n12893), .B0(n7828), .Y(n7929) );
  NOR2X1 U23811 ( .A(n17604), .B(n14512), .Y(n7829) );
  NOR2XL U23812 ( .A(n14956), .B(n7843), .Y(n20000) );
  NAND2X1 U23813 ( .A(n5865), .B(n7843), .Y(n19268) );
  NAND2X1 U23814 ( .A(n14633), .B(n14717), .Y(n7851) );
  NOR2XL U23815 ( .A(n7861), .B(n20333), .Y(n7853) );
  NAND2X1 U23816 ( .A(n12763), .B(n12807), .Y(n12901) );
  AOI21XL U23817 ( .A0(n17304), .A1(n13624), .B0(n13623), .Y(n17302) );
  NAND2X1 U23818 ( .A(n7214), .B(n14108), .Y(n7862) );
  OAI21X4 U23819 ( .A0(n13627), .A1(n13626), .B0(n13625), .Y(n13639) );
  NAND2X1 U23820 ( .A(n13084), .B(n13083), .Y(n13580) );
  NOR2X2 U23821 ( .A(n13856), .B(n13857), .Y(n13872) );
  AND2X2 U23822 ( .A(n13069), .B(n7915), .Y(n7967) );
  AOI21X2 U23823 ( .A0(n13573), .A1(n13071), .B0(n13051), .Y(n7874) );
  OAI21X4 U23824 ( .A0(n13633), .A1(n13632), .B0(n13631), .Y(n13646) );
  NOR2X1 U23825 ( .A(n17324), .B(n13562), .Y(n13563) );
  XOR2X2 U23826 ( .A(n7925), .B(n13091), .Y(n19259) );
  NAND2X1 U23827 ( .A(n13565), .B(n13570), .Y(n13598) );
  INVX1 U23828 ( .A(n14780), .Y(n7883) );
  NAND2X1 U23829 ( .A(n14654), .B(n14655), .Y(n14780) );
  NAND2X1 U23830 ( .A(n14666), .B(n14667), .Y(n14805) );
  XOR2X1 U23831 ( .A(n19568), .B(n19567), .Y(n7902) );
  NAND2X1 U23832 ( .A(n17341), .B(n17345), .Y(n17324) );
  NAND2X1 U23833 ( .A(n19565), .B(n19566), .Y(n19575) );
  NOR2XL U23834 ( .A(n13087), .B(n13086), .Y(n7909) );
  NOR2XL U23835 ( .A(n13046), .B(n13041), .Y(n13599) );
  OAI21X2 U23836 ( .A0(n12949), .A1(n12948), .B0(n12947), .Y(n12998) );
  NAND2XL U23837 ( .A(n7915), .B(n14957), .Y(n17340) );
  OAI21X2 U23838 ( .A0(n13060), .A1(n13061), .B0(n13059), .Y(n7926) );
  NOR2X4 U23839 ( .A(n13061), .B(n13056), .Y(n7927) );
  AND2X4 U23840 ( .A(n12981), .B(n12980), .Y(n7928) );
  NOR2X4 U23841 ( .A(n12986), .B(n12987), .Y(n13056) );
  NOR2X4 U23842 ( .A(n12988), .B(n12989), .Y(n13061) );
  XOR2X2 U23843 ( .A(n7936), .B(n6959), .Y(U1_U0_z0[11]) );
  OAI21XL U23844 ( .A0(n9108), .A1(n9105), .B0(n9109), .Y(n9058) );
  NAND2X1 U23845 ( .A(n9056), .B(n9057), .Y(n9109) );
  INVX1 U23846 ( .A(U2_B_i[4]), .Y(n8313) );
  NOR2X1 U23847 ( .A(n10634), .B(n10639), .Y(n10627) );
  NOR2X2 U23848 ( .A(n10621), .B(n10624), .Y(n8273) );
  NOR2X4 U23849 ( .A(W0[6]), .B(W0[22]), .Y(n9833) );
  NOR2X4 U23850 ( .A(W0[23]), .B(W0[7]), .Y(n9831) );
  NAND2X1 U23851 ( .A(n12394), .B(n25337), .Y(n25324) );
  AOI21X1 U23852 ( .A0(n18707), .A1(n18706), .B0(n18705), .Y(n18815) );
  NOR2X1 U23853 ( .A(n14922), .B(n14900), .Y(n17140) );
  XNOR2X1 U23854 ( .A(n24428), .B(n24427), .Y(n24429) );
  XNOR2X1 U23855 ( .A(n24443), .B(n24442), .Y(n24444) );
  OR2X2 U23856 ( .A(n22949), .B(n24666), .Y(n23006) );
  CMPR22X1 U23857 ( .A(U2_U0_y2[35]), .B(U2_U0_y0[35]), .CO(n24289), .S(n24249) );
  NAND2X1 U23858 ( .A(n18054), .B(n18053), .Y(n18138) );
  OAI211X4 U23859 ( .A0(n28752), .A1(n27772), .B0(n27083), .C0(n27082), .Y(
        A0_addr[0]) );
  AOI21X4 U23860 ( .A0(n8284), .A1(n11156), .B0(n8283), .Y(n11139) );
  INVX1 U23861 ( .A(n24421), .Y(n24447) );
  XOR2X4 U23862 ( .A(n11525), .B(n11524), .Y(U2_U0_z0[17]) );
  AOI21X1 U23863 ( .A0(n24469), .A1(n13520), .B0(n13519), .Y(n13999) );
  AOI21X1 U23864 ( .A0(n5788), .A1(n19642), .B0(n19533), .Y(n19534) );
  NOR2X2 U23865 ( .A(n18191), .B(n18190), .Y(n18248) );
  OAI21XL U23866 ( .A0(n10574), .A1(n10583), .B0(n10575), .Y(n9560) );
  NAND2X1 U23867 ( .A(n8171), .B(BOPB[44]), .Y(n10583) );
  NOR2X1 U23868 ( .A(n8093), .B(AOPC[48]), .Y(n11256) );
  AOI21X1 U23869 ( .A0(n13025), .A1(n17657), .B0(n13036), .Y(n17644) );
  OAI21XL U23870 ( .A0(n11224), .A1(n11263), .B0(n11223), .Y(n11251) );
  INVXL U23871 ( .A(n12601), .Y(n12611) );
  AOI21XL U23872 ( .A0(n19648), .A1(n19310), .B0(n19642), .Y(n19645) );
  INVX1 U23873 ( .A(n22744), .Y(n22767) );
  XNOR2X2 U23874 ( .A(n10425), .B(n10424), .Y(U0_U0_z0[15]) );
  INVX1 U23875 ( .A(n11549), .Y(n9636) );
  INVX1 U23876 ( .A(n11552), .Y(n9637) );
  ADDHX2 U23877 ( .A(U1_U1_y0[30]), .B(U1_U1_y2[30]), .CO(n13065), .S(n12988)
         );
  NAND2XL U23878 ( .A(n23017), .B(n23022), .Y(n23003) );
  AOI21X1 U23879 ( .A0(n23017), .A1(n23015), .B0(n22948), .Y(n23002) );
  NOR2X1 U23880 ( .A(n13462), .B(n24453), .Y(n13464) );
  OAI21XL U23881 ( .A0(n22836), .A1(n22809), .B0(n22808), .Y(n22818) );
  INVX1 U23882 ( .A(n9999), .Y(n9727) );
  NAND2X1 U23883 ( .A(n8121), .B(BOPD[34]), .Y(n10814) );
  NAND2X1 U23884 ( .A(n8118), .B(BOPD[35]), .Y(n10809) );
  NAND2X1 U23885 ( .A(n21426), .B(n21425), .Y(n21520) );
  OAI21XL U23886 ( .A0(n24535), .A1(n24505), .B0(n24504), .Y(n24515) );
  NAND2X1 U23887 ( .A(n22494), .B(n5818), .Y(n22433) );
  NOR2X1 U23888 ( .A(n23636), .B(n23635), .Y(n23685) );
  INVX1 U23889 ( .A(n24160), .Y(n18768) );
  INVX1 U23890 ( .A(n22357), .Y(n22351) );
  NOR2X2 U23891 ( .A(n21019), .B(n21018), .Y(n21066) );
  INVX1 U23892 ( .A(n25129), .Y(n25153) );
  NAND2X1 U23893 ( .A(n25377), .B(n6992), .Y(n12382) );
  NOR2X1 U23894 ( .A(n8157), .B(BOPB[48]), .Y(n10550) );
  AOI21X1 U23895 ( .A0(n22649), .A1(n22647), .B0(n12613), .Y(n22633) );
  INVX1 U23896 ( .A(n12606), .Y(n22649) );
  AND2X2 U23897 ( .A(n14562), .B(n22932), .Y(n8105) );
  OAI21X1 U23898 ( .A0(n11389), .A1(n11255), .B0(n11254), .Y(n11260) );
  CMPR22X1 U23899 ( .A(U0_U0_y2[35]), .B(U0_U0_y0[35]), .CO(n14262), .S(n14257) );
  AOI21X1 U23900 ( .A0(n13169), .A1(n6987), .B0(n13168), .Y(n22304) );
  OAI21XL U23901 ( .A0(n19662), .A1(n19641), .B0(n19640), .Y(n19648) );
  ADDHX2 U23902 ( .A(U0_U0_y2[31]), .B(U0_U0_y0[31]), .CO(n14251), .S(n14248)
         );
  XNOR2X4 U23903 ( .A(n11239), .B(n11238), .Y(U0_U1_z0[24]) );
  OAI21X2 U23904 ( .A0(n11389), .A1(n11236), .B0(n11235), .Y(n11239) );
  ADDHX2 U23905 ( .A(U0_U1_y2[21]), .B(U0_U1_y0[21]), .CO(n12532), .S(n12477)
         );
  AOI21XL U23906 ( .A0(n22370), .A1(n22365), .B0(n22364), .Y(n22367) );
  CMPR22X1 U23907 ( .A(U1_U0_y1[35]), .B(U1_U0_y0[35]), .CO(n9337), .S(n9333)
         );
  NAND2X1 U23908 ( .A(n24745), .B(n5794), .Y(n24732) );
  NOR2X1 U23909 ( .A(n24036), .B(n24039), .Y(n24091) );
  ADDHX2 U23910 ( .A(U0_U0_y1[20]), .B(U0_U0_y0[20]), .CO(n13256), .S(n13254)
         );
  AOI21X1 U23911 ( .A0(n25705), .A1(n12232), .B0(n12231), .Y(n12233) );
  XNOR2X4 U23912 ( .A(n11309), .B(n11308), .Y(U0_U1_z0[14]) );
  ADDHX2 U23913 ( .A(U1_U0_y2[30]), .B(U1_U0_y0[30]), .CO(n8439), .S(n8436) );
  INVX1 U23914 ( .A(n13112), .Y(n22365) );
  NOR2XL U23915 ( .A(n22918), .B(n14533), .Y(n13112) );
  AOI21X1 U23916 ( .A0(n12575), .A1(n12574), .B0(n12573), .Y(n22658) );
  NOR2X1 U23917 ( .A(n13147), .B(n13150), .Y(n13152) );
  INVX1 U23918 ( .A(n25550), .Y(n25592) );
  OAI21X1 U23919 ( .A0(n10559), .A1(n10566), .B0(n10560), .Y(n10547) );
  ADDHX2 U23920 ( .A(U1_U0_y1[30]), .B(U1_U0_y0[30]), .CO(n9325), .S(n9322) );
  OAI211X4 U23921 ( .A0(n28752), .A1(n27379), .B0(n27072), .C0(n27071), .Y(
        A2_addr[0]) );
  NAND2X1 U23922 ( .A(n14647), .B(n14646), .Y(n14766) );
  OAI211X4 U23923 ( .A0(n28753), .A1(n27379), .B0(n27075), .C0(n27074), .Y(
        A2_addr[1]) );
  CMPR22X1 U23924 ( .A(U2_U0_y2[33]), .B(U2_U0_y0[33]), .CO(n24206), .S(n24160) );
  OAI21X1 U23925 ( .A0(n10997), .A1(n10959), .B0(n10958), .Y(n10964) );
  NOR2X1 U23926 ( .A(n11128), .B(n11134), .Y(n11120) );
  OAI211X4 U23927 ( .A0(n28755), .A1(n27379), .B0(n27077), .C0(n27076), .Y(
        A2_addr[2]) );
  OAI211X4 U23928 ( .A0(n28754), .A1(n27379), .B0(n27080), .C0(n27079), .Y(
        A2_addr[4]) );
  ADDHX2 U23929 ( .A(U2_U0_y1[31]), .B(U2_U0_y0[31]), .CO(n26759), .S(n26703)
         );
  ADDHX2 U23930 ( .A(U2_U0_y2[31]), .B(U2_U0_y0[31]), .CO(n24097), .S(n24041)
         );
  NOR2X2 U23931 ( .A(BOPA[32]), .B(BOPA[30]), .Y(n8355) );
  NOR2X4 U23932 ( .A(n14244), .B(n14243), .Y(n14397) );
  NAND2X1 U23933 ( .A(n22434), .B(n22443), .Y(n22445) );
  OAI21X1 U23934 ( .A0(n11316), .A1(n11323), .B0(n11317), .Y(n11301) );
  NAND2X1 U23935 ( .A(n7062), .B(AOPC[38]), .Y(n11323) );
  NAND2X1 U23936 ( .A(n22506), .B(n22510), .Y(n14046) );
  OAI21XL U23937 ( .A0(n22044), .A1(n22374), .B0(n22045), .Y(n13115) );
  OAI21X1 U23938 ( .A0(n18815), .A1(n18814), .B0(n18813), .Y(n18859) );
  NOR2XL U23939 ( .A(n18807), .B(n18814), .Y(n18856) );
  AOI21X1 U23940 ( .A0(n9507), .A1(n9506), .B0(n9505), .Y(n9508) );
  OAI21XL U23941 ( .A0(n19332), .A1(n19303), .B0(n19302), .Y(n19313) );
  NOR2X1 U23942 ( .A(n14643), .B(n14642), .Y(n14696) );
  NAND2XL U23943 ( .A(n26347), .B(n26353), .Y(n26593) );
  AOI21X1 U23944 ( .A0(n26353), .A1(n26352), .B0(n26351), .Y(n26602) );
  AOI21X1 U23945 ( .A0(n9697), .A1(n9696), .B0(n9695), .Y(n9698) );
  NOR2X2 U23946 ( .A(n11168), .B(n11163), .Y(n11155) );
  OAI21XL U23947 ( .A0(n17257), .A1(n17234), .B0(n17233), .Y(n17240) );
  XNOR2X1 U23948 ( .A(n17332), .B(n17331), .Y(n17333) );
  AOI21X1 U23949 ( .A0(n11372), .A1(n11351), .B0(n11350), .Y(n11361) );
  XNOR2X2 U23950 ( .A(n10719), .B(n10718), .Y(U1_U2_z0[23]) );
  XNOR2X4 U23951 ( .A(n8281), .B(n8280), .Y(U1_U0_z0[15]) );
  AOI21X1 U23952 ( .A0(n24781), .A1(n25051), .B0(n9008), .Y(n9009) );
  AOI21X1 U23953 ( .A0(n19631), .A1(n19629), .B0(n19543), .Y(n19617) );
  ADDHX2 U23954 ( .A(U2_U0_y1[27]), .B(U2_U0_y0[27]), .CO(n26515), .S(n26461)
         );
  NAND2X1 U23955 ( .A(n9992), .B(n9995), .Y(n9998) );
  NOR2X1 U23956 ( .A(n8095), .B(AOPB[48]), .Y(n10359) );
  OAI21XL U23957 ( .A0(n19472), .A1(n19452), .B0(n19451), .Y(n19458) );
  OAI21X2 U23958 ( .A0(n14351), .A1(n14355), .B0(n14352), .Y(n14367) );
  ADDHX2 U23959 ( .A(U1_U0_y2[23]), .B(U1_U0_y0[23]), .CO(n8424), .S(n8421) );
  NAND2X1 U23960 ( .A(n25552), .B(n25510), .Y(n25512) );
  XNOR2X4 U23961 ( .A(n10380), .B(n10379), .Y(U0_U0_z0[21]) );
  CMPR22X1 U23962 ( .A(U0_U1_y2[15]), .B(U0_U1_y0[15]), .CO(n12457), .S(n12454) );
  NOR2X2 U23963 ( .A(n26762), .B(n26761), .Y(n26817) );
  INVXL U23964 ( .A(n11584), .Y(n8314) );
  OAI21XL U23965 ( .A0(n22745), .A1(n14155), .B0(n14154), .Y(n14156) );
  NAND2X1 U23966 ( .A(n8185), .B(BOPC[38]), .Y(n11142) );
  NAND2X1 U23967 ( .A(n19103), .B(n9709), .Y(n9711) );
  NAND2X1 U23968 ( .A(W2[12]), .B(W2[28]), .Y(n9942) );
  AOI21X1 U23969 ( .A0(n14117), .A1(n14116), .B0(n14115), .Y(n14118) );
  OAI21XL U23970 ( .A0(n19344), .A1(n19350), .B0(n19345), .Y(n19335) );
  NAND2X1 U23971 ( .A(n24661), .B(n24660), .Y(n24748) );
  AND2X2 U23972 ( .A(n9512), .B(U1_A_r_d0[19]), .Y(n19106) );
  XNOR2X2 U23973 ( .A(n11059), .B(n11058), .Y(U1_U1_z0[23]) );
  AOI21X1 U23974 ( .A0(n20230), .A1(n20214), .B0(n20213), .Y(n20221) );
  INVX1 U23975 ( .A(n20225), .Y(n20230) );
  CMPR22X1 U23976 ( .A(U2_U0_y1[35]), .B(U2_U0_y0[35]), .CO(n26948), .S(n26909) );
  INVXL U23977 ( .A(n11196), .Y(n11206) );
  XNOR2X1 U23978 ( .A(n17630), .B(n17629), .Y(n17631) );
  NAND2X2 U23979 ( .A(n11447), .B(n11513), .Y(n11449) );
  OAI21X1 U23980 ( .A0(n20069), .A1(n20058), .B0(n20057), .Y(n20067) );
  NAND2X1 U23981 ( .A(n24451), .B(n13464), .Y(n13466) );
  NAND2X2 U23982 ( .A(n9822), .B(n9821), .Y(n10173) );
  OAI21X1 U23983 ( .A0(n9699), .A1(n19128), .B0(n9698), .Y(n19102) );
  NAND2X1 U23984 ( .A(n13702), .B(U1_A_r_d0[19]), .Y(n19414) );
  CMPR22X1 U23985 ( .A(U0_U1_y2[35]), .B(U0_U1_y0[35]), .CO(n13157), .S(n13142) );
  NAND2X2 U23986 ( .A(n6989), .B(n11545), .Y(n11433) );
  NAND2X2 U23987 ( .A(n9970), .B(n9969), .Y(n10234) );
  OAI21XL U23988 ( .A0(n24422), .A1(n13491), .B0(n13490), .Y(n13492) );
  AOI21X1 U23989 ( .A0(n24431), .A1(n13489), .B0(n13488), .Y(n24422) );
  NAND2X2 U23990 ( .A(U2_B_r[6]), .B(n9626), .Y(n11579) );
  INVX2 U23991 ( .A(U2_B_i[6]), .Y(n9626) );
  INVXL U23992 ( .A(n10501), .Y(n10511) );
  NOR2X2 U23993 ( .A(n7060), .B(BOPC[39]), .Y(n11134) );
  OAI21X1 U23994 ( .A0(n22946), .A1(n23027), .B0(n22945), .Y(n23000) );
  AOI21X1 U23995 ( .A0(n6984), .A1(n24766), .B0(n24651), .Y(n24753) );
  OAI21X2 U23996 ( .A0(n10502), .A1(n10508), .B0(n10503), .Y(n8211) );
  OAI21X1 U23997 ( .A0(n10997), .A1(n10948), .B0(n10947), .Y(n10953) );
  NAND2X1 U23998 ( .A(n19557), .B(n14507), .Y(n17622) );
  OAI21X1 U23999 ( .A0(n22952), .A1(n23002), .B0(n22951), .Y(n22953) );
  NAND2X1 U24000 ( .A(n23006), .B(n23010), .Y(n22952) );
  AOI21X1 U24001 ( .A0(n23006), .A1(n23004), .B0(n22950), .Y(n22951) );
  AOI21X1 U24002 ( .A0(n22030), .A1(n22364), .B0(n13118), .Y(n13119) );
  AOI21X1 U24003 ( .A0(n17524), .A1(n17478), .B0(n17477), .Y(n17491) );
  XNOR2X4 U24004 ( .A(n10753), .B(n10752), .Y(U1_U2_z0[18]) );
  AOI21X1 U24005 ( .A0(n18251), .A1(n18250), .B0(n18249), .Y(n18492) );
  NAND2X1 U24006 ( .A(n8950), .B(n8949), .Y(n8968) );
  NOR2X1 U24007 ( .A(n8747), .B(n8746), .Y(n8821) );
  ADDHX2 U24008 ( .A(U0_U2_y1[18]), .B(U0_U2_y0[18]), .CO(n8747), .S(n8744) );
  AOI21X1 U24009 ( .A0(n8233), .A1(n10357), .B0(n8232), .Y(n8234) );
  ADDHX2 U24010 ( .A(U1_U1_y1[21]), .B(U1_U1_y0[21]), .CO(n14649), .S(n14646)
         );
  OAI21X2 U24011 ( .A0(n10456), .A1(n10465), .B0(n10457), .Y(n8217) );
  NAND2X2 U24012 ( .A(n8205), .B(AOPB[36]), .Y(n10465) );
  NOR2X2 U24013 ( .A(n8124), .B(BOPC[32]), .Y(n11181) );
  OAI21X2 U24014 ( .A0(n10524), .A1(n10527), .B0(n10525), .Y(n10501) );
  NOR2X1 U24015 ( .A(n9717), .B(U1_A_i_d0[24]), .Y(n9541) );
  NAND2X2 U24016 ( .A(n8064), .B(AOPB[34]), .Y(n10475) );
  NOR2X1 U24017 ( .A(n14538), .B(n22040), .Y(n14541) );
  XNOR2X4 U24018 ( .A(n10604), .B(n10603), .Y(U1_U0_z0[14]) );
  OAI21X2 U24019 ( .A0(n10965), .A1(n8324), .B0(n8323), .Y(n8325) );
  ADDHX2 U24020 ( .A(U1_U0_y2[28]), .B(U1_U0_y0[28]), .CO(n8435), .S(n8432) );
  OAI21XL U24021 ( .A0(n22440), .A1(n22439), .B0(n22438), .Y(n22441) );
  NAND2X1 U24022 ( .A(n9814), .B(n9825), .Y(n9864) );
  OAI21X1 U24023 ( .A0(n11321), .A1(n8340), .B0(n8339), .Y(n8341) );
  CMPR22X1 U24024 ( .A(U2_U0_y2[19]), .B(U2_U0_y0[19]), .CO(n23428), .S(n23366) );
  OAI21X1 U24025 ( .A0(n10446), .A1(n8222), .B0(n8221), .Y(n8223) );
  CMPR22X1 U24026 ( .A(U1_U0_y1[37]), .B(U1_U0_y0[37]), .CO(n9343), .S(n9339)
         );
  AOI21X1 U24027 ( .A0(n14958), .A1(n16824), .B0(n8051), .Y(n16810) );
  OAI21X1 U24028 ( .A0(n12529), .A1(n22687), .B0(n7042), .Y(n22657) );
  AND2XL U24029 ( .A(U0_U0_y1[0]), .B(U0_U0_y0[0]), .Y(n7958) );
  AND2X1 U24030 ( .A(n14961), .B(n20041), .Y(n7960) );
  OR2X2 U24031 ( .A(n14564), .B(n24640), .Y(n7963) );
  AND2X2 U24032 ( .A(n24685), .B(n24684), .Y(n7966) );
  OR2X2 U24033 ( .A(n5797), .B(n19243), .Y(n7969) );
  OR2X2 U24034 ( .A(n24634), .B(n24633), .Y(n7999) );
  XNOR2X1 U24035 ( .A(n14992), .B(n14991), .Y(n8044) );
  AND2X2 U24036 ( .A(n5855), .B(n14957), .Y(n8051) );
  AND2X2 U24037 ( .A(n17297), .B(n17296), .Y(n8052) );
  OR2X2 U24038 ( .A(n25199), .B(U2_A_i_d[14]), .Y(n8057) );
  OR2X2 U24039 ( .A(n21774), .B(U2_A_i_d[14]), .Y(n8058) );
  OR2X2 U24040 ( .A(n14133), .B(U2_A_r_d[20]), .Y(n8078) );
  NOR2X1 U24041 ( .A(n8063), .B(AOPD[34]), .Y(n10994) );
  OR2X2 U24042 ( .A(n14575), .B(n24676), .Y(n8083) );
  OR2X2 U24043 ( .A(n8451), .B(n8450), .Y(n8149) );
  AND2XL U24044 ( .A(U1_U2_y1[0]), .B(U1_U2_y0[0]), .Y(n12707) );
  AOI21X1 U24045 ( .A0(n8338), .A1(n11301), .B0(n8337), .Y(n8339) );
  AOI21XL U24046 ( .A0(n12029), .A1(n12028), .B0(n12027), .Y(n12030) );
  AOI21XL U24047 ( .A0(n9248), .A1(n9247), .B0(n9246), .Y(n9249) );
  AOI21XL U24048 ( .A0(n9281), .A1(n9280), .B0(n9279), .Y(n9282) );
  CMPR22X1 U24049 ( .A(U0_U2_y1[36]), .B(U0_U2_y0[36]), .CO(n9205), .S(n9191)
         );
  ADDHX2 U24050 ( .A(U0_U1_y2[20]), .B(U0_U1_y0[20]), .CO(n12478), .S(n12466)
         );
  OR2X2 U24051 ( .A(n13235), .B(U0_U0_y0[13]), .Y(n13238) );
  AOI21XL U24052 ( .A0(n5779), .A1(n8787), .B0(n8786), .Y(n8788) );
  NOR2X1 U24053 ( .A(n11451), .B(U2_B_r[21]), .Y(n11497) );
  OAI21X1 U24054 ( .A0(n11389), .A1(n11262), .B0(n11261), .Y(n11266) );
  INVX8 U24055 ( .A(n8242), .Y(n11428) );
  OR2X2 U24056 ( .A(n8791), .B(U0_U1_y0[13]), .Y(n8794) );
  OAI21X1 U24057 ( .A0(n13081), .A1(n13080), .B0(n13079), .Y(n13583) );
  ADDHX2 U24058 ( .A(U2_U0_y1[30]), .B(U2_U0_y0[30]), .CO(n26702), .S(n26646)
         );
  INVX1 U24059 ( .A(n23525), .Y(n18143) );
  AOI21XL U24060 ( .A0(n12495), .A1(n12494), .B0(n12493), .Y(n12496) );
  AOI21XL U24061 ( .A0(n14719), .A1(n14718), .B0(n14717), .Y(n14720) );
  AOI21XL U24062 ( .A0(n26056), .A1(n26055), .B0(n26054), .Y(n26057) );
  AOI21XL U24063 ( .A0(n21298), .A1(n21328), .B0(n21327), .Y(n21383) );
  AOI21XL U24064 ( .A0(n18640), .A1(n18565), .B0(n18639), .Y(n18670) );
  NOR2X1 U24065 ( .A(n26406), .B(n26405), .Y(n26456) );
  AOI21XL U24066 ( .A0(n19054), .A1(n19053), .B0(n19052), .Y(n19061) );
  AND2X1 U24067 ( .A(n14150), .B(U2_A_r_d[23]), .Y(n13488) );
  OAI21XL U24068 ( .A0(n22081), .A1(n22079), .B0(n22082), .Y(n14523) );
  NAND2X1 U24069 ( .A(n14132), .B(n14140), .Y(n14143) );
  AND2X1 U24070 ( .A(n19775), .B(U1_A_i_d0[23]), .Y(n8685) );
  XOR2XL U24071 ( .A(U1_U2_y0[40]), .B(U1_U2_y2[40]), .Y(n13993) );
  XNOR2X1 U24072 ( .A(n12934), .B(n12933), .Y(n19330) );
  AOI21X1 U24073 ( .A0(n9602), .A1(n17191), .B0(n9601), .Y(n17181) );
  AOI21XL U24074 ( .A0(n23255), .A1(n23254), .B0(n23253), .Y(n23458) );
  AOI21XL U24075 ( .A0(n26770), .A1(n26714), .B0(n26769), .Y(n26771) );
  AOI21XL U24076 ( .A0(n26537), .A1(n26536), .B0(n26535), .Y(n26773) );
  AOI21X1 U24077 ( .A0(n21571), .A1(n5765), .B0(n21570), .Y(n21572) );
  AOI21X1 U24078 ( .A0(n22236), .A1(n22200), .B0(n22199), .Y(n22212) );
  OR2X2 U24079 ( .A(n24632), .B(n24631), .Y(n24779) );
  INVX1 U24080 ( .A(n25173), .Y(n25503) );
  OR2X2 U24081 ( .A(n12378), .B(n22918), .Y(n22028) );
  AOI21X1 U24082 ( .A0(n21879), .A1(n21841), .B0(n21840), .Y(n21851) );
  AOI21X1 U24083 ( .A0(n12170), .A1(n12169), .B0(n12168), .Y(n25724) );
  AOI21XL U24084 ( .A0(n13884), .A1(n13883), .B0(n13882), .Y(n17108) );
  AOI21XL U24085 ( .A0(n12850), .A1(n12849), .B0(n12848), .Y(n12855) );
  AOI21XL U24086 ( .A0(OP2_done0), .A1(Q3[1]), .B0(n27820), .Y(n28289) );
  AOI21XL U24087 ( .A0(B4_q[30]), .A1(n5925), .B0(n5924), .Y(n15857) );
  AOI21XL U24088 ( .A0(B2_q[10]), .A1(n15958), .B0(n5924), .Y(n15183) );
  AOI21XL U24089 ( .A0(B0_q[32]), .A1(n15557), .B0(n16051), .Y(n16052) );
  AOI21XL U24090 ( .A0(B0_q[41]), .A1(n15687), .B0(n28985), .Y(n16203) );
  AOI21XL U24091 ( .A0(B3_q[42]), .A1(n7127), .B0(n5924), .Y(n16397) );
  AOI21XL U24092 ( .A0(B0_q[9]), .A1(n5925), .B0(n5924), .Y(n15187) );
  AOI21XL U24093 ( .A0(n26735), .A1(n26791), .B0(n26794), .Y(n26740) );
  AOI21XL U24094 ( .A0(n25961), .A1(n25907), .B0(n25906), .Y(n25912) );
  AOI21XL U24095 ( .A0(n23313), .A1(n23233), .B0(n23232), .Y(n23238) );
  AOI21XL U24096 ( .A0(n26924), .A1(n26883), .B0(n26923), .Y(n26980) );
  AOI21XL U24097 ( .A0(n23665), .A1(n23664), .B0(n23663), .Y(n23670) );
  AOI21XL U24098 ( .A0(n24051), .A1(n23893), .B0(n23991), .Y(n23947) );
  AOI21XL U24099 ( .A0(n26829), .A1(n26774), .B0(n26828), .Y(n26874) );
  AOI21XL U24100 ( .A0(n26014), .A1(n26111), .B0(n26116), .Y(n26065) );
  AOI21XL U24101 ( .A0(n24364), .A1(n24322), .B0(n24363), .Y(n24390) );
  AOI21XL U24102 ( .A0(n23534), .A1(n23533), .B0(n23532), .Y(n23539) );
  AOI21XL U24103 ( .A0(B4_q[0]), .A1(n5925), .B0(n5924), .Y(n15983) );
  AOI21XL U24104 ( .A0(B4_q[13]), .A1(n15969), .B0(n16496), .Y(n15925) );
  AOI21XL U24105 ( .A0(B6_q[20]), .A1(n15958), .B0(n5924), .Y(n15897) );
  AOI21XL U24106 ( .A0(B5_q[25]), .A1(n16165), .B0(n5924), .Y(n15482) );
  AOI21XL U24107 ( .A0(n18274), .A1(n18273), .B0(n18272), .Y(n18279) );
  AOI21XL U24108 ( .A0(n20185), .A1(n20184), .B0(n20183), .Y(n20491) );
  AOI21XL U24109 ( .A0(n21582), .A1(n21539), .B0(n21581), .Y(n21624) );
  AOI21XL U24110 ( .A0(n18660), .A1(n18716), .B0(n18719), .Y(n18665) );
  XOR2XL U24111 ( .A(n28988), .B(U1_pipe15[27]), .Y(n18993) );
  AOI21XL U24112 ( .A0(n18388), .A1(n18387), .B0(n18386), .Y(n18393) );
  AOI21XL U24113 ( .A0(n21686), .A1(n21649), .B0(n21685), .Y(n21725) );
  AOI21XL U24114 ( .A0(n20623), .A1(n20711), .B0(n20716), .Y(n20667) );
  AOI21XL U24115 ( .A0(n21015), .A1(n21014), .B0(n21013), .Y(n21022) );
  OAI21XL U24116 ( .A0(n25070), .A1(n25059), .B0(n25058), .Y(n25067) );
  AOI21XL U24117 ( .A0(n25218), .A1(n25211), .B0(n25210), .Y(n25214) );
  OAI21XL U24118 ( .A0(n23081), .A1(n23065), .B0(n23064), .Y(n23077) );
  AOI21XL U24119 ( .A0(n25422), .A1(n25420), .B0(n25412), .Y(n25417) );
  OAI21XL U24120 ( .A0(n17697), .A1(n17681), .B0(n17680), .Y(n17693) );
  OAI21XL U24121 ( .A0(n16887), .A1(n16870), .B0(n16869), .Y(n16883) );
  OAI21XL U24122 ( .A0(n19184), .A1(n19154), .B0(n19153), .Y(n19164) );
  AOI21XL U24123 ( .A0(n19313), .A1(n19304), .B0(n8146), .Y(n19308) );
  AOI21XL U24124 ( .A0(n7685), .A1(n19444), .B0(n19443), .Y(n19446) );
  OAI21XL U24125 ( .A0(n28981), .A1(n27976), .B0(n27265), .Y(n27793) );
  AOI21XL U24126 ( .A0(n11885), .A1(n11999), .B0(n28637), .Y(n11883) );
  AOI21XL U24127 ( .A0(n15982), .A1(B3_q[47]), .B0(n15056), .Y(n15058) );
  XNOR2XL U24128 ( .A(n26845), .B(n26801), .Y(n26802) );
  XOR2XL U24129 ( .A(n26003), .B(n25965), .Y(n25966) );
  XOR2XL U24130 ( .A(n24858), .B(n25808), .Y(n24859) );
  XOR2XL U24131 ( .A(n23661), .B(n23660), .Y(n23662) );
  XOR2XL U24132 ( .A(n26980), .B(n26928), .Y(n26929) );
  XOR2XL U24133 ( .A(n26341), .B(n26102), .Y(n26103) );
  XOR2XL U24134 ( .A(n24078), .B(n24077), .Y(n24079) );
  XOR2XL U24135 ( .A(n23247), .B(n23246), .Y(n23248) );
  XNOR2XL U24136 ( .A(n24051), .B(n23896), .Y(n23897) );
  XOR2XL U24137 ( .A(n22733), .B(n23153), .Y(n22734) );
  XOR2XL U24138 ( .A(n26417), .B(n26309), .Y(n26310) );
  XOR2XL U24139 ( .A(n25455), .B(n25823), .Y(n25456) );
  XNOR2XL U24140 ( .A(n24062), .B(n23865), .Y(n23866) );
  XOR2XL U24141 ( .A(n23266), .B(n23265), .Y(n23267) );
  XOR2XL U24142 ( .A(n26696), .B(n26695), .Y(n26697) );
  XOR2XL U24143 ( .A(n21389), .B(n21388), .Y(n21390) );
  XNOR2XL U24144 ( .A(n18090), .B(n18089), .Y(n18091) );
  XOR2XL U24145 ( .A(n18937), .B(n18901), .Y(n18902) );
  XOR2XL U24146 ( .A(n21082), .B(n20976), .Y(n20977) );
  XOR2XL U24147 ( .A(n17452), .B(n17774), .Y(n17453) );
  XNOR2XL U24148 ( .A(n18660), .B(n18518), .Y(n18519) );
  XOR2XL U24149 ( .A(n17864), .B(n17863), .Y(n17865) );
  XOR2XL U24150 ( .A(n18687), .B(n18686), .Y(n18688) );
  XOR2XL U24151 ( .A(n20986), .B(n20772), .Y(n20773) );
  XOR2XL U24152 ( .A(n21648), .B(n21594), .Y(n21595) );
  XNOR2XL U24153 ( .A(n18178), .B(n18134), .Y(n18135) );
  XOR2XL U24154 ( .A(n18834), .B(n18804), .Y(n18805) );
  XNOR2XL U24155 ( .A(n20824), .B(n20823), .Y(n20825) );
  XOR2XL U24156 ( .A(n21049), .B(n20930), .Y(n20931) );
  XOR2XL U24157 ( .A(n24924), .B(n24923), .Y(n24925) );
  XNOR2XL U24158 ( .A(n22413), .B(n22412), .Y(n22414) );
  XOR2XL U24159 ( .A(n22228), .B(n22227), .Y(n22229) );
  XOR2XL U24160 ( .A(n24823), .B(n24822), .Y(n24824) );
  XNOR2XL U24161 ( .A(n24556), .B(n24555), .Y(n24557) );
  XOR2XL U24162 ( .A(n25617), .B(n25616), .Y(n25618) );
  XNOR2XL U24163 ( .A(n22085), .B(n22084), .Y(n22086) );
  XOR2XL U24164 ( .A(n21936), .B(n21935), .Y(n21937) );
  XNOR2XL U24165 ( .A(n25258), .B(n25257), .Y(n25259) );
  XOR2XL U24166 ( .A(n23113), .B(n23112), .Y(n23114) );
  XOR2XL U24167 ( .A(n25718), .B(n25717), .Y(n25719) );
  XOR2XL U24168 ( .A(n22527), .B(n22812), .Y(n22528) );
  XNOR2XL U24169 ( .A(n20163), .B(n20162), .Y(n20164) );
  XOR2XL U24170 ( .A(n17248), .B(n17545), .Y(n17250) );
  XNOR2XL U24171 ( .A(n20447), .B(n20446), .Y(n20448) );
  XOR2XL U24172 ( .A(n17570), .B(n17569), .Y(n17571) );
  XNOR2XL U24173 ( .A(n17115), .B(n17114), .Y(n17116) );
  XNOR2XL U24174 ( .A(n19487), .B(n19486), .Y(n19488) );
  XOR2XL U24175 ( .A(n19662), .B(n19661), .Y(n19663) );
  AOI21XL U24176 ( .A0(n11993), .A1(n11992), .B0(n11994), .Y(A7_CEN) );
  AOI21XL U24177 ( .A0(n11993), .A1(n11645), .B0(n11994), .Y(A6_CEN) );
  AOI21XL U24178 ( .A0(n11992), .A1(n11646), .B0(n11994), .Y(A5_CEN) );
  AOI21XL U24179 ( .A0(n11993), .A1(n11992), .B0(n29241), .Y(A3_CEN) );
  AOI21XL U24180 ( .A0(n11993), .A1(n11645), .B0(n29241), .Y(A2_CEN) );
  AOI21XL U24181 ( .A0(n11992), .A1(n11646), .B0(n29241), .Y(A1_CEN) );
  NOR2X1 U24182 ( .A(n8075), .B(AOPD[30]), .Y(n11003) );
  NAND2X1 U24183 ( .A(n8075), .B(AOPD[30]), .Y(n11010) );
  INVXL U24184 ( .A(n8318), .Y(n8209) );
  NOR2X2 U24185 ( .A(n8208), .B(AOPB[26]), .Y(n10527) );
  NAND2X1 U24186 ( .A(n8081), .B(AOPB[29]), .Y(n10503) );
  AOI21X4 U24187 ( .A0(n8212), .A1(n10501), .B0(n8211), .Y(n10478) );
  NAND2X1 U24188 ( .A(n8076), .B(AOPB[30]), .Y(n10497) );
  OAI21X2 U24189 ( .A0(n10492), .A1(n10497), .B0(n10493), .Y(n10479) );
  AOI21X2 U24190 ( .A0(n8214), .A1(n10479), .B0(n8213), .Y(n8215) );
  OAI21X4 U24191 ( .A0(n8216), .A1(n10478), .B0(n8215), .Y(n10414) );
  NOR2X2 U24192 ( .A(n7990), .B(AOPB[40]), .Y(n10430) );
  NOR2X1 U24193 ( .A(n8197), .B(AOPB[41]), .Y(n10421) );
  NOR2X1 U24194 ( .A(n10430), .B(n10421), .Y(n8220) );
  NAND2X1 U24195 ( .A(n10427), .B(n8220), .Y(n8222) );
  NOR2X1 U24196 ( .A(n8064), .B(AOPB[34]), .Y(n10474) );
  NOR2X2 U24197 ( .A(n8061), .B(AOPB[35]), .Y(n10469) );
  NOR2X2 U24198 ( .A(n8205), .B(AOPB[36]), .Y(n10452) );
  NAND2X1 U24199 ( .A(n8061), .B(AOPB[35]), .Y(n10470) );
  AOI21X4 U24200 ( .A0(n8218), .A1(n10462), .B0(n8217), .Y(n10446) );
  NAND2XL U24201 ( .A(n8197), .B(AOPB[41]), .Y(n10422) );
  OAI21XL U24202 ( .A0(n10421), .A1(n10431), .B0(n10422), .Y(n8219) );
  AOI21X4 U24203 ( .A0(n10414), .A1(n8224), .B0(n8223), .Y(n10413) );
  BUFX12 U24204 ( .A(n10413), .Y(n10522) );
  NOR2X1 U24205 ( .A(n7057), .B(AOPB[42]), .Y(n10409) );
  NOR2XL U24206 ( .A(n10409), .B(n10404), .Y(n10396) );
  NAND2X1 U24207 ( .A(n10396), .B(n8226), .Y(n10382) );
  INVXL U24208 ( .A(n10382), .Y(n10371) );
  NAND2XL U24209 ( .A(n8110), .B(AOPB[44]), .Y(n10400) );
  NAND2XL U24210 ( .A(n8108), .B(AOPB[45]), .Y(n10392) );
  OAI21XL U24211 ( .A0(n10391), .A1(n10400), .B0(n10392), .Y(n8225) );
  NAND2XL U24212 ( .A(n8098), .B(AOPB[47]), .Y(n10377) );
  NAND2XL U24213 ( .A(n8095), .B(AOPB[48]), .Y(n10358) );
  NAND2X1 U24214 ( .A(n8229), .B(n10358), .Y(n8230) );
  XNOR2X4 U24215 ( .A(n8231), .B(n8230), .Y(U0_U0_z0[22]) );
  NOR2XL U24216 ( .A(n10359), .B(n10365), .Y(n8233) );
  NOR2X1 U24217 ( .A(n10382), .B(n8235), .Y(n10513) );
  INVXL U24218 ( .A(n10513), .Y(n8237) );
  NAND2XL U24219 ( .A(n8092), .B(AOPB[49]), .Y(n10366) );
  OAI21XL U24220 ( .A0(n10365), .A1(n10358), .B0(n10366), .Y(n8232) );
  OAI21X2 U24221 ( .A0(n10522), .A1(n8237), .B0(n8236), .Y(n8239) );
  NAND2X1 U24222 ( .A(n10349), .B(n10515), .Y(n8238) );
  XNOR2X4 U24223 ( .A(n8239), .B(n8238), .Y(U0_U0_z0[24]) );
  NOR2X4 U24224 ( .A(BOPA[29]), .B(BOPA[27]), .Y(n8354) );
  NOR2X2 U24225 ( .A(BOPA[33]), .B(BOPA[31]), .Y(n8240) );
  INVX8 U24226 ( .A(n11428), .Y(n11427) );
  INVX8 U24227 ( .A(n8242), .Y(n11430) );
  NAND2XL U24228 ( .A(BOPA[11]), .B(n11430), .Y(n8243) );
  OAI21XL U24229 ( .A0(n28747), .A1(n11430), .B0(n8243), .Y(U2_B_r[11]) );
  NOR2X1 U24230 ( .A(n8268), .B(BOPA[36]), .Y(n8244) );
  CLKINVX4 U24231 ( .A(U2_factor_reg), .Y(n11418) );
  XNOR2X1 U24232 ( .A(n8247), .B(BOPA[43]), .Y(n8249) );
  NAND2X2 U24233 ( .A(n8139), .B(BOPD[28]), .Y(n10862) );
  NOR2X1 U24234 ( .A(n8134), .B(BOPD[30]), .Y(n10830) );
  NOR2X1 U24235 ( .A(n10830), .B(n10832), .Y(n10819) );
  NOR2X2 U24236 ( .A(n8118), .B(BOPD[35]), .Y(n10808) );
  NOR2X1 U24237 ( .A(n10813), .B(n10808), .Y(n10803) );
  NOR2X1 U24238 ( .A(n8192), .B(BOPD[36]), .Y(n10794) );
  NOR2X2 U24239 ( .A(n8189), .B(BOPD[37]), .Y(n10798) );
  NOR2X2 U24240 ( .A(n10794), .B(n10798), .Y(n8253) );
  NAND2X1 U24241 ( .A(n10803), .B(n8253), .Y(n10790) );
  OAI21X2 U24242 ( .A0(n10808), .A1(n10814), .B0(n10809), .Y(n10804) );
  NAND2XL U24243 ( .A(n8189), .B(BOPD[37]), .Y(n10799) );
  OAI21X1 U24244 ( .A0(n10798), .A1(n10805), .B0(n10799), .Y(n8252) );
  AOI21X4 U24245 ( .A0(n8253), .A1(n10804), .B0(n8252), .Y(n10789) );
  NAND2XL U24246 ( .A(n7058), .B(BOPD[41]), .Y(n10769) );
  NOR2X1 U24247 ( .A(n8172), .B(BOPD[44]), .Y(n10737) );
  NOR2X1 U24248 ( .A(n8170), .B(BOPD[45]), .Y(n10741) );
  NOR2X1 U24249 ( .A(n10737), .B(n10741), .Y(n8258) );
  NAND2XL U24250 ( .A(n10746), .B(n8258), .Y(n10732) );
  INVXL U24251 ( .A(n10732), .Y(n10720) );
  NOR2XL U24252 ( .A(n8165), .B(BOPD[46]), .Y(n10691) );
  NAND2XL U24253 ( .A(n10720), .B(n10734), .Y(n8261) );
  NAND2XL U24254 ( .A(n8170), .B(BOPD[45]), .Y(n10742) );
  INVXL U24255 ( .A(n10731), .Y(n10723) );
  NAND2XL U24256 ( .A(n8165), .B(BOPD[46]), .Y(n10733) );
  INVXL U24257 ( .A(n10733), .Y(n8259) );
  AOI21XL U24258 ( .A0(n10723), .A1(n10734), .B0(n8259), .Y(n8260) );
  INVXL U24259 ( .A(n10693), .Y(n8262) );
  NAND2XL U24260 ( .A(n8162), .B(BOPD[47]), .Y(n10692) );
  NAND2X1 U24261 ( .A(n8262), .B(n10692), .Y(n8263) );
  NAND2XL U24262 ( .A(n11633), .B(n11979), .Y(n28638) );
  OAI21XL U24263 ( .A0(cnt[0]), .A1(cnt[2]), .B0(n11963), .Y(n8265) );
  AOI22XL U24264 ( .A0(n11878), .A1(cnt[2]), .B0(cnt[0]), .B1(n29107), .Y(
        n8266) );
  AOI22XL U24265 ( .A0(n7305), .A1(n28704), .B0(n8266), .B1(n11633), .Y(n28636) );
  AOI21XL U24266 ( .A0(n11885), .A1(n15024), .B0(n28636), .Y(n8267) );
  NAND2X1 U24267 ( .A(n11418), .B(BOPA[10]), .Y(n8269) );
  NOR2X1 U24268 ( .A(n8184), .B(BOPB[38]), .Y(n10605) );
  NOR2X2 U24269 ( .A(n8183), .B(BOPB[39]), .Y(n10611) );
  NOR2X2 U24270 ( .A(n10605), .B(n10611), .Y(n10597) );
  INVXL U24271 ( .A(n10597), .Y(n8271) );
  NOR2XL U24272 ( .A(n8271), .B(n10600), .Y(n8276) );
  NAND2X1 U24273 ( .A(n8184), .B(BOPB[38]), .Y(n10618) );
  NAND2XL U24274 ( .A(n8183), .B(BOPB[39]), .Y(n10612) );
  OAI21X1 U24275 ( .A0(n10611), .A1(n10618), .B0(n10612), .Y(n10596) );
  INVXL U24276 ( .A(n10596), .Y(n8274) );
  NAND2X1 U24277 ( .A(n6944), .B(BOPB[40]), .Y(n10601) );
  OAI21XL U24278 ( .A0(n8274), .A1(n10600), .B0(n10601), .Y(n8275) );
  NOR2X2 U24279 ( .A(n8179), .B(BOPB[41]), .Y(n9555) );
  INVXL U24280 ( .A(n9555), .Y(n8279) );
  NAND2X1 U24281 ( .A(n8279), .B(n9554), .Y(n8280) );
  NAND2X1 U24282 ( .A(n8167), .B(BOPC[27]), .Y(n11219) );
  NOR2X1 U24283 ( .A(n8133), .B(BOPC[30]), .Y(n11185) );
  NAND2XL U24284 ( .A(n8282), .B(BOPC[33]), .Y(n11177) );
  NOR2X1 U24285 ( .A(n8120), .B(BOPC[34]), .Y(n11168) );
  NAND2X1 U24286 ( .A(n8181), .B(BOPC[40]), .Y(n11124) );
  OAI21XL U24287 ( .A0(n11114), .A1(n11124), .B0(n11115), .Y(n8285) );
  AOI21XL U24288 ( .A0(n8286), .A1(n11119), .B0(n8285), .Y(n8287) );
  NOR2XL U24289 ( .A(n8164), .B(BOPC[46]), .Y(n11069) );
  NOR2XL U24290 ( .A(n11069), .B(n11075), .Y(n11061) );
  NOR2XL U24291 ( .A(n11064), .B(n11055), .Y(n8292) );
  NAND2XL U24292 ( .A(n11061), .B(n8292), .Y(n8294) );
  INVXL U24293 ( .A(n11208), .Y(n8296) );
  NAND2XL U24294 ( .A(n7061), .B(BOPC[45]), .Y(n11088) );
  NAND2XL U24295 ( .A(n8164), .B(BOPC[46]), .Y(n11081) );
  NAND2XL U24296 ( .A(n8161), .B(BOPC[47]), .Y(n11076) );
  OAI21XL U24297 ( .A0(n11075), .A1(n11081), .B0(n11076), .Y(n11060) );
  OAI21XL U24298 ( .A0(n11055), .A1(n11065), .B0(n11056), .Y(n8291) );
  AOI21XL U24299 ( .A0(n8292), .A1(n11060), .B0(n8291), .Y(n8293) );
  INVXL U24300 ( .A(n11214), .Y(n8295) );
  NAND2X1 U24301 ( .A(n11043), .B(n11210), .Y(n8297) );
  XNOR2X4 U24302 ( .A(n8298), .B(n8297), .Y(U1_U1_z0[24]) );
  NAND2XL U24303 ( .A(BOPA[4]), .B(n11430), .Y(n8299) );
  OAI21XL U24304 ( .A0(n29104), .A1(n11428), .B0(n8299), .Y(U2_B_r[4]) );
  NAND2X1 U24305 ( .A(n11418), .B(BOPA[1]), .Y(n8300) );
  MXI2X2 U24306 ( .A(n28751), .B(n28676), .S0(n11430), .Y(U2_B_r[0]) );
  NAND2XL U24307 ( .A(BOPA[3]), .B(n11430), .Y(n8303) );
  OAI21XL U24308 ( .A0(n29103), .A1(n11428), .B0(n8303), .Y(U2_B_r[3]) );
  NAND2XL U24309 ( .A(BOPA[2]), .B(n11430), .Y(n8306) );
  NOR2X4 U24310 ( .A(U2_B_r[0]), .B(n11603), .Y(n11601) );
  NAND2X1 U24311 ( .A(n8311), .B(U2_B_r[2]), .Y(n11596) );
  INVX1 U24312 ( .A(n11596), .Y(n11591) );
  INVXL U24313 ( .A(n11592), .Y(n8312) );
  NOR2X1 U24314 ( .A(n8313), .B(U2_B_r[4]), .Y(n11584) );
  NOR2X2 U24315 ( .A(n8324), .B(n10966), .Y(n8326) );
  NAND2X1 U24316 ( .A(n8199), .B(AOPD[38]), .Y(n10967) );
  NAND2XL U24317 ( .A(n7989), .B(AOPD[39]), .Y(n10961) );
  OAI21X1 U24318 ( .A0(n10960), .A1(n10967), .B0(n10961), .Y(n10945) );
  OAI21XL U24319 ( .A0(n10940), .A1(n10950), .B0(n10941), .Y(n8321) );
  AOI21X1 U24320 ( .A0(n8322), .A1(n10945), .B0(n8321), .Y(n8323) );
  NOR2X1 U24321 ( .A(n8115), .B(AOPD[42]), .Y(n10930) );
  NOR2X1 U24322 ( .A(n8107), .B(AOPD[45]), .Y(n10915) );
  NAND2XL U24323 ( .A(n10920), .B(n8328), .Y(n10906) );
  INVXL U24324 ( .A(n10906), .Y(n10894) );
  NAND2XL U24325 ( .A(n10894), .B(n10908), .Y(n8331) );
  NAND2X1 U24326 ( .A(n8115), .B(AOPD[42]), .Y(n10931) );
  OAI21X2 U24327 ( .A0(n10926), .A1(n10931), .B0(n10927), .Y(n10921) );
  NAND2XL U24328 ( .A(n6950), .B(AOPD[44]), .Y(n10924) );
  NAND2XL U24329 ( .A(n8107), .B(AOPD[45]), .Y(n10916) );
  OAI21XL U24330 ( .A0(n10915), .A1(n10924), .B0(n10916), .Y(n8327) );
  AOI21X2 U24331 ( .A0(n8328), .A1(n10921), .B0(n8327), .Y(n10905) );
  AOI21X1 U24332 ( .A0(n10897), .A1(n10908), .B0(n8329), .Y(n8330) );
  NAND2XL U24333 ( .A(n8097), .B(AOPD[47]), .Y(n10867) );
  NAND2X1 U24334 ( .A(n8332), .B(n10867), .Y(n8333) );
  XNOR2X4 U24335 ( .A(n8334), .B(n8333), .Y(U0_U2_z0[21]) );
  NAND2X1 U24336 ( .A(n8084), .B(AOPC[28]), .Y(n11392) );
  NAND2X1 U24337 ( .A(n8079), .B(AOPC[29]), .Y(n11375) );
  NOR2X2 U24338 ( .A(n8067), .B(AOPC[32]), .Y(n11357) );
  NOR2X2 U24339 ( .A(n8059), .B(AOPC[35]), .Y(n9646) );
  NOR2X1 U24340 ( .A(n11344), .B(n9646), .Y(n11336) );
  NOR2X1 U24341 ( .A(n11322), .B(n8340), .Y(n8342) );
  OAI21X2 U24342 ( .A0(n9646), .A1(n11345), .B0(n9647), .Y(n11337) );
  NAND2X1 U24343 ( .A(n8200), .B(AOPC[37]), .Y(n11332) );
  AOI21X2 U24344 ( .A0(n8336), .A1(n11337), .B0(n8335), .Y(n11321) );
  NAND2X1 U24345 ( .A(n7954), .B(AOPC[39]), .Y(n11317) );
  AOI21X2 U24346 ( .A0(n9645), .A1(n8342), .B0(n8341), .Y(n8343) );
  NOR2X1 U24347 ( .A(n8114), .B(AOPC[42]), .Y(n11288) );
  NOR2X1 U24348 ( .A(n8111), .B(AOPC[43]), .Y(n11284) );
  NOR2XL U24349 ( .A(n8109), .B(AOPC[44]), .Y(n11267) );
  NOR2X1 U24350 ( .A(n11267), .B(n11271), .Y(n8345) );
  INVXL U24351 ( .A(n11262), .Y(n11250) );
  NOR2XL U24352 ( .A(n8099), .B(AOPC[46]), .Y(n11222) );
  NAND2XL U24353 ( .A(n11250), .B(n11264), .Y(n8348) );
  NAND2XL U24354 ( .A(n8111), .B(AOPC[43]), .Y(n11285) );
  NAND2XL U24355 ( .A(n8109), .B(AOPC[44]), .Y(n11280) );
  NAND2XL U24356 ( .A(n8106), .B(AOPC[45]), .Y(n11272) );
  OAI21XL U24357 ( .A0(n11271), .A1(n11280), .B0(n11272), .Y(n8344) );
  NAND2XL U24358 ( .A(n8096), .B(AOPC[47]), .Y(n11223) );
  NAND2X1 U24359 ( .A(n8349), .B(n11223), .Y(n8350) );
  XNOR2X4 U24360 ( .A(n8351), .B(n8350), .Y(U0_U1_z0[21]) );
  NOR2X1 U24361 ( .A(W0[8]), .B(W0[24]), .Y(n9810) );
  INVXL U24362 ( .A(n9810), .Y(n9855) );
  NAND2X1 U24363 ( .A(W0[8]), .B(W0[24]), .Y(n9854) );
  INVXL U24364 ( .A(n9854), .Y(n8352) );
  NAND4X1 U24365 ( .A(n7031), .B(n8356), .C(n8355), .D(n29100), .Y(n8357) );
  XOR2X1 U24366 ( .A(n8357), .B(n6932), .Y(n8359) );
  NAND2XL U24367 ( .A(n11418), .B(BOPA[9]), .Y(n8358) );
  CMPR22X1 U24368 ( .A(U1_U0_y2[18]), .B(U1_U0_y0[18]), .CO(n8414), .S(n8411)
         );
  NOR2X1 U24369 ( .A(n8414), .B(n8413), .Y(n8468) );
  AND2XL U24370 ( .A(U1_U0_y2[0]), .B(U1_U0_y0[0]), .Y(n8361) );
  OR2X1 U24371 ( .A(U1_U0_y2[3]), .B(U1_U0_y0[3]), .Y(n8366) );
  NAND2XL U24372 ( .A(n8363), .B(n8366), .Y(n8368) );
  AOI21XL U24373 ( .A0(n8366), .A1(n8365), .B0(n8364), .Y(n8367) );
  OAI21XL U24374 ( .A0(n8369), .A1(n8368), .B0(n8367), .Y(n8384) );
  OR2X2 U24375 ( .A(U1_U0_y2[5]), .B(U1_U0_y0[5]), .Y(n8375) );
  OR2X2 U24376 ( .A(U1_U0_y2[6]), .B(U1_U0_y0[6]), .Y(n8372) );
  OR2X2 U24377 ( .A(U1_U0_y2[7]), .B(U1_U0_y0[7]), .Y(n8378) );
  AOI21X1 U24378 ( .A0(n8378), .A1(n8377), .B0(n8376), .Y(n8379) );
  OAI21XL U24379 ( .A0(n8381), .A1(n8380), .B0(n8379), .Y(n8382) );
  CMPR22X1 U24380 ( .A(U1_U0_y2[14]), .B(U1_U0_y0[14]), .CO(n8406), .S(n8400)
         );
  OR2X2 U24381 ( .A(U1_U0_y2[9]), .B(U1_U0_y0[9]), .Y(n8391) );
  OR2X2 U24382 ( .A(U1_U0_y2[10]), .B(U1_U0_y0[10]), .Y(n8387) );
  OR2X2 U24383 ( .A(U1_U0_y2[11]), .B(U1_U0_y0[11]), .Y(n8394) );
  OAI21XL U24384 ( .A0(n8397), .A1(n8396), .B0(n8395), .Y(n8494) );
  NAND2XL U24385 ( .A(n8400), .B(U1_U0_y2[13]), .Y(n8504) );
  OAI21XL U24386 ( .A0(n8499), .A1(n8503), .B0(n8504), .Y(n8401) );
  NAND2XL U24387 ( .A(n8408), .B(n8407), .Y(n8516) );
  ADDHX2 U24388 ( .A(U1_U0_y2[24]), .B(U1_U0_y0[24]), .CO(n8426), .S(n8423) );
  CMPR22X1 U24389 ( .A(U1_U0_y2[25]), .B(U1_U0_y0[25]), .CO(n8428), .S(n8425)
         );
  ADDHX2 U24390 ( .A(U1_U0_y2[26]), .B(U1_U0_y0[26]), .CO(n8431), .S(n8427) );
  CMPR22X1 U24391 ( .A(U1_U0_y2[34]), .B(U1_U0_y0[34]), .CO(n8448), .S(n8444)
         );
  NAND2X1 U24392 ( .A(n8424), .B(n8423), .Y(n8528) );
  INVX1 U24393 ( .A(n8624), .Y(n8452) );
  CMPR22X1 U24394 ( .A(U1_U0_y2[36]), .B(U1_U0_y0[36]), .CO(n8454), .S(n8450)
         );
  NOR2X1 U24395 ( .A(n8454), .B(n8453), .Y(n8626) );
  CMPR22X1 U24396 ( .A(U1_U0_y2[37]), .B(U1_U0_y0[37]), .CO(n8456), .S(n8453)
         );
  CMPR22X1 U24397 ( .A(U1_U0_y2[38]), .B(U1_U0_y0[38]), .CO(n8458), .S(n8455)
         );
  NAND2XL U24398 ( .A(n8470), .B(n8469), .Y(n8471) );
  NOR2XL U24399 ( .A(n12295), .B(U1_A_i_d0[5]), .Y(n16753) );
  NAND2XL U24400 ( .A(n8476), .B(n8533), .Y(n8477) );
  OR2X2 U24401 ( .A(n12296), .B(U1_A_i_d0[7]), .Y(n16740) );
  NAND2XL U24402 ( .A(n17020), .B(n16740), .Y(n8524) );
  INVXL U24403 ( .A(n8479), .Y(n8480) );
  OAI21XL U24404 ( .A0(n8514), .A1(n8481), .B0(n8480), .Y(n8492) );
  AOI21XL U24405 ( .A0(n8492), .A1(n8490), .B0(n8483), .Y(n8488) );
  INVXL U24406 ( .A(n8484), .Y(n8486) );
  NOR2XL U24407 ( .A(n12292), .B(U1_A_i_d0[4]), .Y(n16760) );
  XNOR2X1 U24408 ( .A(n8492), .B(n8491), .Y(n12291) );
  NOR2XL U24409 ( .A(n12291), .B(U1_A_i_d0[3]), .Y(n17036) );
  NOR2XL U24410 ( .A(n16760), .B(n17036), .Y(n8521) );
  INVXL U24411 ( .A(n8493), .Y(n8496) );
  AOI21XL U24412 ( .A0(n8496), .A1(n8495), .B0(n8494), .Y(n8497) );
  INVXL U24413 ( .A(n8497), .Y(n8502) );
  INVXL U24414 ( .A(n8498), .Y(n8501) );
  AOI21XL U24415 ( .A0(n8502), .A1(n8501), .B0(n8500), .Y(n8507) );
  NAND2XL U24416 ( .A(n12288), .B(U1_A_i_d0[1]), .Y(n16776) );
  INVXL U24417 ( .A(n16776), .Y(n8511) );
  AOI21XL U24418 ( .A0(n17046), .A1(n8510), .B0(n8511), .Y(n17043) );
  OAI21XL U24419 ( .A0(n8514), .A1(n8513), .B0(n8512), .Y(n8519) );
  INVXL U24420 ( .A(n8515), .Y(n8517) );
  NOR2XL U24421 ( .A(n12290), .B(U1_A_i_d0[2]), .Y(n16770) );
  OAI21XL U24422 ( .A0(n17043), .A1(n16770), .B0(n16771), .Y(n17034) );
  NAND2XL U24423 ( .A(n12291), .B(U1_A_i_d0[3]), .Y(n17035) );
  NAND2XL U24424 ( .A(n12292), .B(U1_A_i_d0[4]), .Y(n16761) );
  OAI21XL U24425 ( .A0(n16760), .A1(n17035), .B0(n16761), .Y(n8520) );
  AOI21XL U24426 ( .A0(n8521), .A1(n17034), .B0(n8520), .Y(n17018) );
  NAND2XL U24427 ( .A(n12295), .B(U1_A_i_d0[5]), .Y(n17024) );
  NAND2XL U24428 ( .A(n12296), .B(U1_A_i_d0[7]), .Y(n16739) );
  INVXL U24429 ( .A(n16739), .Y(n8522) );
  AOI21XL U24430 ( .A0(n17019), .A1(n16740), .B0(n8522), .Y(n8523) );
  INVXL U24431 ( .A(n8527), .Y(n8529) );
  NOR2XL U24432 ( .A(n19732), .B(U1_A_i_d0[9]), .Y(n16728) );
  NOR2XL U24433 ( .A(n12301), .B(U1_A_i_d0[8]), .Y(n17005) );
  INVXL U24434 ( .A(n17005), .Y(n16732) );
  NAND2XL U24435 ( .A(n8556), .B(n16732), .Y(n16996) );
  INVXL U24436 ( .A(n8543), .Y(n8545) );
  NAND2X1 U24437 ( .A(n8545), .B(n8544), .Y(n8546) );
  NOR2XL U24438 ( .A(n19734), .B(U1_A_i_d0[12]), .Y(n8547) );
  INVX1 U24439 ( .A(n8547), .Y(n16708) );
  NAND2XL U24440 ( .A(n12301), .B(U1_A_i_d0[8]), .Y(n17004) );
  INVXL U24441 ( .A(n17004), .Y(n8555) );
  NAND2XL U24442 ( .A(n19732), .B(U1_A_i_d0[9]), .Y(n17006) );
  OAI21XL U24443 ( .A0(n16722), .A1(n17006), .B0(n16723), .Y(n8554) );
  AOI21XL U24444 ( .A0(n8556), .A1(n8555), .B0(n8554), .Y(n16995) );
  NAND2XL U24445 ( .A(n19736), .B(U1_A_i_d0[11]), .Y(n16712) );
  INVXL U24446 ( .A(n16712), .Y(n16997) );
  NAND2XL U24447 ( .A(n19734), .B(U1_A_i_d0[12]), .Y(n16707) );
  INVXL U24448 ( .A(n16707), .Y(n8557) );
  OAI21XL U24449 ( .A0(n16995), .A1(n8559), .B0(n8558), .Y(n8560) );
  NOR2XL U24450 ( .A(n12313), .B(U1_A_i_d0[15]), .Y(n16980) );
  INVXL U24451 ( .A(n16980), .Y(n16688) );
  INVXL U24452 ( .A(n8570), .Y(n8572) );
  INVXL U24453 ( .A(n8576), .Y(n8578) );
  OR2X2 U24454 ( .A(n12311), .B(U1_A_i_d0[13]), .Y(n16988) );
  NAND2XL U24455 ( .A(n8580), .B(n16988), .Y(n16975) );
  INVXL U24456 ( .A(n8589), .Y(n8591) );
  OAI21X2 U24457 ( .A0(n8620), .A1(n8601), .B0(n8602), .Y(n8600) );
  NAND2X1 U24458 ( .A(n8598), .B(n8597), .Y(n8599) );
  NAND2XL U24459 ( .A(n8174), .B(n16674), .Y(n16959) );
  NAND2XL U24460 ( .A(n12311), .B(U1_A_i_d0[13]), .Y(n16698) );
  INVXL U24461 ( .A(n16698), .Y(n16987) );
  NAND2XL U24462 ( .A(n19754), .B(U1_A_i_d0[14]), .Y(n16694) );
  INVXL U24463 ( .A(n16694), .Y(n8605) );
  INVXL U24464 ( .A(n16979), .Y(n8607) );
  INVXL U24465 ( .A(n16684), .Y(n8606) );
  AOI21XL U24466 ( .A0(n8574), .A1(n8607), .B0(n8606), .Y(n8608) );
  OAI21XL U24467 ( .A0(n8609), .A1(n16976), .B0(n8608), .Y(n16957) );
  NAND2XL U24468 ( .A(n19756), .B(U1_A_i_d0[17]), .Y(n16967) );
  INVXL U24469 ( .A(n16967), .Y(n8611) );
  INVXL U24470 ( .A(n16670), .Y(n8610) );
  INVXL U24471 ( .A(n16961), .Y(n8612) );
  NOR2XL U24472 ( .A(n12327), .B(U1_A_i_d0[21]), .Y(n16951) );
  INVXL U24473 ( .A(n16951), .Y(n16650) );
  NAND2XL U24474 ( .A(n16650), .B(n8148), .Y(n16946) );
  NOR2XL U24475 ( .A(n19774), .B(U1_A_i_d0[23]), .Y(n16643) );
  NOR2XL U24476 ( .A(n16946), .B(n16643), .Y(n8631) );
  INVXL U24477 ( .A(n16950), .Y(n8629) );
  NAND2XL U24478 ( .A(n19773), .B(U1_A_i_d0[22]), .Y(n16648) );
  INVXL U24479 ( .A(n16648), .Y(n8628) );
  NAND2XL U24480 ( .A(n19774), .B(U1_A_i_d0[23]), .Y(n16644) );
  OAI21XL U24481 ( .A0(n16945), .A1(n16643), .B0(n16644), .Y(n8630) );
  NOR2XL U24482 ( .A(n12332), .B(U1_A_i_d0[24]), .Y(n16635) );
  NAND2XL U24483 ( .A(n12334), .B(U1_A_i_d0[25]), .Y(n16628) );
  MXI2X1 U24484 ( .A(U1_pipe4[27]), .B(n8640), .S0(n5812), .Y(n5095) );
  NOR2XL U24485 ( .A(n19724), .B(U1_A_i_d0[6]), .Y(n8652) );
  NOR2XL U24486 ( .A(n19723), .B(U1_A_i_d0[5]), .Y(n16744) );
  NAND2XL U24487 ( .A(n16738), .B(n8641), .Y(n8655) );
  INVX1 U24488 ( .A(n12292), .Y(n19718) );
  NOR2XL U24489 ( .A(n19718), .B(U1_A_i_d0[4]), .Y(n8648) );
  NOR2XL U24490 ( .A(n8648), .B(n16759), .Y(n8650) );
  NOR2XL U24491 ( .A(n16780), .B(U1_A_i_d0[0]), .Y(n16777) );
  OR2XL U24492 ( .A(n19711), .B(U1_A_i_d0[1]), .Y(n8643) );
  AOI21XL U24493 ( .A0(n8644), .A1(n8643), .B0(n8642), .Y(n16773) );
  OAI21XL U24494 ( .A0(n16773), .A1(n8646), .B0(n8645), .Y(n16757) );
  NAND2XL U24495 ( .A(n19718), .B(U1_A_i_d0[4]), .Y(n8647) );
  OAI21XL U24496 ( .A0(n8648), .A1(n16758), .B0(n8647), .Y(n8649) );
  AOI21XL U24497 ( .A0(n8650), .A1(n16757), .B0(n8649), .Y(n16736) );
  NAND2XL U24498 ( .A(n19723), .B(U1_A_i_d0[5]), .Y(n16745) );
  NAND2XL U24499 ( .A(n19724), .B(U1_A_i_d0[6]), .Y(n8651) );
  OAI21XL U24500 ( .A0(n8652), .A1(n16745), .B0(n8651), .Y(n16737) );
  AOI21XL U24501 ( .A0(n16737), .A1(n8641), .B0(n8653), .Y(n8654) );
  NOR2XL U24502 ( .A(n8657), .B(U1_A_i_d0[9]), .Y(n16718) );
  NOR2XL U24503 ( .A(n19737), .B(U1_A_i_d0[8]), .Y(n16717) );
  INVXL U24504 ( .A(n16717), .Y(n8656) );
  OR2X2 U24505 ( .A(n19744), .B(U1_A_i_d0[11]), .Y(n16706) );
  NOR2XL U24506 ( .A(n16704), .B(n8665), .Y(n8667) );
  NAND2XL U24507 ( .A(n19737), .B(U1_A_i_d0[8]), .Y(n16716) );
  INVXL U24508 ( .A(n16716), .Y(n8661) );
  NAND2XL U24509 ( .A(n8657), .B(U1_A_i_d0[9]), .Y(n16719) );
  NAND2XL U24510 ( .A(n19738), .B(U1_A_i_d0[10]), .Y(n8658) );
  OAI21XL U24511 ( .A0(n8659), .A1(n16719), .B0(n8658), .Y(n8660) );
  AOI21XL U24512 ( .A0(n8663), .A1(n16705), .B0(n8662), .Y(n8664) );
  OAI21XL U24513 ( .A0(n16703), .A1(n8665), .B0(n8664), .Y(n8666) );
  NOR2XL U24514 ( .A(n19760), .B(U1_A_i_d0[15]), .Y(n16683) );
  INVXL U24515 ( .A(n16683), .Y(n8668) );
  NAND2XL U24516 ( .A(n8672), .B(n8668), .Y(n8674) );
  INVX1 U24517 ( .A(n12311), .Y(n19757) );
  OR2X2 U24518 ( .A(n19757), .B(U1_A_i_d0[13]), .Y(n16693) );
  NAND2XL U24519 ( .A(n5786), .B(n16693), .Y(n16678) );
  NOR2XL U24520 ( .A(n8674), .B(n16678), .Y(n16656) );
  OR2X2 U24521 ( .A(n19767), .B(U1_A_i_d0[19]), .Y(n16660) );
  OR2X2 U24522 ( .A(n19765), .B(U1_A_i_d0[17]), .Y(n16669) );
  AND2X2 U24523 ( .A(n19757), .B(U1_A_i_d0[13]), .Y(n16692) );
  AOI21XL U24524 ( .A0(n5786), .A1(n16692), .B0(n8669), .Y(n16679) );
  NAND2XL U24525 ( .A(n19760), .B(U1_A_i_d0[15]), .Y(n16682) );
  INVXL U24526 ( .A(n16682), .Y(n8671) );
  AND2X2 U24527 ( .A(n19761), .B(U1_A_i_d0[16]), .Y(n8670) );
  AOI21XL U24528 ( .A0(n8672), .A1(n8671), .B0(n8670), .Y(n8673) );
  OAI21XL U24529 ( .A0(n8678), .A1(n16657), .B0(n8677), .Y(n8679) );
  NOR2XL U24530 ( .A(n19776), .B(U1_A_i_d0[21]), .Y(n16647) );
  NOR2XL U24531 ( .A(n19777), .B(U1_A_i_d0[22]), .Y(n8684) );
  NOR2XL U24532 ( .A(n16647), .B(n8684), .Y(n16640) );
  NOR2XL U24533 ( .A(n19775), .B(U1_A_i_d0[23]), .Y(n8682) );
  INVXL U24534 ( .A(n8682), .Y(n8686) );
  NAND2XL U24535 ( .A(n16640), .B(n8686), .Y(n16634) );
  INVX1 U24536 ( .A(n12332), .Y(n19782) );
  NAND2XL U24537 ( .A(n19777), .B(U1_A_i_d0[22]), .Y(n8683) );
  NAND2XL U24538 ( .A(n19782), .B(U1_A_i_d0[24]), .Y(n8687) );
  NAND2XL U24539 ( .A(n19786), .B(U1_A_i_d0[25]), .Y(n8688) );
  NOR2XL U24540 ( .A(U0_U2_y1[1]), .B(U0_U2_y0[1]), .Y(n8691) );
  INVXL U24541 ( .A(n8691), .Y(n8693) );
  AND2XL U24542 ( .A(U0_U2_y1[0]), .B(U0_U2_y0[0]), .Y(n8692) );
  AOI21XL U24543 ( .A0(n8693), .A1(n8692), .B0(n7995), .Y(n8701) );
  NOR2XL U24544 ( .A(U0_U2_y1[2]), .B(U0_U2_y0[2]), .Y(n8694) );
  INVXL U24545 ( .A(n8694), .Y(n8696) );
  NOR2XL U24546 ( .A(U0_U2_y1[3]), .B(U0_U2_y0[3]), .Y(n8695) );
  INVXL U24547 ( .A(n8695), .Y(n8698) );
  NAND2XL U24548 ( .A(n8696), .B(n8698), .Y(n8700) );
  AND2XL U24549 ( .A(U0_U2_y1[2]), .B(U0_U2_y0[2]), .Y(n8697) );
  AOI21XL U24550 ( .A0(n8698), .A1(n8697), .B0(n7993), .Y(n8699) );
  OAI21XL U24551 ( .A0(n8701), .A1(n8700), .B0(n8699), .Y(n8718) );
  NOR2XL U24552 ( .A(U0_U2_y1[5]), .B(U0_U2_y0[5]), .Y(n8703) );
  INVXL U24553 ( .A(n8703), .Y(n8710) );
  NAND2XL U24554 ( .A(n8704), .B(n8710), .Y(n8708) );
  NOR2XL U24555 ( .A(U0_U2_y1[6]), .B(U0_U2_y0[6]), .Y(n8705) );
  INVXL U24556 ( .A(n8705), .Y(n8707) );
  NOR2XL U24557 ( .A(U0_U2_y1[7]), .B(U0_U2_y0[7]), .Y(n8706) );
  INVXL U24558 ( .A(n8706), .Y(n8712) );
  NAND2XL U24559 ( .A(n8707), .B(n8712), .Y(n8714) );
  NOR2XL U24560 ( .A(n8708), .B(n8714), .Y(n8717) );
  AND2XL U24561 ( .A(U0_U2_y1[4]), .B(U0_U2_y0[4]), .Y(n8709) );
  AOI21XL U24562 ( .A0(n8710), .A1(n8709), .B0(n7943), .Y(n8715) );
  AOI21XL U24563 ( .A0(n8712), .A1(n8711), .B0(n7944), .Y(n8713) );
  OAI21XL U24564 ( .A0(n8715), .A1(n8714), .B0(n8713), .Y(n8716) );
  OR2X2 U24565 ( .A(n8732), .B(U0_U2_y0[13]), .Y(n8734) );
  NAND2XL U24566 ( .A(n8734), .B(n8719), .Y(n8864) );
  NOR2X1 U24567 ( .A(n8735), .B(U0_U2_y1[13]), .Y(n8869) );
  NOR2X1 U24568 ( .A(n8864), .B(n8869), .Y(n8737) );
  OR2X2 U24569 ( .A(U0_U2_y1[9]), .B(U0_U2_y0[9]), .Y(n8725) );
  OR2X2 U24570 ( .A(U0_U2_y1[11]), .B(U0_U2_y0[11]), .Y(n8728) );
  OAI21XL U24571 ( .A0(n8731), .A1(n8730), .B0(n8729), .Y(n8860) );
  OAI21XL U24572 ( .A0(n8865), .A1(n8869), .B0(n8870), .Y(n8736) );
  CMPR22X1 U24573 ( .A(U0_U2_y1[17]), .B(U0_U2_y0[17]), .CO(n8745), .S(n8742)
         );
  CMPR22X1 U24574 ( .A(U0_U2_y1[19]), .B(U0_U2_y0[19]), .CO(n8749), .S(n8746)
         );
  NOR2X2 U24575 ( .A(n8749), .B(n8748), .Y(n8824) );
  INVXL U24576 ( .A(n8824), .Y(n8750) );
  XNOR2X2 U24577 ( .A(n8752), .B(n8751), .Y(n24608) );
  OR2XL U24578 ( .A(U0_U1_y1[1]), .B(U0_U1_y0[1]), .Y(n8755) );
  AND2XL U24579 ( .A(U0_U1_y1[0]), .B(U0_U1_y0[0]), .Y(n8754) );
  AOI21XL U24580 ( .A0(n8755), .A1(n8754), .B0(n8753), .Y(n8762) );
  NAND2XL U24581 ( .A(n8756), .B(n8759), .Y(n8761) );
  AND2XL U24582 ( .A(U0_U1_y1[2]), .B(U0_U1_y0[2]), .Y(n8758) );
  AOI21XL U24583 ( .A0(n8759), .A1(n8758), .B0(n8757), .Y(n8760) );
  OAI21XL U24584 ( .A0(n8762), .A1(n8761), .B0(n8760), .Y(n8777) );
  OR2X2 U24585 ( .A(U0_U1_y1[7]), .B(U0_U1_y0[7]), .Y(n8771) );
  AOI21XL U24586 ( .A0(n8768), .A1(n8767), .B0(n8766), .Y(n8774) );
  AOI21XL U24587 ( .A0(n8771), .A1(n8770), .B0(n8769), .Y(n8772) );
  OAI21XL U24588 ( .A0(n8774), .A1(n8773), .B0(n8772), .Y(n8775) );
  AOI21XL U24589 ( .A0(n8777), .A1(n8776), .B0(n8775), .Y(n8874) );
  OR2X2 U24590 ( .A(U0_U1_y1[12]), .B(U0_U1_y0[12]), .Y(n8778) );
  NAND2XL U24591 ( .A(n8794), .B(n8778), .Y(n8879) );
  OR2X2 U24592 ( .A(U0_U1_y1[10]), .B(U0_U1_y0[10]), .Y(n8781) );
  OAI21XL U24593 ( .A0(n8790), .A1(n8789), .B0(n8788), .Y(n8875) );
  NAND2XL U24594 ( .A(n8795), .B(U0_U1_y1[13]), .Y(n8885) );
  OAI21XL U24595 ( .A0(n8880), .A1(n8884), .B0(n8885), .Y(n8796) );
  CMPR22X1 U24596 ( .A(U0_U1_y1[14]), .B(U0_U1_y0[14]), .CO(n8801), .S(n8795)
         );
  NOR2XL U24597 ( .A(n8855), .B(n8845), .Y(n8905) );
  NAND2X1 U24598 ( .A(n8905), .B(n8809), .Y(n8931) );
  NAND2XL U24599 ( .A(n8803), .B(n8802), .Y(n8846) );
  OAI21XL U24600 ( .A0(n8845), .A1(n8856), .B0(n8846), .Y(n8906) );
  NAND2XL U24601 ( .A(n8807), .B(n8806), .Y(n8913) );
  OAI21XL U24602 ( .A0(n8912), .A1(n8921), .B0(n8913), .Y(n8808) );
  CMPR22X1 U24603 ( .A(U0_U1_y1[18]), .B(U0_U1_y0[18]), .CO(n8811), .S(n8806)
         );
  INVXL U24604 ( .A(n8833), .Y(n8814) );
  NOR2XL U24605 ( .A(n24608), .B(n24582), .Y(n25081) );
  INVXL U24606 ( .A(n8830), .Y(n8818) );
  NAND2XL U24607 ( .A(n8818), .B(n8832), .Y(n8819) );
  NOR2XL U24608 ( .A(n25081), .B(n25079), .Y(n25074) );
  ADDHX2 U24609 ( .A(U0_U2_y1[20]), .B(U0_U2_y0[20]), .CO(n8827), .S(n8748) );
  AOI21XL U24610 ( .A0(n8834), .A1(n8930), .B0(n8935), .Y(n8973) );
  XOR2X1 U24611 ( .A(n8973), .B(n8838), .Y(n24584) );
  NAND2XL U24612 ( .A(n25074), .B(n8839), .Y(n8929) );
  OAI21XL U24613 ( .A0(n8897), .A1(n8851), .B0(n8852), .Y(n8844) );
  XNOR2X1 U24614 ( .A(n8844), .B(n8843), .Y(n24596) );
  OAI21XL U24615 ( .A0(n8909), .A1(n8855), .B0(n8856), .Y(n8849) );
  INVXL U24616 ( .A(n8851), .Y(n8853) );
  NAND2XL U24617 ( .A(n8853), .B(n8852), .Y(n8854) );
  XOR2X1 U24618 ( .A(n8909), .B(n8858), .Y(n24588) );
  NOR2XL U24619 ( .A(n24590), .B(n24588), .Y(n25107) );
  INVXL U24620 ( .A(n25107), .Y(n24847) );
  NAND2XL U24621 ( .A(n8850), .B(n24847), .Y(n8892) );
  INVXL U24622 ( .A(n8859), .Y(n8862) );
  AOI21XL U24623 ( .A0(n8862), .A1(n8861), .B0(n8860), .Y(n8863) );
  INVXL U24624 ( .A(n8863), .Y(n8868) );
  AOI21XL U24625 ( .A0(n8868), .A1(n8867), .B0(n8866), .Y(n8873) );
  INVXL U24626 ( .A(n8869), .Y(n8871) );
  INVXL U24627 ( .A(n8874), .Y(n8877) );
  AOI21XL U24628 ( .A0(n8877), .A1(n8876), .B0(n8875), .Y(n8878) );
  INVXL U24629 ( .A(n8878), .Y(n8883) );
  AOI21XL U24630 ( .A0(n8883), .A1(n8882), .B0(n8881), .Y(n8888) );
  NAND2XL U24631 ( .A(n24590), .B(n24588), .Y(n25106) );
  INVXL U24632 ( .A(n25106), .Y(n8890) );
  NAND2XL U24633 ( .A(n24596), .B(n24595), .Y(n24843) );
  INVXL U24634 ( .A(n24843), .Y(n8889) );
  AOI21XL U24635 ( .A0(n8850), .A1(n8890), .B0(n8889), .Y(n8891) );
  INVXL U24636 ( .A(n8893), .Y(n8896) );
  INVXL U24637 ( .A(n8894), .Y(n8895) );
  AOI21XL U24638 ( .A0(n8920), .A1(n8918), .B0(n8899), .Y(n8904) );
  NAND2XL U24639 ( .A(n8902), .B(n8901), .Y(n8903) );
  INVXL U24640 ( .A(n8905), .Y(n8908) );
  INVXL U24641 ( .A(n8906), .Y(n8907) );
  OAI21XL U24642 ( .A0(n8909), .A1(n8908), .B0(n8907), .Y(n8924) );
  AOI21XL U24643 ( .A0(n8924), .A1(n8922), .B0(n8911), .Y(n8916) );
  XOR2X1 U24644 ( .A(n8916), .B(n8915), .Y(n24586) );
  NOR2XL U24645 ( .A(n24602), .B(n24586), .Y(n25096) );
  NAND2XL U24646 ( .A(n8918), .B(n8917), .Y(n8919) );
  NOR2XL U24647 ( .A(n24600), .B(n24587), .Y(n25095) );
  NOR2XL U24648 ( .A(n25096), .B(n25095), .Y(n8926) );
  NAND2XL U24649 ( .A(n24600), .B(n24587), .Y(n25094) );
  NAND2XL U24650 ( .A(n24602), .B(n24586), .Y(n25097) );
  OAI21XL U24651 ( .A0(n25096), .A1(n25094), .B0(n25097), .Y(n8925) );
  NAND2XL U24652 ( .A(n24606), .B(n24583), .Y(n25087) );
  NAND2XL U24653 ( .A(n24608), .B(n24582), .Y(n25082) );
  OAI21XL U24654 ( .A0(n25081), .A1(n25087), .B0(n25082), .Y(n25073) );
  NAND2XL U24655 ( .A(n24610), .B(n24584), .Y(n25075) );
  INVXL U24656 ( .A(n25075), .Y(n8927) );
  AOI21XL U24657 ( .A0(n25073), .A1(n8839), .B0(n8927), .Y(n8928) );
  NOR2X2 U24658 ( .A(n8933), .B(n8932), .Y(n8974) );
  OAI21XL U24659 ( .A0(n8974), .A1(n8971), .B0(n8975), .Y(n8934) );
  CMPR22X1 U24660 ( .A(U0_U1_y1[22]), .B(U0_U1_y0[22]), .CO(n8940), .S(n8932)
         );
  INVXL U24661 ( .A(n8982), .Y(n8944) );
  CMPR22X1 U24662 ( .A(U0_U2_y1[21]), .B(U0_U2_y0[21]), .CO(n8950), .S(n8826)
         );
  NAND2X1 U24663 ( .A(n8955), .B(n8954), .Y(n8992) );
  AOI21X2 U24664 ( .A0(n5821), .A1(n8963), .B0(n8956), .Y(n8960) );
  CMPR22X1 U24665 ( .A(U0_U2_y1[23]), .B(U0_U2_y0[23]), .CO(n8957), .S(n8954)
         );
  INVXL U24666 ( .A(n8993), .Y(n8958) );
  NAND2XL U24667 ( .A(n8961), .B(n8981), .Y(n8962) );
  XNOR2X1 U24668 ( .A(n9062), .B(n8962), .Y(n24616) );
  NAND2XL U24669 ( .A(n8963), .B(n8992), .Y(n8964) );
  NOR2XL U24670 ( .A(n24616), .B(n24623), .Y(n24802) );
  OAI21XL U24671 ( .A0(n8973), .A1(n8972), .B0(n8971), .Y(n8978) );
  NOR2XL U24672 ( .A(n24621), .B(n24617), .Y(n25059) );
  INVXL U24673 ( .A(n25059), .Y(n24806) );
  NAND2XL U24674 ( .A(n9007), .B(n24806), .Y(n25050) );
  NOR2X1 U24675 ( .A(n8984), .B(n8983), .Y(n9042) );
  NOR2X2 U24676 ( .A(n8986), .B(n8985), .Y(n9046) );
  INVXL U24677 ( .A(n9046), .Y(n8987) );
  NAND2XL U24678 ( .A(n8986), .B(n8985), .Y(n9044) );
  NAND2X1 U24679 ( .A(n8987), .B(n9044), .Y(n8988) );
  XNOR2X2 U24680 ( .A(n8989), .B(n8988), .Y(n24619) );
  CMPR22X1 U24681 ( .A(U0_U2_y1[25]), .B(U0_U2_y0[25]), .CO(n8996), .S(n8994)
         );
  INVXL U24682 ( .A(n9016), .Y(n8997) );
  INVXL U24683 ( .A(n9042), .Y(n8999) );
  INVXL U24684 ( .A(n25058), .Y(n9006) );
  NAND2XL U24685 ( .A(n24616), .B(n24623), .Y(n25060) );
  OAI21XL U24686 ( .A0(n24796), .A1(n25060), .B0(n24797), .Y(n9005) );
  AOI21XL U24687 ( .A0(n9007), .A1(n9006), .B0(n9005), .Y(n25049) );
  NAND2XL U24688 ( .A(n24619), .B(n24633), .Y(n24780) );
  INVXL U24689 ( .A(n24780), .Y(n9008) );
  CMPR22X1 U24690 ( .A(U0_U2_y1[27]), .B(U0_U2_y0[27]), .CO(n9021), .S(n9018)
         );
  CMPR22X1 U24691 ( .A(U0_U2_y1[30]), .B(U0_U2_y0[30]), .CO(n9030), .S(n9024)
         );
  INVXL U24692 ( .A(n9153), .Y(n9040) );
  NAND2X1 U24693 ( .A(n9040), .B(n9151), .Y(n9041) );
  NOR2X2 U24694 ( .A(n9042), .B(n9046), .Y(n9049) );
  NAND2X1 U24695 ( .A(n9043), .B(n9049), .Y(n9094) );
  ADDHX2 U24696 ( .A(U0_U1_y1[28]), .B(U0_U1_y0[28]), .CO(n9055), .S(n9052) );
  AOI21X2 U24697 ( .A0(n9059), .A1(n9095), .B0(n9058), .Y(n9060) );
  INVXL U24698 ( .A(n9166), .Y(n9071) );
  INVXL U24699 ( .A(n25011), .Y(n9078) );
  NAND2X1 U24700 ( .A(n8035), .B(n9078), .Y(n9144) );
  NAND2X1 U24701 ( .A(n9082), .B(n9081), .Y(n9083) );
  INVXL U24702 ( .A(n9084), .Y(n9086) );
  NAND2X1 U24703 ( .A(n5793), .B(n9088), .Y(n9089) );
  XOR2X2 U24704 ( .A(n9107), .B(n9098), .Y(n24645) );
  NOR2XL U24705 ( .A(n24645), .B(n24652), .Y(n25031) );
  INVXL U24706 ( .A(n25031), .Y(n25034) );
  INVXL U24707 ( .A(n9115), .Y(n9117) );
  NAND2XL U24708 ( .A(n25034), .B(n7014), .Y(n9140) );
  NAND2X1 U24709 ( .A(n9121), .B(n9120), .Y(n9122) );
  INVXL U24710 ( .A(n9124), .Y(n9126) );
  XOR2X1 U24711 ( .A(n9135), .B(n9134), .Y(n24649) );
  NAND2XL U24712 ( .A(n25040), .B(n9136), .Y(n25027) );
  NAND2XL U24713 ( .A(n24647), .B(n24649), .Y(n25044) );
  INVXL U24714 ( .A(n25044), .Y(n25038) );
  INVXL U24715 ( .A(n25039), .Y(n9137) );
  INVXL U24716 ( .A(n25033), .Y(n9138) );
  AOI21XL U24717 ( .A0(n7014), .A1(n9138), .B0(n8086), .Y(n9139) );
  NAND2XL U24718 ( .A(n24661), .B(n24643), .Y(n25024) );
  INVXL U24719 ( .A(n25024), .Y(n9141) );
  AOI21X1 U24720 ( .A0(n9146), .A1(n25007), .B0(n9145), .Y(n9147) );
  INVXL U24721 ( .A(n9183), .Y(n9157) );
  AOI21XL U24722 ( .A0(n7738), .A1(n9157), .B0(n9156), .Y(n9161) );
  CMPR22X1 U24723 ( .A(U0_U2_y1[34]), .B(U0_U2_y0[34]), .CO(n9159), .S(n9038)
         );
  CMPR22X1 U24724 ( .A(U0_U1_y1[34]), .B(U0_U1_y0[34]), .CO(n9171), .S(n9069)
         );
  NOR2X1 U24725 ( .A(n9171), .B(n9170), .Y(n9178) );
  NOR2XL U24726 ( .A(n24679), .B(n24674), .Y(n24997) );
  INVXL U24727 ( .A(n24997), .Y(n25002) );
  CMPR22X1 U24728 ( .A(U0_U1_y1[35]), .B(U0_U1_y0[35]), .CO(n9182), .S(n9170)
         );
  NOR2XL U24729 ( .A(n24675), .B(n24680), .Y(n9194) );
  NAND2XL U24730 ( .A(n25002), .B(n24721), .Y(n24993) );
  CMPR22X1 U24731 ( .A(U0_U1_y1[36]), .B(U0_U1_y0[36]), .CO(n9198), .S(n9181)
         );
  NOR2X1 U24732 ( .A(n9198), .B(n9197), .Y(n9213) );
  NOR2X1 U24733 ( .A(n9205), .B(n9204), .Y(n9220) );
  NOR2XL U24734 ( .A(n24676), .B(n24684), .Y(n24714) );
  NAND2XL U24735 ( .A(n24679), .B(n24674), .Y(n25001) );
  INVXL U24736 ( .A(n25001), .Y(n9209) );
  NAND2XL U24737 ( .A(n24675), .B(n24680), .Y(n24720) );
  INVXL U24738 ( .A(n24720), .Y(n9208) );
  AOI21XL U24739 ( .A0(n9209), .A1(n24721), .B0(n9208), .Y(n24992) );
  NAND2XL U24740 ( .A(n24676), .B(n24684), .Y(n24715) );
  CMPR22X1 U24741 ( .A(U0_U1_y1[37]), .B(U0_U1_y0[37]), .CO(n9217), .S(n9197)
         );
  CMPR22X1 U24742 ( .A(U0_U2_y1[37]), .B(U0_U2_y0[37]), .CO(n9223), .S(n9204)
         );
  CMPR22X1 U24743 ( .A(U0_U1_y1[38]), .B(U0_U1_y0[38]), .CO(n9229), .S(n9216)
         );
  NOR2X1 U24744 ( .A(n9229), .B(n9228), .Y(n12344) );
  CMPR22X1 U24745 ( .A(U0_U2_y1[38]), .B(U0_U2_y0[38]), .CO(n9235), .S(n9222)
         );
  CLKINVX3 U24746 ( .A(n5837), .Y(n25101) );
  CMPR22X1 U24747 ( .A(U1_U0_y1[17]), .B(U1_U0_y0[17]), .CO(n9297), .S(n9294)
         );
  CMPR22X1 U24748 ( .A(U1_U0_y1[20]), .B(U1_U0_y0[20]), .CO(n9305), .S(n9302)
         );
  OR2X2 U24749 ( .A(U1_U0_y1[3]), .B(U1_U0_y0[3]), .Y(n9248) );
  NAND2XL U24750 ( .A(n9245), .B(n9248), .Y(n9250) );
  OAI21XL U24751 ( .A0(n9251), .A1(n9250), .B0(n9249), .Y(n9268) );
  OR2X2 U24752 ( .A(U1_U0_y1[5]), .B(U1_U0_y0[5]), .Y(n9259) );
  OR2X2 U24753 ( .A(U1_U0_y1[7]), .B(U1_U0_y0[7]), .Y(n9262) );
  OAI21XL U24754 ( .A0(n9265), .A1(n9264), .B0(n9263), .Y(n9266) );
  NOR2XL U24755 ( .A(U1_U0_y1[12]), .B(U1_U0_y0[12]), .Y(n9269) );
  INVXL U24756 ( .A(n9269), .Y(n9270) );
  CMPR22X1 U24757 ( .A(U1_U0_y1[14]), .B(U1_U0_y0[14]), .CO(n9291), .S(n9287)
         );
  OR2X2 U24758 ( .A(U1_U0_y1[9]), .B(U1_U0_y0[9]), .Y(n9278) );
  NAND2XL U24759 ( .A(n9288), .B(n9382), .Y(n9289) );
  OAI21XL U24760 ( .A0(n9284), .A1(n9283), .B0(n9282), .Y(n9381) );
  AOI21XL U24761 ( .A0(n9286), .A1(n9285), .B0(n8141), .Y(n9385) );
  NAND2XL U24762 ( .A(n9293), .B(n9292), .Y(n9405) );
  NAND2X1 U24763 ( .A(n9297), .B(n9296), .Y(n9373) );
  CMPR22X1 U24764 ( .A(U1_U0_y1[23]), .B(U1_U0_y0[23]), .CO(n9311), .S(n9308)
         );
  CMPR22X1 U24765 ( .A(U1_U0_y1[31]), .B(U1_U0_y0[31]), .CO(n9327), .S(n9324)
         );
  NOR2X2 U24766 ( .A(n9327), .B(n9326), .Y(n9492) );
  CMPR22X1 U24767 ( .A(U1_U0_y1[32]), .B(U1_U0_y0[32]), .CO(n9329), .S(n9326)
         );
  CMPR22X1 U24768 ( .A(U1_U0_y1[33]), .B(U1_U0_y0[33]), .CO(n9331), .S(n9328)
         );
  CMPR22X1 U24769 ( .A(U1_U0_y1[34]), .B(U1_U0_y0[34]), .CO(n9334), .S(n9330)
         );
  NAND2X2 U24770 ( .A(n9325), .B(n9324), .Y(n9498) );
  OR2X2 U24771 ( .A(n9337), .B(n9336), .Y(n9527) );
  NAND2X1 U24772 ( .A(n9337), .B(n9336), .Y(n9526) );
  CMPR22X1 U24773 ( .A(U1_U0_y1[36]), .B(U1_U0_y0[36]), .CO(n9340), .S(n9336)
         );
  NAND2X1 U24774 ( .A(n9340), .B(n9339), .Y(n9529) );
  CMPR22X1 U24775 ( .A(U1_U0_y1[38]), .B(U1_U0_y0[38]), .CO(n9346), .S(n9342)
         );
  NOR2X1 U24776 ( .A(n9346), .B(n9345), .Y(n9542) );
  XOR2X1 U24777 ( .A(U1_U0_y0[40]), .B(U1_U0_y1[40]), .Y(n9348) );
  INVXL U24778 ( .A(n9353), .Y(n9355) );
  NOR2XL U24779 ( .A(n9665), .B(U1_A_i_d0[6]), .Y(n9416) );
  NOR2XL U24780 ( .A(n9664), .B(U1_A_i_d0[5]), .Y(n17564) );
  NOR2XL U24781 ( .A(n9416), .B(n17564), .Y(n17559) );
  INVXL U24782 ( .A(n9431), .Y(n9363) );
  NAND2XL U24783 ( .A(n9363), .B(n9430), .Y(n9364) );
  XOR2X1 U24784 ( .A(n9432), .B(n9364), .Y(n13676) );
  INVX1 U24785 ( .A(n13676), .Y(n9668) );
  NAND2XL U24786 ( .A(n17559), .B(n9365), .Y(n9419) );
  INVXL U24787 ( .A(n9372), .Y(n9374) );
  NOR2XL U24788 ( .A(n9659), .B(U1_A_i_d0[4]), .Y(n9412) );
  NOR2XL U24789 ( .A(n9658), .B(U1_A_i_d0[3]), .Y(n17578) );
  NOR2XL U24790 ( .A(n9412), .B(n17578), .Y(n9414) );
  INVXL U24791 ( .A(n13667), .Y(n9397) );
  NOR2XL U24792 ( .A(n9397), .B(U1_A_i_d0[1]), .Y(n9396) );
  INVXL U24793 ( .A(n9396), .Y(n9399) );
  AOI21XL U24794 ( .A0(n9400), .A1(n9399), .B0(n9398), .Y(n17588) );
  OAI21XL U24795 ( .A0(n17588), .A1(n9410), .B0(n9409), .Y(n17576) );
  NAND2XL U24796 ( .A(n9659), .B(U1_A_i_d0[4]), .Y(n9411) );
  OAI21XL U24797 ( .A0(n9412), .A1(n17577), .B0(n9411), .Y(n9413) );
  AOI21XL U24798 ( .A0(n9414), .A1(n17576), .B0(n9413), .Y(n17557) );
  NAND2XL U24799 ( .A(n9664), .B(U1_A_i_d0[5]), .Y(n17565) );
  OAI21XL U24800 ( .A0(n9416), .A1(n17565), .B0(n9415), .Y(n17558) );
  AOI21XL U24801 ( .A0(n17558), .A1(n9365), .B0(n9417), .Y(n9418) );
  AOI21X2 U24802 ( .A0(n7628), .A1(n9428), .B0(n9421), .Y(n9426) );
  INVXL U24803 ( .A(n9422), .Y(n9424) );
  NOR2XL U24804 ( .A(n9449), .B(U1_A_i_d0[9]), .Y(n17541) );
  NOR2X1 U24805 ( .A(n9452), .B(n17541), .Y(n9455) );
  INVX1 U24806 ( .A(n13681), .Y(n9674) );
  NOR2XL U24807 ( .A(n9674), .B(U1_A_i_d0[8]), .Y(n17540) );
  INVXL U24808 ( .A(n17540), .Y(n9436) );
  NAND2XL U24809 ( .A(n9455), .B(n9436), .Y(n17528) );
  OAI21X1 U24810 ( .A0(n9448), .A1(n9444), .B0(n9445), .Y(n9443) );
  INVXL U24811 ( .A(n9439), .Y(n9441) );
  INVXL U24812 ( .A(n9444), .Y(n9446) );
  NAND2XL U24813 ( .A(n9674), .B(U1_A_i_d0[8]), .Y(n17539) );
  INVXL U24814 ( .A(n17539), .Y(n9454) );
  NAND2XL U24815 ( .A(n9449), .B(U1_A_i_d0[9]), .Y(n17542) );
  NAND2XL U24816 ( .A(n9450), .B(U1_A_i_d0[10]), .Y(n9451) );
  AOI21XL U24817 ( .A0(n7007), .A1(n17529), .B0(n9456), .Y(n9457) );
  INVXL U24818 ( .A(n9464), .Y(n9466) );
  NAND2X1 U24819 ( .A(n9466), .B(n9465), .Y(n9467) );
  INVXL U24820 ( .A(n17507), .Y(n9471) );
  OR2X2 U24821 ( .A(n9690), .B(U1_A_i_d0[13]), .Y(n17517) );
  NAND2XL U24822 ( .A(n9503), .B(n17517), .Y(n17502) );
  INVXL U24823 ( .A(n9486), .Y(n9488) );
  NAND2X1 U24824 ( .A(n9488), .B(n9487), .Y(n9489) );
  OR2X2 U24825 ( .A(n9512), .B(U1_A_i_d0[19]), .Y(n17482) );
  NAND2X1 U24826 ( .A(n9513), .B(n17482), .Y(n9515) );
  INVXL U24827 ( .A(n9492), .Y(n9494) );
  XNOR2X4 U24828 ( .A(n9496), .B(n9495), .Y(n13699) );
  INVXL U24829 ( .A(n9497), .Y(n9499) );
  OR2X2 U24830 ( .A(n9700), .B(U1_A_i_d0[17]), .Y(n17493) );
  NAND2X1 U24831 ( .A(n9511), .B(n17493), .Y(n17480) );
  NOR2X1 U24832 ( .A(n9515), .B(n17480), .Y(n9517) );
  AOI21XL U24833 ( .A0(n9503), .A1(n17516), .B0(n9502), .Y(n17503) );
  NAND2XL U24834 ( .A(n9504), .B(U1_A_i_d0[15]), .Y(n17506) );
  INVXL U24835 ( .A(n17506), .Y(n9506) );
  AND2X2 U24836 ( .A(n9700), .B(U1_A_i_d0[17]), .Y(n17492) );
  AND2X2 U24837 ( .A(n9701), .B(U1_A_i_d0[18]), .Y(n9510) );
  AOI21X1 U24838 ( .A0(n9511), .A1(n17492), .B0(n9510), .Y(n17479) );
  OAI21XL U24839 ( .A0(n9515), .A1(n17479), .B0(n9514), .Y(n9516) );
  NOR2X1 U24840 ( .A(n5848), .B(U1_A_i_d0[21]), .Y(n17470) );
  NOR2X1 U24841 ( .A(n9712), .B(U1_A_i_d0[22]), .Y(n9536) );
  NOR2X1 U24842 ( .A(n17470), .B(n9536), .Y(n17461) );
  INVXL U24843 ( .A(n9528), .Y(n9530) );
  XOR2X4 U24844 ( .A(n9532), .B(n9531), .Y(n13713) );
  NAND2X1 U24845 ( .A(n13713), .B(n8156), .Y(n9539) );
  NAND2XL U24846 ( .A(n9712), .B(U1_A_i_d0[22]), .Y(n9535) );
  NAND2XL U24847 ( .A(n9717), .B(U1_A_i_d0[24]), .Y(n9540) );
  NOR2XL U24848 ( .A(n9720), .B(U1_A_i_d0[25]), .Y(n9548) );
  MXI2X1 U24849 ( .A(U1_pipe10[27]), .B(n9549), .S0(n24784), .Y(n4865) );
  XNOR2X1 U24850 ( .A(n9552), .B(BOPA[32]), .Y(n9551) );
  NAND2XL U24851 ( .A(n11418), .B(BOPA[6]), .Y(n9550) );
  NAND2X1 U24852 ( .A(n11418), .B(BOPA[7]), .Y(n9553) );
  OAI21XL U24853 ( .A0(n9555), .A1(n10601), .B0(n9554), .Y(n9556) );
  AOI21X1 U24854 ( .A0(n9557), .A1(n10596), .B0(n9556), .Y(n9558) );
  NOR2X1 U24855 ( .A(n7055), .B(BOPB[42]), .Y(n10592) );
  NOR2X1 U24856 ( .A(n8175), .B(BOPB[43]), .Y(n10587) );
  NOR2XL U24857 ( .A(n10592), .B(n10587), .Y(n10579) );
  NOR2X1 U24858 ( .A(n8171), .B(BOPB[44]), .Y(n10570) );
  NOR2X1 U24859 ( .A(n8169), .B(BOPB[45]), .Y(n10574) );
  NOR2X1 U24860 ( .A(n10570), .B(n10574), .Y(n9561) );
  NOR2XL U24861 ( .A(n10550), .B(n10542), .Y(n9563) );
  NAND2XL U24862 ( .A(n10548), .B(n9563), .Y(n9565) );
  NOR2XL U24863 ( .A(n10565), .B(n9565), .Y(n10671) );
  NAND2X1 U24864 ( .A(n7055), .B(BOPB[42]), .Y(n10593) );
  AOI21X2 U24865 ( .A0(n9561), .A1(n10580), .B0(n9560), .Y(n10564) );
  NAND2XL U24866 ( .A(n8160), .B(BOPB[47]), .Y(n10560) );
  NAND2XL U24867 ( .A(n8157), .B(BOPB[48]), .Y(n10551) );
  NAND2XL U24868 ( .A(n8153), .B(BOPB[49]), .Y(n10543) );
  OAI21XL U24869 ( .A0(n10542), .A1(n10551), .B0(n10543), .Y(n9562) );
  AOI21XL U24870 ( .A0(n9563), .A1(n10547), .B0(n9562), .Y(n9564) );
  OAI21XL U24871 ( .A0(n10564), .A1(n9565), .B0(n9564), .Y(n10677) );
  INVXL U24872 ( .A(n10677), .Y(n9566) );
  NAND2X1 U24873 ( .A(n10530), .B(n10673), .Y(n9568) );
  NOR2XL U24874 ( .A(n13675), .B(U1_A_i_d0[6]), .Y(n17268) );
  NOR2XL U24875 ( .A(n17268), .B(n17266), .Y(n17261) );
  OR2X2 U24876 ( .A(n13676), .B(U1_A_i_d0[7]), .Y(n17263) );
  NAND2XL U24877 ( .A(n17261), .B(n17263), .Y(n9576) );
  NOR2XL U24878 ( .A(n17278), .B(n17283), .Y(n9573) );
  NAND2XL U24879 ( .A(n13667), .B(U1_A_i_d0[1]), .Y(n17293) );
  INVXL U24880 ( .A(n17293), .Y(n9571) );
  AOI21XL U24881 ( .A0(n17294), .A1(n9570), .B0(n9571), .Y(n17291) );
  OAI21XL U24882 ( .A0(n17291), .A1(n17288), .B0(n17289), .Y(n17277) );
  NAND2XL U24883 ( .A(n13670), .B(U1_A_i_d0[3]), .Y(n17284) );
  NAND2XL U24884 ( .A(n13671), .B(U1_A_i_d0[4]), .Y(n17279) );
  AOI21XL U24885 ( .A0(n9573), .A1(n17277), .B0(n9572), .Y(n17259) );
  NAND2XL U24886 ( .A(n13674), .B(U1_A_i_d0[5]), .Y(n17273) );
  NAND2XL U24887 ( .A(n13675), .B(U1_A_i_d0[6]), .Y(n17269) );
  OAI21XL U24888 ( .A0(n17268), .A1(n17273), .B0(n17269), .Y(n17260) );
  AOI21XL U24889 ( .A0(n17260), .A1(n17263), .B0(n9574), .Y(n9575) );
  OAI21XL U24890 ( .A0(n9576), .A1(n17259), .B0(n9575), .Y(n17232) );
  NOR2XL U24891 ( .A(n13682), .B(U1_A_i_d0[9]), .Y(n17243) );
  NAND2XL U24892 ( .A(n9580), .B(n17256), .Y(n17234) );
  NAND2XL U24893 ( .A(n13681), .B(U1_A_i_d0[8]), .Y(n17255) );
  INVXL U24894 ( .A(n17255), .Y(n9579) );
  NAND2XL U24895 ( .A(n13682), .B(U1_A_i_d0[9]), .Y(n17251) );
  NAND2XL U24896 ( .A(n13683), .B(U1_A_i_d0[10]), .Y(n17246) );
  OAI21XL U24897 ( .A0(n17245), .A1(n17251), .B0(n17246), .Y(n9578) );
  NAND2XL U24898 ( .A(n13687), .B(U1_A_i_d0[11]), .Y(n17239) );
  INVXL U24899 ( .A(n17236), .Y(n9581) );
  OR2X2 U24900 ( .A(n13691), .B(U1_A_i_d0[13]), .Y(n17229) );
  NOR2XL U24901 ( .A(n13702), .B(U1_A_i_d0[19]), .Y(n13726) );
  INVXL U24902 ( .A(n13726), .Y(n17199) );
  NOR2XL U24903 ( .A(n13698), .B(U1_A_i_d0[17]), .Y(n17202) );
  INVXL U24904 ( .A(n17202), .Y(n17208) );
  NAND2X1 U24905 ( .A(n13721), .B(n9598), .Y(n9600) );
  NAND2XL U24906 ( .A(n13691), .B(U1_A_i_d0[13]), .Y(n17228) );
  INVXL U24907 ( .A(n17228), .Y(n17224) );
  NAND2XL U24908 ( .A(n13692), .B(U1_A_i_d0[14]), .Y(n17225) );
  INVXL U24909 ( .A(n17225), .Y(n9586) );
  AOI21XL U24910 ( .A0(n6996), .A1(n17224), .B0(n9586), .Y(n17212) );
  INVXL U24911 ( .A(n17220), .Y(n9588) );
  INVXL U24912 ( .A(n17216), .Y(n9587) );
  AOI21XL U24913 ( .A0(n17217), .A1(n9588), .B0(n9587), .Y(n9589) );
  OAI21X1 U24914 ( .A0(n9590), .A1(n17212), .B0(n9589), .Y(n13720) );
  NAND2X1 U24915 ( .A(n13698), .B(U1_A_i_d0[17]), .Y(n17207) );
  INVXL U24916 ( .A(n17207), .Y(n9592) );
  NAND2XL U24917 ( .A(n13699), .B(U1_A_i_d0[18]), .Y(n17204) );
  INVXL U24918 ( .A(n17204), .Y(n9591) );
  AOI21X1 U24919 ( .A0(n7001), .A1(n9592), .B0(n9591), .Y(n13723) );
  NAND2X1 U24920 ( .A(n13702), .B(U1_A_i_d0[19]), .Y(n17198) );
  INVXL U24921 ( .A(n17198), .Y(n9594) );
  NAND2XL U24922 ( .A(n7696), .B(U1_A_i_d0[20]), .Y(n13727) );
  INVXL U24923 ( .A(n13727), .Y(n9593) );
  AOI21X2 U24924 ( .A0(n13720), .A1(n9598), .B0(n9597), .Y(n9599) );
  OAI21X4 U24925 ( .A0(n13719), .A1(n9600), .B0(n9599), .Y(n17180) );
  INVX1 U24926 ( .A(n17189), .Y(n17195) );
  OR2X2 U24927 ( .A(n13710), .B(U1_A_i_d0[22]), .Y(n17191) );
  NOR2X1 U24928 ( .A(n13713), .B(U1_A_i_d0[23]), .Y(n17183) );
  NOR2XL U24929 ( .A(n17182), .B(n17183), .Y(n9604) );
  NAND2X1 U24930 ( .A(n13709), .B(U1_A_i_d0[21]), .Y(n17194) );
  NAND2XL U24931 ( .A(n13710), .B(U1_A_i_d0[22]), .Y(n17190) );
  INVXL U24932 ( .A(n17190), .Y(n9601) );
  NAND2X1 U24933 ( .A(n13716), .B(U1_A_i_d0[24]), .Y(n17177) );
  OR2X2 U24934 ( .A(n13717), .B(U1_A_i_d0[25]), .Y(n17175) );
  NAND2XL U24935 ( .A(n13717), .B(U1_A_i_d0[25]), .Y(n17174) );
  INVXL U24936 ( .A(n17174), .Y(n9605) );
  INVX4 U24937 ( .A(n7096), .Y(n17187) );
  OAI21XL U24938 ( .A0(n28710), .A1(n11430), .B0(n9609), .Y(U2_B_r[22]) );
  NAND2X1 U24939 ( .A(n11418), .B(BOPA[8]), .Y(n9610) );
  NAND2XL U24940 ( .A(BOPA[6]), .B(n11430), .Y(n9612) );
  NAND2XL U24941 ( .A(BOPA[8]), .B(n11430), .Y(n9613) );
  OAI21XL U24942 ( .A0(n6910), .A1(n11430), .B0(n9613), .Y(U2_B_r[8]) );
  NAND2XL U24943 ( .A(BOPA[9]), .B(n11430), .Y(n9614) );
  NAND2X1 U24944 ( .A(n11418), .B(BOPA[5]), .Y(n9616) );
  NAND2XL U24945 ( .A(BOPA[5]), .B(n11428), .Y(n9617) );
  OAI21XL U24946 ( .A0(n29105), .A1(n11428), .B0(n9617), .Y(U2_B_r[5]) );
  NOR2X2 U24947 ( .A(n9629), .B(U2_B_r[9]), .Y(n11562) );
  NOR2X2 U24948 ( .A(n11568), .B(n11562), .Y(n9631) );
  NOR2X2 U24949 ( .A(n9623), .B(n7088), .Y(n11586) );
  NOR2X1 U24950 ( .A(n11586), .B(n11584), .Y(n9625) );
  OAI21X1 U24951 ( .A0(n11586), .A1(n11583), .B0(n11587), .Y(n9624) );
  NAND2X2 U24952 ( .A(n9627), .B(U2_B_r[7]), .Y(n11575) );
  NAND2X1 U24953 ( .A(n9628), .B(n7130), .Y(n11569) );
  NAND2XL U24954 ( .A(n9629), .B(U2_B_r[9]), .Y(n11563) );
  AOI21X2 U24955 ( .A0(n11558), .A1(n9631), .B0(n9630), .Y(n9632) );
  OAI21X4 U24956 ( .A0(n9633), .A1(n11557), .B0(n9632), .Y(n11436) );
  CLKINVX3 U24957 ( .A(U2_B_i[10]), .Y(n9635) );
  NAND2X2 U24958 ( .A(n8147), .B(n11553), .Y(n11543) );
  INVXL U24959 ( .A(n11543), .Y(n9634) );
  NAND2XL U24960 ( .A(n9634), .B(n11545), .Y(n9641) );
  NAND2X1 U24961 ( .A(n9635), .B(U2_B_r[10]), .Y(n11552) );
  AOI21X2 U24962 ( .A0(n8147), .A1(n9637), .B0(n9636), .Y(n11542) );
  INVXL U24963 ( .A(n11542), .Y(n9639) );
  OAI21X1 U24964 ( .A0(n11555), .A1(n9641), .B0(n9640), .Y(n9644) );
  NOR2BX1 U24965 ( .AN(U2_B_r[13]), .B(U2_B_i[13]), .Y(n11431) );
  INVX4 U24966 ( .A(n9645), .Y(n11348) );
  NOR2XL U24967 ( .A(n9665), .B(U1_A_r_d0[6]), .Y(n9667) );
  NOR2XL U24968 ( .A(n9664), .B(U1_A_r_d0[5]), .Y(n19193) );
  NOR2XL U24969 ( .A(n9667), .B(n19193), .Y(n19188) );
  OR2X2 U24970 ( .A(n9668), .B(U1_A_r_d0[7]), .Y(n9670) );
  NAND2XL U24971 ( .A(n19188), .B(n9670), .Y(n9672) );
  NOR2XL U24972 ( .A(n9659), .B(U1_A_r_d0[4]), .Y(n9661) );
  NOR2XL U24973 ( .A(n9658), .B(U1_A_r_d0[3]), .Y(n19209) );
  NOR2XL U24974 ( .A(n9661), .B(n19209), .Y(n9663) );
  NOR2XL U24975 ( .A(n9397), .B(U1_A_r_d0[1]), .Y(n9651) );
  INVXL U24976 ( .A(n9651), .Y(n9653) );
  AOI21XL U24977 ( .A0(n9654), .A1(n9653), .B0(n9652), .Y(n19224) );
  OAI21XL U24978 ( .A0(n19224), .A1(n9657), .B0(n9656), .Y(n19207) );
  NAND2XL U24979 ( .A(n9659), .B(U1_A_r_d0[4]), .Y(n9660) );
  OAI21XL U24980 ( .A0(n9661), .A1(n19208), .B0(n9660), .Y(n9662) );
  AOI21XL U24981 ( .A0(n9663), .A1(n19207), .B0(n9662), .Y(n19186) );
  NAND2XL U24982 ( .A(n9664), .B(U1_A_r_d0[5]), .Y(n19194) );
  OAI21XL U24983 ( .A0(n9667), .A1(n19194), .B0(n9666), .Y(n19187) );
  AOI21XL U24984 ( .A0(n19187), .A1(n9670), .B0(n9669), .Y(n9671) );
  NOR2XL U24985 ( .A(n9674), .B(U1_A_r_d0[8]), .Y(n19167) );
  INVXL U24986 ( .A(n19167), .Y(n9673) );
  NAND2XL U24987 ( .A(n9679), .B(n9673), .Y(n19154) );
  OR2X2 U24988 ( .A(n9680), .B(U1_A_r_d0[11]), .Y(n19156) );
  NAND2XL U24989 ( .A(n9674), .B(U1_A_r_d0[8]), .Y(n19166) );
  INVXL U24990 ( .A(n19166), .Y(n9678) );
  NAND2XL U24991 ( .A(n9449), .B(U1_A_r_d0[9]), .Y(n19169) );
  NAND2XL U24992 ( .A(n9450), .B(U1_A_r_d0[10]), .Y(n9675) );
  OAI21XL U24993 ( .A0(n9676), .A1(n19169), .B0(n9675), .Y(n9677) );
  NOR2XL U24994 ( .A(n9693), .B(U1_A_r_d0[15]), .Y(n19132) );
  OR2X2 U24995 ( .A(n9690), .B(U1_A_r_d0[13]), .Y(n19143) );
  NAND2XL U24996 ( .A(n9692), .B(n19143), .Y(n19127) );
  NOR2X1 U24997 ( .A(n9707), .B(n19105), .Y(n9709) );
  AND2X2 U24998 ( .A(n9690), .B(U1_A_r_d0[13]), .Y(n19142) );
  AOI21XL U24999 ( .A0(n9692), .A1(n19142), .B0(n9691), .Y(n19128) );
  NAND2XL U25000 ( .A(n9693), .B(U1_A_r_d0[15]), .Y(n19131) );
  INVXL U25001 ( .A(n19131), .Y(n9696) );
  AND2X2 U25002 ( .A(n9694), .B(U1_A_r_d0[16]), .Y(n9695) );
  AND2X2 U25003 ( .A(n9701), .B(U1_A_r_d0[18]), .Y(n9702) );
  AND2X2 U25004 ( .A(n9703), .B(U1_A_r_d0[20]), .Y(n9704) );
  AOI21X2 U25005 ( .A0(n19102), .A1(n9709), .B0(n9708), .Y(n9710) );
  NOR2X1 U25006 ( .A(n5848), .B(U1_A_r_d0[21]), .Y(n19092) );
  NOR2XL U25007 ( .A(n9712), .B(U1_A_r_d0[22]), .Y(n9714) );
  NAND2XL U25008 ( .A(n19081), .B(n9716), .Y(n19074) );
  NOR2X1 U25009 ( .A(n9717), .B(U1_A_r_d0[24]), .Y(n9719) );
  NAND2X1 U25010 ( .A(n5848), .B(U1_A_r_d0[21]), .Y(n19091) );
  NAND2XL U25011 ( .A(n9712), .B(U1_A_r_d0[22]), .Y(n9713) );
  AOI21X1 U25012 ( .A0(n19082), .A1(n9716), .B0(n9715), .Y(n19073) );
  NAND2XL U25013 ( .A(n9717), .B(U1_A_r_d0[24]), .Y(n9718) );
  NOR2XL U25014 ( .A(n9720), .B(U1_A_r_d0[25]), .Y(n9722) );
  NAND2XL U25015 ( .A(n9720), .B(U1_A_r_d0[25]), .Y(n9721) );
  MXI2X1 U25016 ( .A(U1_pipe2[27]), .B(n9724), .S0(n5812), .Y(n5039) );
  NOR2X2 U25017 ( .A(n9974), .B(n9972), .Y(n9967) );
  NAND2X1 U25018 ( .A(W1[7]), .B(W1[23]), .Y(n9969) );
  NAND2X1 U25019 ( .A(W1[8]), .B(W1[24]), .Y(n9980) );
  OAI21X2 U25020 ( .A0(n9963), .A1(n9980), .B0(n9964), .Y(n9956) );
  NOR2X1 U25021 ( .A(W1[12]), .B(W1[28]), .Y(n9952) );
  NOR2XL U25022 ( .A(n9948), .B(n9952), .Y(n9992) );
  INVXL U25023 ( .A(n9992), .Y(n9729) );
  NAND2X1 U25024 ( .A(W1[12]), .B(W1[28]), .Y(n9953) );
  NAND2XL U25025 ( .A(W1[13]), .B(W1[29]), .Y(n9949) );
  OAI21XL U25026 ( .A0(n9948), .A1(n9953), .B0(n9949), .Y(n9996) );
  INVXL U25027 ( .A(n9996), .Y(n9728) );
  OAI21X1 U25028 ( .A0(n9955), .A1(n9729), .B0(n9728), .Y(n9732) );
  NOR2XL U25029 ( .A(W1[14]), .B(W1[30]), .Y(n9730) );
  INVXL U25030 ( .A(n9730), .Y(n9995) );
  NAND2XL U25031 ( .A(W1[14]), .B(W1[30]), .Y(n9993) );
  NAND2X1 U25032 ( .A(n9995), .B(n9993), .Y(n9731) );
  MXI2X1 U25033 ( .A(U1_pipe10[26]), .B(n9733), .S0(n17641), .Y(n4864) );
  NAND2X1 U25034 ( .A(W3[3]), .B(W3[19]), .Y(n9765) );
  NAND2X1 U25035 ( .A(W3[6]), .B(W3[22]), .Y(n9800) );
  NOR2XL U25036 ( .A(n9786), .B(n9784), .Y(n9768) );
  NAND2XL U25037 ( .A(n9768), .B(n9735), .Y(n9752) );
  INVXL U25038 ( .A(n9752), .Y(n9737) );
  NAND2XL U25039 ( .A(W3[8]), .B(W3[24]), .Y(n9797) );
  NAND2XL U25040 ( .A(W3[10]), .B(W3[26]), .Y(n9790) );
  NAND2X1 U25041 ( .A(W3[11]), .B(W3[27]), .Y(n9770) );
  OAI21XL U25042 ( .A0(n9769), .A1(n9790), .B0(n9770), .Y(n9734) );
  INVXL U25043 ( .A(n9758), .Y(n9736) );
  INVXL U25044 ( .A(n9755), .Y(n9738) );
  OAI21XL U25045 ( .A0(n9806), .A1(n9739), .B0(n9738), .Y(n9741) );
  XNOR2X1 U25046 ( .A(n9741), .B(n10034), .Y(U2_U0_z2[14]) );
  AOI21X1 U25047 ( .A0(n9755), .A1(n9740), .B0(n9754), .Y(n9756) );
  INVXL U25048 ( .A(n9761), .Y(n9773) );
  CLKINVX3 U25049 ( .A(n9762), .Y(U2_U0_z2[16]) );
  INVXL U25050 ( .A(n9769), .Y(n9771) );
  XNOR2X2 U25051 ( .A(n9772), .B(n10078), .Y(U2_U0_z2[11]) );
  ADDFX2 U25052 ( .A(n8000), .B(n7986), .CI(n9773), .CO(n9762), .S(
        U2_U0_z2[15]) );
  XOR2X1 U25053 ( .A(n10048), .B(n9777), .Y(U2_U0_z2[1]) );
  INVXL U25054 ( .A(n9786), .Y(n9788) );
  INVXL U25055 ( .A(n9789), .Y(n9791) );
  XOR2X1 U25056 ( .A(n9802), .B(n10104), .Y(U2_U0_z2[6]) );
  XNOR2X1 U25057 ( .A(n9809), .B(n10087), .Y(U2_U0_z2[4]) );
  NOR2XL U25058 ( .A(n9820), .B(n9859), .Y(n9863) );
  INVXL U25059 ( .A(n9863), .Y(n9817) );
  NAND2X1 U25060 ( .A(W0[13]), .B(W0[29]), .Y(n9821) );
  INVXL U25061 ( .A(n9867), .Y(n9816) );
  OAI21X1 U25062 ( .A0(n9862), .A1(n9817), .B0(n9816), .Y(n9819) );
  NOR2XL U25063 ( .A(W0[14]), .B(W0[30]), .Y(n9818) );
  OAI21X2 U25064 ( .A0(n9862), .A1(n9859), .B0(n9860), .Y(n9823) );
  XNOR2X4 U25065 ( .A(n9823), .B(n10173), .Y(U0_U0_z2[13]) );
  INVXL U25066 ( .A(n9833), .Y(n9835) );
  XOR2X2 U25067 ( .A(n9836), .B(n10168), .Y(U0_U0_z2[6]) );
  AOI21X2 U25068 ( .A0(n9844), .A1(n9843), .B0(n9838), .Y(n9841) );
  XOR2X4 U25069 ( .A(n9841), .B(n10150), .Y(U0_U0_z2[5]) );
  OAI21XL U25070 ( .A0(n9853), .A1(n9850), .B0(n9851), .Y(n9849) );
  XNOR2X2 U25071 ( .A(n9849), .B(n10156), .Y(U0_U0_z2[3]) );
  XOR2X1 U25072 ( .A(n9853), .B(n10191), .Y(U0_U0_z2[2]) );
  NAND2XL U25073 ( .A(n9855), .B(n9854), .Y(n10164) );
  XNOR2X1 U25074 ( .A(n9870), .B(n10164), .Y(U0_U0_z2[8]) );
  XOR2X1 U25075 ( .A(n9862), .B(n10166), .Y(U0_U0_z2[12]) );
  ADDFHX4 U25076 ( .A(n8006), .B(n7987), .CI(n9872), .CO(n9873), .S(
        U0_U0_z2[15]) );
  NOR2X4 U25077 ( .A(W2[5]), .B(W2[21]), .Y(n9907) );
  NOR2X2 U25078 ( .A(W2[7]), .B(W2[23]), .Y(n9897) );
  OAI21XL U25079 ( .A0(n9886), .A1(n9939), .B0(n9887), .Y(n9874) );
  NOR2XL U25080 ( .A(n9881), .B(n9941), .Y(n9919) );
  INVXL U25081 ( .A(n9919), .Y(n9879) );
  INVXL U25082 ( .A(n9924), .Y(n9878) );
  OAI21X1 U25083 ( .A0(n9944), .A1(n9879), .B0(n9878), .Y(n9880) );
  OR2X2 U25084 ( .A(W2[14]), .B(W2[30]), .Y(n9923) );
  NAND2XL U25085 ( .A(W2[14]), .B(W2[30]), .Y(n9921) );
  NAND2X1 U25086 ( .A(n9923), .B(n9921), .Y(n10292) );
  XNOR2X2 U25087 ( .A(n9880), .B(n10292), .Y(U1_U2_z2[14]) );
  INVXL U25088 ( .A(n9881), .Y(n9883) );
  AOI21X2 U25089 ( .A0(n9934), .A1(n9933), .B0(n9891), .Y(n9895) );
  XNOR2X4 U25090 ( .A(n9900), .B(n7129), .Y(U1_U2_z2[7]) );
  XOR2X1 U25091 ( .A(n9904), .B(n10337), .Y(U1_U2_z2[6]) );
  INVXL U25092 ( .A(n9911), .Y(n9906) );
  AOI21XL U25093 ( .A0(n9913), .A1(n9912), .B0(n9906), .Y(n9910) );
  XOR2X2 U25094 ( .A(n9910), .B(n10319), .Y(U1_U2_z2[5]) );
  XNOR2X1 U25095 ( .A(n9913), .B(n10322), .Y(U1_U2_z2[4]) );
  OAI21XL U25096 ( .A0(n9947), .A1(n9945), .B0(n9946), .Y(n9918) );
  NAND2X1 U25097 ( .A(n9917), .B(n9916), .Y(n10342) );
  XNOR2X2 U25098 ( .A(n9918), .B(n10342), .Y(U1_U2_z2[3]) );
  NAND2XL U25099 ( .A(n9919), .B(n9923), .Y(n9926) );
  NOR2XL U25100 ( .A(n9920), .B(n9926), .Y(n9930) );
  INVXL U25101 ( .A(n9921), .Y(n9922) );
  OAI21XL U25102 ( .A0(n9927), .A1(n9926), .B0(n9925), .Y(n9928) );
  INVXL U25103 ( .A(n9928), .Y(n9929) );
  XNOR2X1 U25104 ( .A(n9934), .B(n10329), .Y(U1_U2_z2[8]) );
  INVXL U25105 ( .A(n9941), .Y(n9943) );
  XOR2X1 U25106 ( .A(n9947), .B(n10345), .Y(U1_U2_z2[2]) );
  OAI21X2 U25107 ( .A0(n9955), .A1(n9952), .B0(n9953), .Y(n9951) );
  INVXL U25108 ( .A(n9948), .Y(n9950) );
  XOR2X1 U25109 ( .A(n9955), .B(n10244), .Y(U1_U1_z2[12]) );
  XNOR2X4 U25110 ( .A(n9960), .B(n10220), .Y(U1_U1_z2[11]) );
  OAI21X2 U25111 ( .A0(n9985), .A1(n9982), .B0(n9983), .Y(n9971) );
  XNOR2X4 U25112 ( .A(n9971), .B(n10234), .Y(U1_U1_z2[7]) );
  XNOR2X1 U25113 ( .A(n9991), .B(n10238), .Y(U1_U1_z2[4]) );
  INVXL U25114 ( .A(n9993), .Y(n9994) );
  AOI21XL U25115 ( .A0(n9996), .A1(n9995), .B0(n9994), .Y(n9997) );
  INVX8 U25116 ( .A(n10001), .Y(U1_U1_z2[16]) );
  INVX1 U25117 ( .A(n10002), .Y(n10004) );
  XOR2X2 U25118 ( .A(n12004), .B(n10005), .Y(U1_U1_z2[1]) );
  XOR2X1 U25119 ( .A(n10009), .B(n10264), .Y(U1_U1_z2[2]) );
  NOR2X2 U25120 ( .A(n8019), .B(W3[16]), .Y(n10049) );
  OAI21X2 U25121 ( .A0(n10011), .A1(n10049), .B0(n10010), .Y(n10070) );
  NOR2X2 U25122 ( .A(n8021), .B(W3[19]), .Y(n10013) );
  NOR2X1 U25123 ( .A(n10013), .B(n10072), .Y(n10015) );
  OAI21X2 U25124 ( .A0(n10013), .A1(n10071), .B0(n10012), .Y(n10014) );
  AOI21X4 U25125 ( .A0(n10070), .A1(n10015), .B0(n10014), .Y(n10041) );
  NOR2X1 U25126 ( .A(n8037), .B(W3[22]), .Y(n10045) );
  NAND2X1 U25127 ( .A(n8022), .B(W3[21]), .Y(n10016) );
  OAI21X1 U25128 ( .A0(n10017), .A1(n10059), .B0(n10016), .Y(n10042) );
  NAND2XL U25129 ( .A(n8015), .B(W3[23]), .Y(n10018) );
  OAI21X4 U25130 ( .A0(n10041), .A1(n10021), .B0(n10020), .Y(n10103) );
  NOR2XL U25131 ( .A(n8023), .B(W3[24]), .Y(n10051) );
  NOR2XL U25132 ( .A(n8018), .B(W3[27]), .Y(n10025) );
  NOR2XL U25133 ( .A(n10025), .B(n10077), .Y(n10027) );
  NAND2XL U25134 ( .A(n10038), .B(n10027), .Y(n10092) );
  INVXL U25135 ( .A(n10092), .Y(n10029) );
  OAI21X1 U25136 ( .A0(n10023), .A1(n10052), .B0(n10022), .Y(n10037) );
  NAND2XL U25137 ( .A(n7985), .B(W3[26]), .Y(n10076) );
  OAI21XL U25138 ( .A0(n10025), .A1(n10076), .B0(n10024), .Y(n10026) );
  AOI21X1 U25139 ( .A0(n10037), .A1(n10027), .B0(n10026), .Y(n10097) );
  INVXL U25140 ( .A(n10097), .Y(n10028) );
  AOI21X2 U25141 ( .A0(n10103), .A1(n10029), .B0(n10028), .Y(n10083) );
  NOR2XL U25142 ( .A(n8016), .B(W3[29]), .Y(n10031) );
  NOR2XL U25143 ( .A(n7984), .B(W3[28]), .Y(n10066) );
  NOR2XL U25144 ( .A(n10031), .B(n10066), .Y(n10091) );
  NAND2XL U25145 ( .A(n7984), .B(W3[28]), .Y(n10065) );
  OAI21XL U25146 ( .A0(n10031), .A1(n10065), .B0(n10030), .Y(n10094) );
  XNOR2X1 U25147 ( .A(n10036), .B(n10035), .Y(U2_U0_z1[14]) );
  CLKINVX2 U25148 ( .A(n10041), .Y(n10089) );
  OAI21X1 U25149 ( .A0(n10106), .A1(n10045), .B0(n10044), .Y(n10047) );
  AOI21XL U25150 ( .A0(n10103), .A1(n10054), .B0(n10053), .Y(n10057) );
  INVXL U25151 ( .A(n10058), .Y(n10061) );
  INVXL U25152 ( .A(n10059), .Y(n10060) );
  AOI21XL U25153 ( .A0(n10089), .A1(n10061), .B0(n10060), .Y(n10064) );
  XOR2X2 U25154 ( .A(n10064), .B(n10063), .Y(U2_U0_z1[5]) );
  XNOR2X2 U25155 ( .A(n10069), .B(n10068), .Y(U2_U0_z1[13]) );
  XNOR2X2 U25156 ( .A(n10075), .B(n10074), .Y(U2_U0_z1[3]) );
  XNOR2X2 U25157 ( .A(n10080), .B(n10079), .Y(U2_U0_z1[11]) );
  INVX1 U25158 ( .A(n10081), .Y(n10082) );
  NOR2X1 U25159 ( .A(n7982), .B(W3[30]), .Y(n10090) );
  NOR2XL U25160 ( .A(n10092), .B(n10096), .Y(n10099) );
  AOI21XL U25161 ( .A0(n10094), .A1(n10093), .B0(n7983), .Y(n10095) );
  CLKINVX3 U25162 ( .A(n10101), .Y(U2_U0_z1[16]) );
  XOR2X1 U25163 ( .A(n10106), .B(n10105), .Y(U2_U0_z1[6]) );
  XNOR2XL U25164 ( .A(n8019), .B(W3[16]), .Y(U2_U0_z1[0]) );
  NOR2X2 U25165 ( .A(n10108), .B(n10155), .Y(n10110) );
  NAND2X1 U25166 ( .A(n8026), .B(W0[19]), .Y(n10107) );
  OAI21X2 U25167 ( .A0(n10108), .A1(n10154), .B0(n10107), .Y(n10109) );
  NOR2X4 U25168 ( .A(n10114), .B(n10143), .Y(n10116) );
  NAND2X2 U25169 ( .A(n8039), .B(W0[22]), .Y(n10142) );
  NAND2X1 U25170 ( .A(n8043), .B(W0[23]), .Y(n10113) );
  NOR2X1 U25171 ( .A(n7998), .B(W0[24]), .Y(n10133) );
  NOR2X2 U25172 ( .A(n10117), .B(n10133), .Y(n10129) );
  NAND2XL U25173 ( .A(n8025), .B(W0[27]), .Y(n10118) );
  NOR2XL U25174 ( .A(n8005), .B(W0[29]), .Y(n10123) );
  NAND2X1 U25175 ( .A(n7973), .B(W0[28]), .Y(n10171) );
  NAND2XL U25176 ( .A(n8005), .B(W0[29]), .Y(n10122) );
  INVXL U25177 ( .A(n10182), .Y(n10124) );
  XNOR2X4 U25178 ( .A(n10132), .B(n5763), .Y(U0_U0_z1[11]) );
  INVXL U25179 ( .A(n10133), .Y(n10136) );
  INVX4 U25180 ( .A(n10139), .Y(n10190) );
  AOI21X4 U25181 ( .A0(n10190), .A1(n10141), .B0(n10140), .Y(n10170) );
  OAI21X4 U25182 ( .A0(n10170), .A1(n10143), .B0(n10142), .Y(n10145) );
  XNOR2X4 U25183 ( .A(n10145), .B(n10144), .Y(U0_U0_z1[7]) );
  INVXL U25184 ( .A(n12002), .Y(n10163) );
  XOR2X4 U25185 ( .A(n10174), .B(n10173), .Y(U0_U0_z1[13]) );
  INVX1 U25186 ( .A(n10175), .Y(n10176) );
  NOR2XL U25187 ( .A(n7975), .B(W0[30]), .Y(n10178) );
  INVXL U25188 ( .A(n10178), .Y(n10181) );
  NOR2XL U25189 ( .A(n10180), .B(n10184), .Y(n10186) );
  AOI21X1 U25190 ( .A0(n10182), .A1(n10181), .B0(n7981), .Y(n10183) );
  INVX8 U25191 ( .A(n10187), .Y(U0_U0_z1[16]) );
  XOR2X1 U25192 ( .A(n10193), .B(n10192), .Y(U0_U0_z1[2]) );
  NOR2X1 U25193 ( .A(n8017), .B(W1[24]), .Y(n10223) );
  NOR2X1 U25194 ( .A(n8024), .B(W1[27]), .Y(n10202) );
  NOR2XL U25195 ( .A(n10205), .B(n10214), .Y(n10247) );
  OR2X2 U25196 ( .A(n8004), .B(W1[30]), .Y(n10252) );
  NAND2XL U25197 ( .A(n8024), .B(W1[27]), .Y(n10201) );
  NAND2XL U25198 ( .A(n8007), .B(W1[29]), .Y(n10204) );
  OAI21XL U25199 ( .A0(n10205), .A1(n10213), .B0(n10204), .Y(n10248) );
  AOI21XL U25200 ( .A0(n10248), .A1(n10252), .B0(n10206), .Y(n10207) );
  XNOR2X4 U25201 ( .A(n10222), .B(n10221), .Y(U1_U1_z1[11]) );
  XNOR2X1 U25202 ( .A(n10260), .B(n10239), .Y(U1_U1_z1[4]) );
  XNOR2X2 U25203 ( .A(n10243), .B(n10242), .Y(U1_U1_z1[3]) );
  INVXL U25204 ( .A(n10247), .Y(n10250) );
  INVXL U25205 ( .A(n10248), .Y(n10249) );
  NAND2X1 U25206 ( .A(n10252), .B(n10251), .Y(n10253) );
  XNOR2X2 U25207 ( .A(n10254), .B(n10253), .Y(U1_U1_z1[14]) );
  XNOR2X1 U25208 ( .A(n8009), .B(W1[16]), .Y(U1_U1_z1[0]) );
  NOR2X1 U25209 ( .A(n8011), .B(W2[24]), .Y(n10303) );
  NAND2XL U25210 ( .A(n10299), .B(n10274), .Y(n10284) );
  OR2X2 U25211 ( .A(n8012), .B(W2[30]), .Y(n10277) );
  NOR2XL U25212 ( .A(n10284), .B(n10279), .Y(n10281) );
  NAND2XL U25213 ( .A(n7997), .B(W2[27]), .Y(n10271) );
  OAI21XL U25214 ( .A0(n10272), .A1(n10300), .B0(n10271), .Y(n10273) );
  INVXL U25215 ( .A(n10326), .Y(n10282) );
  NAND2X1 U25216 ( .A(W2[15]), .B(n7978), .Y(n10325) );
  NAND2XL U25217 ( .A(n10282), .B(n10325), .Y(n10283) );
  INVXL U25218 ( .A(n10288), .Y(n10291) );
  XNOR2X4 U25219 ( .A(n10297), .B(n5759), .Y(U1_U2_z1[13]) );
  XNOR2X4 U25220 ( .A(n10302), .B(n5769), .Y(U1_U2_z1[11]) );
  INVXL U25221 ( .A(n10303), .Y(n10306) );
  XNOR2X4 U25222 ( .A(n10314), .B(n6891), .Y(U1_U2_z1[7]) );
  AOI21X1 U25223 ( .A0(n10324), .A1(n10318), .B0(n10317), .Y(n10321) );
  INVX1 U25224 ( .A(n10319), .Y(n10320) );
  XOR2X1 U25225 ( .A(n10336), .B(n10335), .Y(U1_U2_z1[12]) );
  INVX1 U25226 ( .A(n10339), .Y(n10347) );
  OAI21XL U25227 ( .A0(n10347), .A1(n10341), .B0(n10340), .Y(n10344) );
  INVX1 U25228 ( .A(n10342), .Y(n10343) );
  XNOR2X2 U25229 ( .A(n10344), .B(n10343), .Y(U1_U2_z1[3]) );
  INVXL U25230 ( .A(n10345), .Y(n10346) );
  XOR2X1 U25231 ( .A(n10347), .B(n10346), .Y(U1_U2_z1[2]) );
  XNOR2X1 U25232 ( .A(n8008), .B(W2[16]), .Y(U1_U2_z1[0]) );
  NAND2XL U25233 ( .A(n10513), .B(n10349), .Y(n10351) );
  XNOR2X1 U25234 ( .A(n10354), .B(n10353), .Y(U0_U0_z0[25]) );
  INVXL U25235 ( .A(n10355), .Y(n10356) );
  NOR2XL U25236 ( .A(n10356), .B(n10359), .Y(n10362) );
  NAND2XL U25237 ( .A(n10362), .B(n10371), .Y(n10364) );
  INVXL U25238 ( .A(n10357), .Y(n10360) );
  OAI21XL U25239 ( .A0(n10360), .A1(n10359), .B0(n10358), .Y(n10361) );
  AOI21XL U25240 ( .A0(n10373), .A1(n10362), .B0(n10361), .Y(n10363) );
  INVXL U25241 ( .A(n10365), .Y(n10367) );
  NAND2XL U25242 ( .A(n10371), .B(n10384), .Y(n10375) );
  OAI21X2 U25243 ( .A0(n10522), .A1(n10375), .B0(n10374), .Y(n10380) );
  NAND2X1 U25244 ( .A(n10378), .B(n10377), .Y(n10379) );
  OAI21X4 U25245 ( .A0(n10522), .A1(n10382), .B0(n10381), .Y(n10386) );
  NAND2X1 U25246 ( .A(n10384), .B(n10383), .Y(n10385) );
  XNOR2X4 U25247 ( .A(n10386), .B(n10385), .Y(U0_U0_z0[20]) );
  INVXL U25248 ( .A(n10400), .Y(n10388) );
  OAI21X4 U25249 ( .A0(n10522), .A1(n10390), .B0(n10389), .Y(n10395) );
  INVXL U25250 ( .A(n10391), .Y(n10393) );
  NAND2X1 U25251 ( .A(n10393), .B(n10392), .Y(n10394) );
  XNOR2X4 U25252 ( .A(n10395), .B(n10394), .Y(U0_U0_z0[19]) );
  NAND2XL U25253 ( .A(n10411), .B(n10410), .Y(n10412) );
  XOR2X1 U25254 ( .A(n10413), .B(n10412), .Y(U0_U0_z0[16]) );
  INVXL U25255 ( .A(n10427), .Y(n10415) );
  NOR2XL U25256 ( .A(n10415), .B(n10430), .Y(n10418) );
  INVXL U25257 ( .A(n10447), .Y(n10436) );
  INVXL U25258 ( .A(n10426), .Y(n10416) );
  OAI21XL U25259 ( .A0(n10416), .A1(n10430), .B0(n10431), .Y(n10417) );
  AOI21X1 U25260 ( .A0(n10438), .A1(n10418), .B0(n10417), .Y(n10419) );
  INVXL U25261 ( .A(n10421), .Y(n10423) );
  NAND2XL U25262 ( .A(n10436), .B(n10427), .Y(n10429) );
  INVXL U25263 ( .A(n10430), .Y(n10432) );
  XNOR2X2 U25264 ( .A(n10434), .B(n10433), .Y(U0_U0_z0[14]) );
  NAND2XL U25265 ( .A(n10436), .B(n10449), .Y(n10440) );
  XNOR2X2 U25266 ( .A(n10445), .B(n10444), .Y(U0_U0_z0[13]) );
  XNOR2X2 U25267 ( .A(n10451), .B(n10450), .Y(U0_U0_z0[12]) );
  AOI21XL U25268 ( .A0(n10462), .A1(n10466), .B0(n10453), .Y(n10454) );
  OAI21X1 U25269 ( .A0(n10477), .A1(n10455), .B0(n10454), .Y(n10460) );
  XNOR2X1 U25270 ( .A(n10460), .B(n10459), .Y(U0_U0_z0[11]) );
  NAND2X1 U25271 ( .A(n10471), .B(n10470), .Y(n10472) );
  INVXL U25272 ( .A(n10481), .Y(n10483) );
  INVXL U25273 ( .A(n10485), .Y(n10487) );
  INVXL U25274 ( .A(n10490), .Y(n10498) );
  INVXL U25275 ( .A(n10497), .Y(n10491) );
  AOI21X1 U25276 ( .A0(n10500), .A1(n10498), .B0(n10491), .Y(n10496) );
  NAND2XL U25277 ( .A(n10494), .B(n10493), .Y(n10495) );
  XOR2X1 U25278 ( .A(n10496), .B(n10495), .Y(U0_U0_z0[5]) );
  NAND2XL U25279 ( .A(n10498), .B(n10497), .Y(n10499) );
  XNOR2X1 U25280 ( .A(n10500), .B(n10499), .Y(U0_U0_z0[4]) );
  OAI21XL U25281 ( .A0(n10511), .A1(n10507), .B0(n10508), .Y(n10506) );
  NAND2XL U25282 ( .A(n10504), .B(n10503), .Y(n10505) );
  XNOR2X1 U25283 ( .A(n10506), .B(n10505), .Y(U0_U0_z0[3]) );
  NOR2XL U25284 ( .A(n10516), .B(n10512), .Y(n10518) );
  NAND2XL U25285 ( .A(n10513), .B(n10518), .Y(n10521) );
  OAI21XL U25286 ( .A0(n10516), .A1(n10515), .B0(n10514), .Y(n10517) );
  OAI21XL U25287 ( .A0(n10522), .A1(n10521), .B0(n10520), .Y(n10523) );
  INVXL U25288 ( .A(n10523), .Y(U0_U0_z0[26]) );
  NAND2XL U25289 ( .A(n10526), .B(n10525), .Y(n10528) );
  NAND2XL U25290 ( .A(n10671), .B(n10530), .Y(n10532) );
  AOI21XL U25291 ( .A0(n10677), .A1(n10530), .B0(n10529), .Y(n10531) );
  OAI21X1 U25292 ( .A0(n6712), .A1(n10532), .B0(n10531), .Y(n10535) );
  INVXL U25293 ( .A(n10674), .Y(n10533) );
  INVXL U25294 ( .A(n10548), .Y(n10536) );
  NOR2XL U25295 ( .A(n10536), .B(n10550), .Y(n10539) );
  INVXL U25296 ( .A(n10565), .Y(n10554) );
  NAND2XL U25297 ( .A(n10539), .B(n10554), .Y(n10541) );
  INVXL U25298 ( .A(n10547), .Y(n10537) );
  OAI21XL U25299 ( .A0(n10537), .A1(n10550), .B0(n10551), .Y(n10538) );
  AOI21XL U25300 ( .A0(n10556), .A1(n10539), .B0(n10538), .Y(n10540) );
  INVXL U25301 ( .A(n10542), .Y(n10544) );
  NAND2XL U25302 ( .A(n10554), .B(n10548), .Y(n10549) );
  NAND2XL U25303 ( .A(n10554), .B(n10567), .Y(n10558) );
  AOI21XL U25304 ( .A0(n10556), .A1(n10567), .B0(n10555), .Y(n10557) );
  NAND2X1 U25305 ( .A(n10561), .B(n10560), .Y(n10562) );
  OAI21X1 U25306 ( .A0(n6712), .A1(n10565), .B0(n10564), .Y(n10569) );
  NAND2X1 U25307 ( .A(n10567), .B(n10566), .Y(n10568) );
  XNOR2X4 U25308 ( .A(n10569), .B(n10568), .Y(U1_U0_z0[20]) );
  NAND2X1 U25309 ( .A(n10576), .B(n10575), .Y(n10577) );
  XNOR2X4 U25310 ( .A(n10578), .B(n10577), .Y(U1_U0_z0[19]) );
  NAND2XL U25311 ( .A(n10594), .B(n10593), .Y(n10595) );
  XOR2X1 U25312 ( .A(n7148), .B(n10595), .Y(U1_U0_z0[16]) );
  NAND2XL U25313 ( .A(n10606), .B(n10597), .Y(n10599) );
  OAI21X1 U25314 ( .A0(n10643), .A1(n10599), .B0(n10598), .Y(n10604) );
  INVXL U25315 ( .A(n10600), .Y(n10602) );
  NAND2X1 U25316 ( .A(n10602), .B(n10601), .Y(n10603) );
  NAND2XL U25317 ( .A(n10606), .B(n10619), .Y(n10610) );
  NAND2XL U25318 ( .A(n10613), .B(n10612), .Y(n10614) );
  XNOR2X2 U25319 ( .A(n10615), .B(n10614), .Y(U1_U0_z0[13]) );
  INVXL U25320 ( .A(n10630), .Y(n10622) );
  XNOR2X2 U25321 ( .A(n10633), .B(n10632), .Y(U1_U0_z0[10]) );
  NAND2XL U25322 ( .A(n7223), .B(n6912), .Y(n10648) );
  XNOR2X1 U25323 ( .A(n10649), .B(n10648), .Y(U1_U0_z0[7]) );
  INVXL U25324 ( .A(n10650), .Y(n10652) );
  INVXL U25325 ( .A(n10654), .Y(n10662) );
  INVXL U25326 ( .A(n10661), .Y(n10655) );
  NAND2XL U25327 ( .A(n10658), .B(n10657), .Y(n10659) );
  XOR2X1 U25328 ( .A(n10660), .B(n10659), .Y(U1_U0_z0[5]) );
  OAI21XL U25329 ( .A0(n10690), .A1(n10686), .B0(n10687), .Y(n10669) );
  INVXL U25330 ( .A(n10665), .Y(n10667) );
  NAND2XL U25331 ( .A(n10667), .B(n10666), .Y(n10668) );
  NOR2XL U25332 ( .A(n10674), .B(n10670), .Y(n10676) );
  NAND2XL U25333 ( .A(n10671), .B(n10676), .Y(n10679) );
  OAI21XL U25334 ( .A0(n10674), .A1(n10673), .B0(n10672), .Y(n10675) );
  AOI21XL U25335 ( .A0(n10677), .A1(n10676), .B0(n10675), .Y(n10678) );
  OAI21XL U25336 ( .A0(n7148), .A1(n10679), .B0(n10678), .Y(n10680) );
  INVXL U25337 ( .A(n10680), .Y(U1_U0_z0[26]) );
  XNOR2X1 U25338 ( .A(n8193), .B(BOPB[26]), .Y(U1_U0_z0[0]) );
  NAND2XL U25339 ( .A(n10688), .B(n10687), .Y(n10689) );
  NOR2XL U25340 ( .A(n10726), .B(n10715), .Y(n10695) );
  NAND2XL U25341 ( .A(n10722), .B(n10695), .Y(n10697) );
  NOR2XL U25342 ( .A(n10697), .B(n10732), .Y(n10847) );
  NAND2XL U25343 ( .A(n10847), .B(n10706), .Y(n10700) );
  OAI21XL U25344 ( .A0(n10693), .A1(n10733), .B0(n10692), .Y(n10721) );
  NAND2XL U25345 ( .A(n8159), .B(BOPD[48]), .Y(n10727) );
  NAND2XL U25346 ( .A(n8155), .B(BOPD[49]), .Y(n10716) );
  OAI21XL U25347 ( .A0(n10715), .A1(n10727), .B0(n10716), .Y(n10694) );
  AOI21XL U25348 ( .A0(n10695), .A1(n10721), .B0(n10694), .Y(n10696) );
  OAI21XL U25349 ( .A0(n10731), .A1(n10697), .B0(n10696), .Y(n10853) );
  AOI21XL U25350 ( .A0(n10853), .A1(n10706), .B0(n10698), .Y(n10699) );
  INVXL U25351 ( .A(n10847), .Y(n10705) );
  INVXL U25352 ( .A(n10853), .Y(n10704) );
  NAND2X1 U25353 ( .A(n10706), .B(n10849), .Y(n10707) );
  INVXL U25354 ( .A(n10722), .Y(n10709) );
  NOR2XL U25355 ( .A(n10709), .B(n10726), .Y(n10712) );
  NAND2XL U25356 ( .A(n10712), .B(n10720), .Y(n10714) );
  INVXL U25357 ( .A(n10721), .Y(n10710) );
  OAI21XL U25358 ( .A0(n10710), .A1(n10726), .B0(n10727), .Y(n10711) );
  AOI21XL U25359 ( .A0(n10723), .A1(n10712), .B0(n10711), .Y(n10713) );
  INVXL U25360 ( .A(n10715), .Y(n10717) );
  NAND2XL U25361 ( .A(n10720), .B(n10722), .Y(n10725) );
  AOI21XL U25362 ( .A0(n10723), .A1(n10722), .B0(n10721), .Y(n10724) );
  INVXL U25363 ( .A(n10726), .Y(n10728) );
  NAND2X1 U25364 ( .A(n10734), .B(n10733), .Y(n10735) );
  NAND2X1 U25365 ( .A(n10743), .B(n10742), .Y(n10744) );
  NAND2X1 U25366 ( .A(n10751), .B(n10750), .Y(n10752) );
  XNOR2X2 U25367 ( .A(n10760), .B(n10759), .Y(U1_U2_z0[17]) );
  INVXL U25368 ( .A(n10773), .Y(n10762) );
  NOR2XL U25369 ( .A(n10762), .B(n10776), .Y(n10765) );
  INVX1 U25370 ( .A(n10790), .Y(n10780) );
  NAND2X1 U25371 ( .A(n10765), .B(n10780), .Y(n10767) );
  INVX2 U25372 ( .A(n10789), .Y(n10782) );
  INVXL U25373 ( .A(n10772), .Y(n10763) );
  OAI21XL U25374 ( .A0(n10763), .A1(n10776), .B0(n10777), .Y(n10764) );
  AOI21X2 U25375 ( .A0(n10782), .A1(n10765), .B0(n10764), .Y(n10766) );
  NAND2XL U25376 ( .A(n7386), .B(n10769), .Y(n10770) );
  NAND2XL U25377 ( .A(n10780), .B(n10773), .Y(n10775) );
  AOI21XL U25378 ( .A0(n10773), .A1(n10782), .B0(n10772), .Y(n10774) );
  OAI21X1 U25379 ( .A0(n10817), .A1(n10775), .B0(n10774), .Y(n10778) );
  NAND2XL U25380 ( .A(n10780), .B(n10792), .Y(n10784) );
  INVXL U25381 ( .A(n10794), .Y(n10806) );
  NAND2XL U25382 ( .A(n10803), .B(n10806), .Y(n10797) );
  INVXL U25383 ( .A(n10805), .Y(n10795) );
  AOI21XL U25384 ( .A0(n10804), .A1(n10806), .B0(n10795), .Y(n10796) );
  NAND2XL U25385 ( .A(n10800), .B(n10799), .Y(n10801) );
  NAND2X1 U25386 ( .A(n10806), .B(n10805), .Y(n10807) );
  OAI21X1 U25387 ( .A0(n10817), .A1(n10813), .B0(n10814), .Y(n10812) );
  NAND2X1 U25388 ( .A(n10810), .B(n10809), .Y(n10811) );
  XNOR2X4 U25389 ( .A(n10812), .B(n10811), .Y(U1_U2_z0[9]) );
  INVXL U25390 ( .A(n10813), .Y(n10815) );
  NAND2X1 U25391 ( .A(n10815), .B(n10814), .Y(n10816) );
  XOR2X2 U25392 ( .A(n10817), .B(n10816), .Y(U1_U2_z0[8]) );
  XNOR2X2 U25393 ( .A(n10824), .B(n10823), .Y(U1_U2_z0[7]) );
  INVXL U25394 ( .A(n10825), .Y(n10827) );
  INVXL U25395 ( .A(n10836), .Y(n10831) );
  INVXL U25396 ( .A(n10832), .Y(n10834) );
  NAND2XL U25397 ( .A(n10837), .B(n10836), .Y(n10838) );
  INVXL U25398 ( .A(n10840), .Y(n10865) );
  OAI21XL U25399 ( .A0(n10865), .A1(n10861), .B0(n10862), .Y(n10845) );
  INVXL U25400 ( .A(n10841), .Y(n10843) );
  NAND2XL U25401 ( .A(n10843), .B(n10842), .Y(n10844) );
  XNOR2XL U25402 ( .A(n10845), .B(n10844), .Y(U1_U2_z0[3]) );
  NAND2XL U25403 ( .A(n10847), .B(n10852), .Y(n10855) );
  OAI21XL U25404 ( .A0(n10850), .A1(n10849), .B0(n10848), .Y(n10851) );
  AOI21XL U25405 ( .A0(n10853), .A1(n10852), .B0(n10851), .Y(n10854) );
  INVXL U25406 ( .A(n10856), .Y(U1_U2_z0[26]) );
  XNOR2X1 U25407 ( .A(n7991), .B(BOPD[26]), .Y(U1_U2_z0[0]) );
  INVXL U25408 ( .A(n10857), .Y(n10859) );
  INVXL U25409 ( .A(n10861), .Y(n10863) );
  NOR2XL U25410 ( .A(n10900), .B(n10890), .Y(n10870) );
  NOR2XL U25411 ( .A(n10906), .B(n10872), .Y(n11021) );
  NAND2XL U25412 ( .A(n11021), .B(n10881), .Y(n10875) );
  NAND2XL U25413 ( .A(n8094), .B(AOPD[48]), .Y(n10901) );
  NAND2XL U25414 ( .A(n8091), .B(AOPD[49]), .Y(n10891) );
  OAI21XL U25415 ( .A0(n10890), .A1(n10901), .B0(n10891), .Y(n10869) );
  AOI21XL U25416 ( .A0(n11027), .A1(n10881), .B0(n10873), .Y(n10874) );
  INVXL U25417 ( .A(n11021), .Y(n10880) );
  INVXL U25418 ( .A(n11027), .Y(n10879) );
  NAND2X1 U25419 ( .A(n10881), .B(n11023), .Y(n10882) );
  INVXL U25420 ( .A(n10896), .Y(n10884) );
  NOR2XL U25421 ( .A(n10884), .B(n10900), .Y(n10887) );
  NAND2XL U25422 ( .A(n10887), .B(n10894), .Y(n10889) );
  INVXL U25423 ( .A(n10895), .Y(n10885) );
  OAI21XL U25424 ( .A0(n10885), .A1(n10900), .B0(n10901), .Y(n10886) );
  AOI21XL U25425 ( .A0(n10897), .A1(n10887), .B0(n10886), .Y(n10888) );
  OAI21X2 U25426 ( .A0(n7197), .A1(n10889), .B0(n10888), .Y(n10893) );
  INVXL U25427 ( .A(n10890), .Y(n10892) );
  NAND2XL U25428 ( .A(n10894), .B(n10896), .Y(n10899) );
  AOI21XL U25429 ( .A0(n10897), .A1(n10896), .B0(n10895), .Y(n10898) );
  XNOR2X2 U25430 ( .A(n10904), .B(n10903), .Y(U0_U2_z0[22]) );
  NAND2X1 U25431 ( .A(n10908), .B(n10907), .Y(n10909) );
  XNOR2X4 U25432 ( .A(n10910), .B(n10909), .Y(U0_U2_z0[20]) );
  NAND2X1 U25433 ( .A(n10917), .B(n10916), .Y(n10918) );
  XNOR2X4 U25434 ( .A(n10919), .B(n10918), .Y(U0_U2_z0[19]) );
  OAI21X2 U25435 ( .A0(n7197), .A1(n10930), .B0(n10931), .Y(n10929) );
  XOR2X1 U25436 ( .A(n11030), .B(n10933), .Y(U0_U2_z0[16]) );
  INVXL U25437 ( .A(n10946), .Y(n10934) );
  NOR2XL U25438 ( .A(n10934), .B(n10949), .Y(n10937) );
  NAND2X1 U25439 ( .A(n10937), .B(n10955), .Y(n10939) );
  INVXL U25440 ( .A(n10945), .Y(n10935) );
  OAI21XL U25441 ( .A0(n10935), .A1(n10949), .B0(n10950), .Y(n10936) );
  AOI21XL U25442 ( .A0(n10957), .A1(n10937), .B0(n10936), .Y(n10938) );
  INVXL U25443 ( .A(n10940), .Y(n10942) );
  NAND2XL U25444 ( .A(n10955), .B(n10946), .Y(n10948) );
  AOI21X1 U25445 ( .A0(n10957), .A1(n10946), .B0(n10945), .Y(n10947) );
  INVXL U25446 ( .A(n10949), .Y(n10951) );
  XNOR2X2 U25447 ( .A(n10953), .B(n10952), .Y(U0_U2_z0[14]) );
  NAND2XL U25448 ( .A(n10955), .B(n10968), .Y(n10959) );
  AOI21X1 U25449 ( .A0(n10957), .A1(n10968), .B0(n10956), .Y(n10958) );
  NAND2XL U25450 ( .A(n10962), .B(n10961), .Y(n10963) );
  XNOR2X2 U25451 ( .A(n10964), .B(n10963), .Y(U0_U2_z0[13]) );
  INVXL U25452 ( .A(n10970), .Y(n10984) );
  INVXL U25453 ( .A(n10983), .Y(n10971) );
  AOI21XL U25454 ( .A0(n10980), .A1(n10984), .B0(n10971), .Y(n10972) );
  NAND2XL U25455 ( .A(n10976), .B(n10975), .Y(n10977) );
  XNOR2X1 U25456 ( .A(n10978), .B(n10977), .Y(U0_U2_z0[11]) );
  XNOR2X2 U25457 ( .A(n10986), .B(n10985), .Y(U0_U2_z0[10]) );
  NAND2X1 U25458 ( .A(n10991), .B(n10990), .Y(n10992) );
  NAND2X1 U25459 ( .A(n10987), .B(n10995), .Y(n10996) );
  INVXL U25460 ( .A(n10998), .Y(n11000) );
  NAND2XL U25461 ( .A(n11000), .B(n10999), .Y(n11001) );
  XOR2X1 U25462 ( .A(n11002), .B(n11001), .Y(U0_U2_z0[6]) );
  INVXL U25463 ( .A(n11003), .Y(n11011) );
  INVXL U25464 ( .A(n11010), .Y(n11004) );
  AOI21X1 U25465 ( .A0(n11013), .A1(n11011), .B0(n11004), .Y(n11009) );
  INVXL U25466 ( .A(n11005), .Y(n11007) );
  NAND2XL U25467 ( .A(n11007), .B(n11006), .Y(n11008) );
  XOR2X1 U25468 ( .A(n11009), .B(n11008), .Y(U0_U2_z0[5]) );
  NAND2XL U25469 ( .A(n11011), .B(n11010), .Y(n11012) );
  INVXL U25470 ( .A(n11014), .Y(n11041) );
  OAI21XL U25471 ( .A0(n11041), .A1(n11037), .B0(n11038), .Y(n11019) );
  XNOR2X1 U25472 ( .A(n11019), .B(n11018), .Y(U0_U2_z0[3]) );
  NAND2XL U25473 ( .A(n11021), .B(n11026), .Y(n11029) );
  OAI21XL U25474 ( .A0(n11024), .A1(n11023), .B0(n11022), .Y(n11025) );
  AOI21XL U25475 ( .A0(n11027), .A1(n11026), .B0(n11025), .Y(n11028) );
  OAI21XL U25476 ( .A0(n7197), .A1(n11029), .B0(n11028), .Y(n11031) );
  INVXL U25477 ( .A(n11031), .Y(U0_U2_z0[26]) );
  XNOR2X1 U25478 ( .A(n8207), .B(AOPD[26]), .Y(U0_U2_z0[0]) );
  INVXL U25479 ( .A(n11032), .Y(n11034) );
  NAND2XL U25480 ( .A(n11208), .B(n11043), .Y(n11045) );
  AOI21XL U25481 ( .A0(n11214), .A1(n11043), .B0(n11042), .Y(n11044) );
  INVXL U25482 ( .A(n11061), .Y(n11049) );
  NOR2XL U25483 ( .A(n11049), .B(n11064), .Y(n11052) );
  NAND2XL U25484 ( .A(n11052), .B(n11070), .Y(n11054) );
  INVXL U25485 ( .A(n11060), .Y(n11050) );
  OAI21XL U25486 ( .A0(n11050), .A1(n11064), .B0(n11065), .Y(n11051) );
  AOI21XL U25487 ( .A0(n11072), .A1(n11052), .B0(n11051), .Y(n11053) );
  NAND2XL U25488 ( .A(n11070), .B(n11061), .Y(n11063) );
  AOI21XL U25489 ( .A0(n11072), .A1(n11061), .B0(n11060), .Y(n11062) );
  NAND2X1 U25490 ( .A(n11066), .B(n11065), .Y(n11067) );
  XNOR2X2 U25491 ( .A(n11068), .B(n11067), .Y(U1_U1_z0[22]) );
  NAND2XL U25492 ( .A(n11070), .B(n11082), .Y(n11074) );
  AOI21XL U25493 ( .A0(n11072), .A1(n11082), .B0(n11071), .Y(n11073) );
  AOI21XL U25494 ( .A0(n11093), .A1(n11097), .B0(n11084), .Y(n11085) );
  INVXL U25495 ( .A(n11087), .Y(n11089) );
  XNOR2X1 U25496 ( .A(n11091), .B(n11090), .Y(U1_U1_z0[19]) );
  INVXL U25497 ( .A(n11120), .Y(n11108) );
  NOR2XL U25498 ( .A(n11108), .B(n11123), .Y(n11111) );
  INVXL U25499 ( .A(n11140), .Y(n11129) );
  NAND2XL U25500 ( .A(n11111), .B(n11129), .Y(n11113) );
  INVXL U25501 ( .A(n11119), .Y(n11109) );
  OAI21XL U25502 ( .A0(n11109), .A1(n11123), .B0(n11124), .Y(n11110) );
  AOI21XL U25503 ( .A0(n11131), .A1(n11111), .B0(n11110), .Y(n11112) );
  OAI21X2 U25504 ( .A0(n11141), .A1(n11113), .B0(n11112), .Y(n11118) );
  INVXL U25505 ( .A(n11114), .Y(n11116) );
  NAND2X1 U25506 ( .A(n11116), .B(n11115), .Y(n11117) );
  XNOR2X4 U25507 ( .A(n11118), .B(n11117), .Y(U1_U1_z0[15]) );
  NAND2XL U25508 ( .A(n11129), .B(n11120), .Y(n11122) );
  NAND2X1 U25509 ( .A(n11125), .B(n11124), .Y(n11126) );
  XNOR2X4 U25510 ( .A(n11127), .B(n11126), .Y(U1_U1_z0[14]) );
  NAND2XL U25511 ( .A(n11129), .B(n11143), .Y(n11133) );
  NAND2X1 U25512 ( .A(n11136), .B(n11135), .Y(n11137) );
  XNOR2X4 U25513 ( .A(n11138), .B(n11137), .Y(U1_U1_z0[13]) );
  XNOR2X2 U25514 ( .A(n11145), .B(n11144), .Y(U1_U1_z0[12]) );
  INVXL U25515 ( .A(n11159), .Y(n11147) );
  INVXL U25516 ( .A(n11155), .Y(n11158) );
  OAI21X1 U25517 ( .A0(n11172), .A1(n11158), .B0(n11157), .Y(n11162) );
  NAND2XL U25518 ( .A(n11160), .B(n11159), .Y(n11161) );
  XNOR2X1 U25519 ( .A(n11162), .B(n11161), .Y(U1_U1_z0[10]) );
  XOR2X2 U25520 ( .A(n11172), .B(n11171), .Y(U1_U1_z0[8]) );
  INVX2 U25521 ( .A(n11173), .Y(n11195) );
  NAND2XL U25522 ( .A(n11178), .B(n11177), .Y(n11179) );
  INVXL U25523 ( .A(n11181), .Y(n11183) );
  NAND2XL U25524 ( .A(n11183), .B(n11182), .Y(n11184) );
  INVXL U25525 ( .A(n11185), .Y(n11193) );
  AOI21XL U25526 ( .A0(n11195), .A1(n11193), .B0(n11186), .Y(n11191) );
  NAND2XL U25527 ( .A(n11189), .B(n11188), .Y(n11190) );
  XOR2X1 U25528 ( .A(n11191), .B(n11190), .Y(U1_U1_z0[5]) );
  XNOR2X2 U25529 ( .A(n11195), .B(n11194), .Y(U1_U1_z0[4]) );
  OAI21XL U25530 ( .A0(n11206), .A1(n11202), .B0(n11203), .Y(n11201) );
  XNOR2X1 U25531 ( .A(n11201), .B(n11200), .Y(U1_U1_z0[3]) );
  INVXL U25532 ( .A(n11202), .Y(n11204) );
  NAND2XL U25533 ( .A(n11204), .B(n11203), .Y(n11205) );
  NOR2XL U25534 ( .A(n11211), .B(n11207), .Y(n11213) );
  NAND2XL U25535 ( .A(n11208), .B(n11213), .Y(n11216) );
  OAI21XL U25536 ( .A0(n11211), .A1(n11210), .B0(n11209), .Y(n11212) );
  INVXL U25537 ( .A(n11217), .Y(U1_U1_z0[26]) );
  INVXL U25538 ( .A(n11218), .Y(n11220) );
  NAND2XL U25539 ( .A(n11220), .B(n11219), .Y(n11221) );
  NOR2XL U25540 ( .A(n11222), .B(n11224), .Y(n11252) );
  NOR2XL U25541 ( .A(n11256), .B(n11246), .Y(n11226) );
  NOR2XL U25542 ( .A(n11262), .B(n11228), .Y(n11380) );
  NAND2XL U25543 ( .A(n11380), .B(n11237), .Y(n11231) );
  NAND2XL U25544 ( .A(n8093), .B(AOPC[48]), .Y(n11257) );
  NAND2XL U25545 ( .A(n8090), .B(AOPC[49]), .Y(n11247) );
  OAI21XL U25546 ( .A0(n11246), .A1(n11257), .B0(n11247), .Y(n11225) );
  AOI21XL U25547 ( .A0(n11386), .A1(n11237), .B0(n11229), .Y(n11230) );
  INVXL U25548 ( .A(n11380), .Y(n11236) );
  INVXL U25549 ( .A(n11386), .Y(n11235) );
  NAND2X1 U25550 ( .A(n11237), .B(n11382), .Y(n11238) );
  INVXL U25551 ( .A(n11252), .Y(n11240) );
  NOR2XL U25552 ( .A(n11240), .B(n11256), .Y(n11243) );
  NAND2XL U25553 ( .A(n11243), .B(n11250), .Y(n11245) );
  INVXL U25554 ( .A(n11251), .Y(n11241) );
  OAI21XL U25555 ( .A0(n11241), .A1(n11256), .B0(n11257), .Y(n11242) );
  INVXL U25556 ( .A(n11246), .Y(n11248) );
  NAND2XL U25557 ( .A(n11250), .B(n11252), .Y(n11255) );
  AOI21XL U25558 ( .A0(n11253), .A1(n11252), .B0(n11251), .Y(n11254) );
  NAND2X1 U25559 ( .A(n11264), .B(n11263), .Y(n11265) );
  XNOR2X4 U25560 ( .A(n11266), .B(n11265), .Y(U0_U1_z0[20]) );
  NAND2X1 U25561 ( .A(n11273), .B(n11272), .Y(n11274) );
  XNOR2X4 U25562 ( .A(n11275), .B(n11274), .Y(U0_U1_z0[19]) );
  NAND2X1 U25563 ( .A(n11281), .B(n11280), .Y(n11282) );
  NAND2X1 U25564 ( .A(n11290), .B(n11289), .Y(n11291) );
  INVXL U25565 ( .A(n11302), .Y(n11292) );
  NOR2XL U25566 ( .A(n11292), .B(n11305), .Y(n11293) );
  INVXL U25567 ( .A(n11322), .Y(n11311) );
  NAND2XL U25568 ( .A(n11293), .B(n11311), .Y(n11296) );
  INVXL U25569 ( .A(n11301), .Y(n11294) );
  OAI21XL U25570 ( .A0(n11294), .A1(n11305), .B0(n11306), .Y(n11295) );
  NAND2XL U25571 ( .A(n11311), .B(n11302), .Y(n11304) );
  INVX1 U25572 ( .A(n11321), .Y(n11313) );
  AOI21X1 U25573 ( .A0(n11313), .A1(n11302), .B0(n11301), .Y(n11303) );
  NAND2X1 U25574 ( .A(n11307), .B(n11306), .Y(n11308) );
  NAND2XL U25575 ( .A(n11311), .B(n11324), .Y(n11315) );
  AOI21X1 U25576 ( .A0(n11313), .A1(n11324), .B0(n11312), .Y(n11314) );
  NAND2XL U25577 ( .A(n11318), .B(n11317), .Y(n11319) );
  XNOR2X1 U25578 ( .A(n11320), .B(n11319), .Y(U0_U1_z0[13]) );
  OAI21XL U25579 ( .A0(n11348), .A1(n11322), .B0(n11321), .Y(n11326) );
  NAND2XL U25580 ( .A(n11324), .B(n11323), .Y(n11325) );
  XNOR2X1 U25581 ( .A(n11326), .B(n11325), .Y(U0_U1_z0[12]) );
  NAND2XL U25582 ( .A(n11336), .B(n11341), .Y(n11330) );
  AOI21XL U25583 ( .A0(n11337), .A1(n11341), .B0(n11328), .Y(n11329) );
  OAI21XL U25584 ( .A0(n11348), .A1(n11330), .B0(n11329), .Y(n11335) );
  NAND2XL U25585 ( .A(n11333), .B(n11332), .Y(n11334) );
  XNOR2X1 U25586 ( .A(n11335), .B(n11334), .Y(U0_U1_z0[11]) );
  INVXL U25587 ( .A(n11336), .Y(n11339) );
  OAI21X1 U25588 ( .A0(n11348), .A1(n11339), .B0(n11338), .Y(n11343) );
  XNOR2X2 U25589 ( .A(n11343), .B(n11342), .Y(U0_U1_z0[10]) );
  INVXL U25590 ( .A(n11352), .Y(n11354) );
  XNOR2X2 U25591 ( .A(n11356), .B(n11355), .Y(U0_U1_z0[7]) );
  NAND2XL U25592 ( .A(n11359), .B(n11358), .Y(n11360) );
  XOR2X1 U25593 ( .A(n11361), .B(n11360), .Y(U0_U1_z0[6]) );
  INVXL U25594 ( .A(n11362), .Y(n11370) );
  INVXL U25595 ( .A(n11369), .Y(n11363) );
  AOI21X1 U25596 ( .A0(n11372), .A1(n11370), .B0(n11363), .Y(n11368) );
  INVXL U25597 ( .A(n11364), .Y(n11366) );
  NAND2XL U25598 ( .A(n11366), .B(n11365), .Y(n11367) );
  XOR2X1 U25599 ( .A(n11368), .B(n11367), .Y(U0_U1_z0[5]) );
  NAND2XL U25600 ( .A(n11370), .B(n11369), .Y(n11371) );
  OAI21XL U25601 ( .A0(n11395), .A1(n11391), .B0(n11392), .Y(n11378) );
  INVXL U25602 ( .A(n11374), .Y(n11376) );
  NAND2XL U25603 ( .A(n11376), .B(n11375), .Y(n11377) );
  XNOR2X1 U25604 ( .A(n11378), .B(n11377), .Y(U0_U1_z0[3]) );
  NAND2XL U25605 ( .A(n11380), .B(n11385), .Y(n11388) );
  OAI21XL U25606 ( .A0(n11383), .A1(n11382), .B0(n11381), .Y(n11384) );
  AOI21XL U25607 ( .A0(n11386), .A1(n11385), .B0(n11384), .Y(n11387) );
  OAI21XL U25608 ( .A0(n11389), .A1(n11388), .B0(n11387), .Y(n11390) );
  INVXL U25609 ( .A(n11390), .Y(U0_U1_z0[26]) );
  INVXL U25610 ( .A(n11391), .Y(n11393) );
  INVXL U25611 ( .A(n11396), .Y(n11398) );
  NAND2XL U25612 ( .A(n11398), .B(n11397), .Y(n11400) );
  OAI21XL U25613 ( .A0(n28684), .A1(n11428), .B0(n11412), .Y(U2_B_r[23]) );
  OAI21XL U25614 ( .A0(n28708), .A1(n11430), .B0(n11420), .Y(U2_B_r[20]) );
  OAI21XL U25615 ( .A0(n28749), .A1(n11430), .B0(n11429), .Y(U2_B_r[25]) );
  AOI21X4 U25616 ( .A0(n11436), .A1(n11435), .B0(n11434), .Y(n11502) );
  NAND2X1 U25617 ( .A(n11439), .B(U2_B_r[15]), .Y(n11535) );
  NAND2X1 U25618 ( .A(n11441), .B(U2_B_r[16]), .Y(n11530) );
  NAND2XL U25619 ( .A(n5824), .B(U2_B_r[17]), .Y(n11522) );
  INVXL U25620 ( .A(n11522), .Y(n11442) );
  OAI21X4 U25621 ( .A0(n11502), .A1(n11449), .B0(n11448), .Y(n11607) );
  NOR2X1 U25622 ( .A(n11452), .B(n7118), .Y(n11490) );
  INVXL U25623 ( .A(U2_B_i[20]), .Y(n11450) );
  NOR2XL U25624 ( .A(n11450), .B(U2_B_r[20]), .Y(n11495) );
  NOR2X1 U25625 ( .A(n11497), .B(n11495), .Y(n11489) );
  NOR2XL U25626 ( .A(n11471), .B(n11462), .Y(n11458) );
  NAND2X1 U25627 ( .A(n11450), .B(U2_B_r[20]), .Y(n11604) );
  OAI21X2 U25628 ( .A0(n11497), .A1(n11604), .B0(n11498), .Y(n11488) );
  NAND2XL U25629 ( .A(n11453), .B(U2_B_r[23]), .Y(n11484) );
  AOI21X2 U25630 ( .A0(n11607), .A1(n11458), .B0(n11457), .Y(n11461) );
  OR2X2 U25631 ( .A(U2_B_i[25]), .B(n11459), .Y(n11466) );
  NAND2XL U25632 ( .A(U2_B_i[25]), .B(n11459), .Y(n11463) );
  XOR2X4 U25633 ( .A(n11461), .B(n11460), .Y(U2_U0_z0[25]) );
  NAND2XL U25634 ( .A(n11466), .B(n11476), .Y(n11468) );
  NOR2XL U25635 ( .A(n11471), .B(n11468), .Y(n11470) );
  INVXL U25636 ( .A(n11475), .Y(n11465) );
  INVXL U25637 ( .A(n11463), .Y(n11464) );
  AOI21XL U25638 ( .A0(n11466), .A1(n11465), .B0(n11464), .Y(n11467) );
  OAI21XL U25639 ( .A0(n11472), .A1(n11468), .B0(n11467), .Y(n11469) );
  AOI21X2 U25640 ( .A0(n11607), .A1(n11470), .B0(n11469), .Y(U2_U0_z0[26]) );
  INVXL U25641 ( .A(n11471), .Y(n11474) );
  INVXL U25642 ( .A(n11472), .Y(n11473) );
  AOI21X2 U25643 ( .A0(n11607), .A1(n11474), .B0(n11473), .Y(n11478) );
  INVXL U25644 ( .A(n11489), .Y(n11479) );
  NOR2XL U25645 ( .A(n11479), .B(n11490), .Y(n11482) );
  INVXL U25646 ( .A(n11488), .Y(n11480) );
  OAI21XL U25647 ( .A0(n11480), .A1(n11490), .B0(n11491), .Y(n11481) );
  AOI21X2 U25648 ( .A0(n11607), .A1(n11482), .B0(n11481), .Y(n11487) );
  INVXL U25649 ( .A(n11483), .Y(n11485) );
  XOR2X4 U25650 ( .A(n11487), .B(n11486), .Y(U2_U0_z0[23]) );
  INVXL U25651 ( .A(n11490), .Y(n11492) );
  INVXL U25652 ( .A(n11495), .Y(n11605) );
  INVXL U25653 ( .A(n11604), .Y(n11496) );
  INVXL U25654 ( .A(n11497), .Y(n11499) );
  INVXL U25655 ( .A(n11513), .Y(n11503) );
  NOR2XL U25656 ( .A(n11503), .B(n11514), .Y(n11506) );
  INVXL U25657 ( .A(n11512), .Y(n11504) );
  INVXL U25658 ( .A(n11507), .Y(n11509) );
  XOR2X4 U25659 ( .A(n11511), .B(n11510), .Y(U2_U0_z0[19]) );
  INVXL U25660 ( .A(n11514), .Y(n11516) );
  NOR2XL U25661 ( .A(n11526), .B(n11519), .Y(n11521) );
  OAI21XL U25662 ( .A0(n11527), .A1(n11519), .B0(n11530), .Y(n11520) );
  NAND2X1 U25663 ( .A(n11523), .B(n11522), .Y(n11524) );
  INVX1 U25664 ( .A(n11526), .Y(n11529) );
  INVX1 U25665 ( .A(n11527), .Y(n11528) );
  NAND2X1 U25666 ( .A(n11536), .B(n11535), .Y(n11537) );
  NAND2X1 U25667 ( .A(n11540), .B(n11539), .Y(n11541) );
  NAND2X1 U25668 ( .A(n11545), .B(n11544), .Y(n11546) );
  XNOR2X4 U25669 ( .A(n11547), .B(n11546), .Y(U2_U0_z0[12]) );
  NAND2X1 U25670 ( .A(n11549), .B(n8147), .Y(n11550) );
  INVXL U25671 ( .A(n11567), .Y(n11556) );
  NOR2XL U25672 ( .A(n11556), .B(n11568), .Y(n11561) );
  INVXL U25673 ( .A(n11558), .Y(n11559) );
  OAI21XL U25674 ( .A0(n11559), .A1(n11568), .B0(n11569), .Y(n11560) );
  INVXL U25675 ( .A(n11562), .Y(n11564) );
  NAND2XL U25676 ( .A(n11564), .B(n11563), .Y(n11565) );
  XOR2X2 U25677 ( .A(n11566), .B(n11565), .Y(U2_U0_z0[9]) );
  AOI21X1 U25678 ( .A0(n11582), .A1(n11567), .B0(n11558), .Y(n11572) );
  INVXL U25679 ( .A(n11568), .Y(n11570) );
  INVX1 U25680 ( .A(n11573), .Y(n11580) );
  NAND2X1 U25681 ( .A(n11576), .B(n11575), .Y(n11577) );
  XNOR2X4 U25682 ( .A(n11582), .B(n11581), .Y(U2_U0_z0[6]) );
  INVXL U25683 ( .A(n11586), .Y(n11588) );
  XNOR2X4 U25684 ( .A(n11590), .B(n11589), .Y(U2_U0_z0[5]) );
  NAND2X1 U25685 ( .A(n11597), .B(n11596), .Y(n11598) );
  XOR2X2 U25686 ( .A(n11602), .B(n11601), .Y(U2_U0_z0[1]) );
  XNOR2X1 U25687 ( .A(n11603), .B(U2_B_r[0]), .Y(U2_U0_z0[0]) );
  NAND2XL U25688 ( .A(n11605), .B(n11604), .Y(n11606) );
  NAND2XL U25689 ( .A(n11633), .B(n11648), .Y(n28643) );
  OAI21XL U25690 ( .A0(n28679), .A1(n28705), .B0(n11965), .Y(n11611) );
  OAI21XL U25691 ( .A0(n11611), .A1(n11610), .B0(n11609), .Y(n11612) );
  INVX1 U25692 ( .A(n11998), .Y(n11999) );
  OAI222X4 U25693 ( .A0(n11625), .A1(n28673), .B0(n28679), .B1(n11633), .C0(
        n11873), .C1(n11618), .Y(n11874) );
  NAND2XL U25694 ( .A(cnt[6]), .B(n11633), .Y(n11624) );
  OAI21XL U25695 ( .A0(n28709), .A1(n11633), .B0(n11624), .Y(n28665) );
  OAI21XL U25696 ( .A0(n28705), .A1(n11633), .B0(n11618), .Y(n28659) );
  OAI21XL U25697 ( .A0(n11999), .A1(n28666), .B0(n11621), .Y(n11619) );
  OAI21XL U25698 ( .A0(n11913), .A1(n28705), .B0(n11619), .Y(n11620) );
  OAI21XL U25699 ( .A0(n11998), .A1(n28666), .B0(n11621), .Y(n11622) );
  OAI21XL U25700 ( .A0(n11913), .A1(n28705), .B0(n11622), .Y(n11623) );
  OAI222X4 U25701 ( .A0(n11625), .A1(n28680), .B0(n28674), .B1(n11633), .C0(
        n11873), .C1(n11624), .Y(n28642) );
  AOI21XL U25702 ( .A0(n15023), .A1(n11984), .B0(n28642), .Y(n11626) );
  AOI2BB2XL U25703 ( .B0(cs[0]), .B1(n28698), .A0N(in_valid), .A1N(cs[0]), .Y(
        n11631) );
  NAND2X2 U25704 ( .A(cs[1]), .B(n28912), .Y(n11954) );
  INVX1 U25705 ( .A(n11954), .Y(n11628) );
  OAI21XL U25706 ( .A0(n5927), .A1(n29107), .B0(n11951), .Y(n11946) );
  OAI21XL U25707 ( .A0(n11638), .A1(n11629), .B0(n11946), .Y(n11630) );
  AOI21XL U25708 ( .A0(n11636), .A1(n11631), .B0(n11630), .Y(n5681) );
  NAND2XL U25709 ( .A(n11633), .B(n11632), .Y(n11907) );
  AOI21XL U25710 ( .A0(n11908), .A1(n15024), .B0(n28639), .Y(n11634) );
  AOI22X1 U25711 ( .A0(n28699), .A1(cs[2]), .B0(n28986), .B1(n27236), .Y(
        n11974) );
  INVX1 U25712 ( .A(n11974), .Y(n11968) );
  AOI211X1 U25713 ( .A0(n11948), .A1(n11638), .B0(cs[2]), .C0(n11637), .Y(
        n28631) );
  NOR2X1 U25714 ( .A(n28631), .B(n11968), .Y(n28630) );
  AOI21XL U25715 ( .A0(cnt[5]), .A1(n11968), .B0(n11639), .Y(n5674) );
  AOI211XL U25716 ( .A0(n28704), .A1(n11641), .B0(n11973), .C0(n11966), .Y(
        n11642) );
  AOI21XL U25717 ( .A0(cnt[6]), .A1(n11968), .B0(n11642), .Y(n5673) );
  NOR2X1 U25718 ( .A(n28698), .B(S_EN), .Y(n11989) );
  AOI22X2 U25719 ( .A0(cnt[8]), .A1(n15024), .B0(n11984), .B1(n28706), .Y(
        n11992) );
  NOR2X1 U25720 ( .A(n28986), .B(n28698), .Y(n11991) );
  NOR2X1 U25721 ( .A(cnt[8]), .B(n11949), .Y(n11652) );
  AOI21XL U25722 ( .A0(cnt[5]), .A1(n11652), .B0(n11972), .Y(n11651) );
  NOR2X4 U25723 ( .A(n28704), .B(n14979), .Y(T1_rom_addr[0]) );
  NOR2X4 U25724 ( .A(n28703), .B(n14979), .Y(T1_rom_addr[1]) );
  NAND2X1 U25725 ( .A(n15027), .B(out_sel), .Y(n11653) );
  OR2X2 U25726 ( .A(n14993), .B(n11653), .Y(n11679) );
  OR2X2 U25727 ( .A(n14994), .B(n11654), .Y(n11709) );
  OR2X2 U25728 ( .A(n14994), .B(n11653), .Y(n11677) );
  OR2X2 U25729 ( .A(n14993), .B(n11654), .Y(n11684) );
  OR2X2 U25730 ( .A(n14998), .B(n11653), .Y(n11719) );
  OR2X2 U25731 ( .A(n14998), .B(n11654), .Y(n11678) );
  OR2X2 U25732 ( .A(n11655), .B(n11654), .Y(n11710) );
  OAI21XL U25733 ( .A0(n28706), .A1(n11949), .B0(n11948), .Y(n5693) );
  AOI21XL U25734 ( .A0(n11998), .A1(n15023), .B0(n11874), .Y(n11875) );
  AOI22XL U25735 ( .A0(n11878), .A1(cnt[3]), .B0(cnt[1]), .B1(n29107), .Y(
        n11879) );
  AOI21XL U25736 ( .A0(n11998), .A1(n11885), .B0(n28637), .Y(n11880) );
  OAI22X2 U25737 ( .A0(n15025), .A1(cnt[7]), .B0(n11881), .B1(n15027), .Y(
        n11882) );
  OAI2BB2X2 U25738 ( .B0(n15025), .B1(cnt[7]), .A0N(n11883), .A1N(n15025), .Y(
        n11884) );
  AOI21XL U25739 ( .A0(n11885), .A1(n11984), .B0(n28636), .Y(n11886) );
  OAI2BB2X2 U25740 ( .B0(n11887), .B1(n15027), .A0N(n15027), .A1N(n28704), .Y(
        n11888) );
  AOI21XL U25741 ( .A0(n11908), .A1(n11984), .B0(n28639), .Y(n11889) );
  OAI2BB2X2 U25742 ( .B0(n15025), .B1(cnt[4]), .A0N(n11889), .A1N(n15025), .Y(
        n11890) );
  AOI21XL U25743 ( .A0(n28252), .A1(Q0_addr[1]), .B0(n27073), .Y(n11893) );
  NAND3X1 U25744 ( .A(A_sel_reg[0]), .B(C_sel_reg[1]), .C(n5922), .Y(n11930)
         );
  NAND3X2 U25745 ( .A(n27298), .B(n14981), .C(n11930), .Y(n27389) );
  NOR2X2 U25746 ( .A(C_sel_reg[1]), .B(n15003), .Y(n27390) );
  OAI211X4 U25747 ( .A0(n28753), .A1(n5916), .B0(n11893), .C0(n11892), .Y(
        A1_addr[1]) );
  AOI21XL U25748 ( .A0(n28252), .A1(Q0_addr[0]), .B0(n27081), .Y(n11895) );
  OAI211X4 U25749 ( .A0(n28752), .A1(n5916), .B0(n11895), .C0(n11894), .Y(
        A1_addr[0]) );
  AOI32X4 U25750 ( .A0(n15025), .A1(n11899), .A2(n11898), .B0(cnt[0]), .B1(
        n15027), .Y(n11900) );
  AOI21XL U25751 ( .A0(n28252), .A1(Q0_addr[5]), .B0(n15028), .Y(n11902) );
  OAI211X4 U25752 ( .A0(n28757), .A1(n5825), .B0(n11902), .C0(n11901), .Y(
        A1_addr[5]) );
  AOI21XL U25753 ( .A0(n28252), .A1(Q0_addr[3]), .B0(n14988), .Y(n11904) );
  OAI211X4 U25754 ( .A0(n28756), .A1(n5825), .B0(n11904), .C0(n11903), .Y(
        A1_addr[3]) );
  AOI21XL U25755 ( .A0(n28252), .A1(Q0_addr[4]), .B0(n27078), .Y(n11906) );
  OAI211X4 U25756 ( .A0(n28754), .A1(n5916), .B0(n11906), .C0(n11905), .Y(
        A1_addr[4]) );
  AOI21XL U25757 ( .A0(n28252), .A1(Q0_addr[2]), .B0(n27084), .Y(n11915) );
  OAI211X4 U25758 ( .A0(n28755), .A1(n5916), .B0(n11915), .C0(n11914), .Y(
        A1_addr[2]) );
  AOI21XL U25759 ( .A0(n28252), .A1(Q0_addr[7]), .B0(n15038), .Y(n11917) );
  OAI211X4 U25760 ( .A0(n28920), .A1(n5825), .B0(n11917), .C0(n11916), .Y(
        A1_addr[7]) );
  AOI21XL U25761 ( .A0(n28252), .A1(Q0_addr[6]), .B0(n15031), .Y(n11919) );
  OAI211X4 U25762 ( .A0(n28919), .A1(n5825), .B0(n11919), .C0(n11918), .Y(
        A1_addr[6]) );
  AOI21XL U25763 ( .A0(n5921), .A1(Q0_addr[7]), .B0(n15038), .Y(n11922) );
  NAND2X1 U25764 ( .A(n28322), .B(C_sel_reg[1]), .Y(n27386) );
  NAND3BX2 U25765 ( .AN(n11929), .B(n14980), .C(n11931), .Y(n27281) );
  OAI211X4 U25766 ( .A0(n28920), .A1(n27379), .B0(n11922), .C0(n11921), .Y(
        A2_addr[7]) );
  AOI21XL U25767 ( .A0(n5921), .A1(Q0_addr[5]), .B0(n15028), .Y(n11924) );
  OAI211X4 U25768 ( .A0(n28757), .A1(n27379), .B0(n11924), .C0(n11923), .Y(
        A2_addr[5]) );
  AOI21XL U25769 ( .A0(n5921), .A1(Q0_addr[6]), .B0(n15031), .Y(n11926) );
  OAI211X4 U25770 ( .A0(n28919), .A1(n27379), .B0(n11926), .C0(n11925), .Y(
        A2_addr[6]) );
  AOI21XL U25771 ( .A0(n5921), .A1(Q0_addr[3]), .B0(n14988), .Y(n11928) );
  OAI211X4 U25772 ( .A0(n28756), .A1(n27379), .B0(n11928), .C0(n11927), .Y(
        A2_addr[3]) );
  AOI21XL U25773 ( .A0(n27631), .A1(Q0_addr[7]), .B0(n15038), .Y(n11933) );
  NAND3X2 U25774 ( .A(n15003), .B(n11931), .C(n11930), .Y(n27497) );
  OAI211X4 U25775 ( .A0(n28920), .A1(n27772), .B0(n11933), .C0(n11932), .Y(
        A0_addr[7]) );
  AOI21XL U25776 ( .A0(n27631), .A1(Q0_addr[6]), .B0(n15031), .Y(n11935) );
  OAI211X4 U25777 ( .A0(n28919), .A1(n27772), .B0(n11935), .C0(n11934), .Y(
        A0_addr[6]) );
  AOI21XL U25778 ( .A0(n27631), .A1(Q0_addr[5]), .B0(n15028), .Y(n11937) );
  OAI211X4 U25779 ( .A0(n28757), .A1(n27772), .B0(n11937), .C0(n11936), .Y(
        A0_addr[5]) );
  AOI21XL U25780 ( .A0(n27631), .A1(Q0_addr[4]), .B0(n27078), .Y(n11939) );
  OAI211X4 U25781 ( .A0(n28754), .A1(n27772), .B0(n11939), .C0(n11938), .Y(
        A0_addr[4]) );
  AOI21XL U25782 ( .A0(n5798), .A1(Q0_addr[3]), .B0(n14988), .Y(n11942) );
  OAI211X4 U25783 ( .A0(n28756), .A1(n27772), .B0(n11942), .C0(n11941), .Y(
        A0_addr[3]) );
  AOI21XL U25784 ( .A0(n5827), .A1(Q0_addr[1]), .B0(n27073), .Y(n11944) );
  OAI211X4 U25785 ( .A0(n28753), .A1(n27772), .B0(n11944), .C0(n11943), .Y(
        A0_addr[1]) );
  NAND2XL U25786 ( .A(n11945), .B(DATA0[5]), .Y(n5743) );
  NAND2XL U25787 ( .A(n11945), .B(DATA0[27]), .Y(n5721) );
  NAND2XL U25788 ( .A(n11945), .B(DATA0[41]), .Y(n5707) );
  NAND2XL U25789 ( .A(n11945), .B(DATA0[3]), .Y(n5745) );
  NAND2XL U25790 ( .A(n11945), .B(DATA0[39]), .Y(n5709) );
  NAND2XL U25791 ( .A(n11945), .B(DATA0[37]), .Y(n5711) );
  NAND2XL U25792 ( .A(n11945), .B(DATA0[49]), .Y(n5699) );
  NAND2XL U25793 ( .A(n11945), .B(DATA0[31]), .Y(n5717) );
  NAND2XL U25794 ( .A(n11945), .B(DATA0[29]), .Y(n5719) );
  NAND2XL U25795 ( .A(n11945), .B(DATA0[45]), .Y(n5703) );
  NAND2XL U25796 ( .A(n11945), .B(DATA0[19]), .Y(n5729) );
  NAND2XL U25797 ( .A(n11945), .B(DATA0[9]), .Y(n5739) );
  NAND2XL U25798 ( .A(n11945), .B(DATA0[23]), .Y(n5725) );
  NAND2XL U25799 ( .A(n11945), .B(DATA0[21]), .Y(n5727) );
  NAND2XL U25800 ( .A(n11945), .B(DATA0[11]), .Y(n5737) );
  NAND2XL U25801 ( .A(n11945), .B(DATA0[13]), .Y(n5735) );
  NAND2XL U25802 ( .A(n11945), .B(DATA0[1]), .Y(n5747) );
  NAND2XL U25803 ( .A(n11945), .B(DATA0[47]), .Y(n5701) );
  AOI211XL U25804 ( .A0(n27236), .A1(n28698), .B0(n11948), .C0(n11947), .Y(
        n5683) );
  OAI21XL U25805 ( .A0(n11949), .A1(n29012), .B0(n15027), .Y(n5695) );
  OAI21XL U25806 ( .A0(n15025), .A1(n28699), .B0(n5695), .Y(n11950) );
  CLKINVX3 U25807 ( .A(n5808), .Y(n11953) );
  AOI22XL U25808 ( .A0(n5834), .A1(Q3_addr[28]), .B0(Q3_addr[20]), .B1(n5808), 
        .Y(n5480) );
  AOI22XL U25809 ( .A0(n15027), .A1(cnt[10]), .B0(out_sel), .B1(n15025), .Y(
        n5156) );
  AOI22XL U25810 ( .A0(n5834), .A1(Q1_addr[34]), .B0(Q1_addr[26]), .B1(n5808), 
        .Y(n5519) );
  AOI22XL U25811 ( .A0(n5834), .A1(Q1_addr[10]), .B0(Q1_addr[2]), .B1(n5808), 
        .Y(n5516) );
  AOI22XL U25812 ( .A0(n11953), .A1(Q1_addr[33]), .B0(Q1_addr[25]), .B1(n5808), 
        .Y(n5524) );
  AOI21XL U25813 ( .A0(n28629), .A1(n28705), .B0(n28631), .Y(n11955) );
  AOI21XL U25814 ( .A0(n28703), .A1(n11959), .B0(n11975), .Y(n11960) );
  AOI21XL U25815 ( .A0(n11963), .A1(n28679), .B0(n11962), .Y(n11964) );
  AOI21XL U25816 ( .A0(n28680), .A1(n11967), .B0(n11966), .Y(n11970) );
  OAI21XL U25817 ( .A0(n28635), .A1(n11976), .B0(n29107), .Y(n11977) );
  AOI21XL U25818 ( .A0(n7305), .A1(ram_sel_reg[1]), .B0(n11982), .Y(n11983) );
  OAI21XL U25819 ( .A0(ram_sel_reg[0]), .A1(n11633), .B0(n11985), .Y(n11988)
         );
  AOI21XL U25820 ( .A0(n7305), .A1(ram_sel_reg[1]), .B0(n11988), .Y(n11990) );
  AOI22XL U25821 ( .A0(n12000), .A1(A_sel_reg[0]), .B0(A_sel_reg[1]), .B1(
        n5829), .Y(n5417) );
  AOI22XL U25822 ( .A0(n12000), .A1(C_sel_reg[8]), .B0(n15024), .B1(n5829), 
        .Y(n5416) );
  XOR2X1 U25823 ( .A(n12002), .B(n12001), .Y(n12003) );
  NOR2XL U25824 ( .A(U0_U2_y2[1]), .B(U0_U2_y0[1]), .Y(n12006) );
  INVXL U25825 ( .A(n12006), .Y(n12009) );
  AND2XL U25826 ( .A(U0_U2_y2[0]), .B(U0_U2_y0[0]), .Y(n12008) );
  NOR2XL U25827 ( .A(U0_U2_y2[2]), .B(U0_U2_y0[2]), .Y(n12010) );
  INVXL U25828 ( .A(n12010), .Y(n12012) );
  NAND2XL U25829 ( .A(n12012), .B(n12014), .Y(n12016) );
  OAI21XL U25830 ( .A0(n12017), .A1(n12016), .B0(n12015), .Y(n12035) );
  OAI21XL U25831 ( .A0(n12032), .A1(n12031), .B0(n12030), .Y(n12033) );
  INVXL U25832 ( .A(U0_U2_y2[13]), .Y(n12050) );
  NOR2XL U25833 ( .A(n12050), .B(U0_U2_y0[13]), .Y(n12036) );
  INVXL U25834 ( .A(n12036), .Y(n12052) );
  OR2X2 U25835 ( .A(U0_U2_y2[12]), .B(U0_U2_y0[12]), .Y(n12037) );
  OR2X2 U25836 ( .A(U0_U2_y2[9]), .B(U0_U2_y0[9]), .Y(n12043) );
  OR2X2 U25837 ( .A(U0_U2_y2[10]), .B(U0_U2_y0[10]), .Y(n12039) );
  OR2X2 U25838 ( .A(U0_U2_y2[11]), .B(U0_U2_y0[11]), .Y(n12046) );
  NAND2XL U25839 ( .A(n12055), .B(n12104), .Y(n12057) );
  OAI21XL U25840 ( .A0(n12049), .A1(n12048), .B0(n12047), .Y(n12103) );
  AOI21XL U25841 ( .A0(n12052), .A1(n12051), .B0(n7961), .Y(n12107) );
  NAND2XL U25842 ( .A(n12053), .B(U0_U2_y2[13]), .Y(n12112) );
  OAI21XL U25843 ( .A0(n12107), .A1(n12111), .B0(n12112), .Y(n12054) );
  AOI21XL U25844 ( .A0(n12055), .A1(n12103), .B0(n12054), .Y(n12056) );
  OAI21X2 U25845 ( .A0(n12102), .A1(n12057), .B0(n12056), .Y(n12139) );
  CMPR22X1 U25846 ( .A(U0_U2_y2[14]), .B(U0_U2_y0[14]), .CO(n12059), .S(n12053) );
  CMPR22X1 U25847 ( .A(U0_U2_y2[17]), .B(U0_U2_y0[17]), .CO(n12065), .S(n12062) );
  NAND2XL U25848 ( .A(n12059), .B(n12058), .Y(n12120) );
  NAND2XL U25849 ( .A(n12060), .B(n12061), .Y(n12124) );
  OAI21XL U25850 ( .A0(n12123), .A1(n12120), .B0(n12124), .Y(n12089) );
  NOR2X1 U25851 ( .A(n12069), .B(n12068), .Y(n12078) );
  INVXL U25852 ( .A(n12081), .Y(n12072) );
  XNOR2X2 U25853 ( .A(n12074), .B(n12073), .Y(n13107) );
  XOR2X1 U25854 ( .A(n12077), .B(n12076), .Y(n13106) );
  NOR2XL U25855 ( .A(n25764), .B(n25762), .Y(n25757) );
  ADDHX2 U25856 ( .A(U0_U2_y2[20]), .B(U0_U2_y0[20]), .CO(n12084), .S(n12070)
         );
  NAND2XL U25857 ( .A(n12085), .B(n12148), .Y(n12086) );
  XOR2X1 U25858 ( .A(n12150), .B(n12086), .Y(n13108) );
  NAND2XL U25859 ( .A(n25757), .B(n12087), .Y(n12132) );
  INVXL U25860 ( .A(n12088), .Y(n12091) );
  INVXL U25861 ( .A(n12089), .Y(n12090) );
  INVXL U25862 ( .A(n12094), .Y(n12096) );
  NAND2XL U25863 ( .A(n12096), .B(n12095), .Y(n12097) );
  XNOR2X1 U25864 ( .A(n12101), .B(n12100), .Y(n13102) );
  NOR2XL U25865 ( .A(n24587), .B(n13102), .Y(n25777) );
  NOR2XL U25866 ( .A(n25427), .B(n25777), .Y(n12129) );
  AOI21XL U25867 ( .A0(n12105), .A1(n12104), .B0(n12103), .Y(n12106) );
  INVXL U25868 ( .A(n12111), .Y(n12113) );
  XOR2X1 U25869 ( .A(n12122), .B(n12117), .Y(n13099) );
  NAND2XL U25870 ( .A(n24588), .B(n13099), .Y(n25787) );
  INVXL U25871 ( .A(n25787), .Y(n12119) );
  AOI21XL U25872 ( .A0(n25788), .A1(n12118), .B0(n12119), .Y(n25784) );
  OAI21XL U25873 ( .A0(n12122), .A1(n12121), .B0(n12120), .Y(n12127) );
  INVXL U25874 ( .A(n12123), .Y(n12125) );
  NOR2XL U25875 ( .A(n24595), .B(n13101), .Y(n25437) );
  NAND2XL U25876 ( .A(n24595), .B(n13101), .Y(n25438) );
  OAI21XL U25877 ( .A0(n25784), .A1(n25437), .B0(n25438), .Y(n25775) );
  NAND2XL U25878 ( .A(n24587), .B(n13102), .Y(n25776) );
  NAND2XL U25879 ( .A(n24586), .B(n13103), .Y(n25428) );
  OAI21XL U25880 ( .A0(n25427), .A1(n25776), .B0(n25428), .Y(n12128) );
  AOI21XL U25881 ( .A0(n12129), .A1(n25775), .B0(n12128), .Y(n25755) );
  NAND2XL U25882 ( .A(n24583), .B(n13106), .Y(n25770) );
  NAND2XL U25883 ( .A(n24582), .B(n13107), .Y(n25765) );
  OAI21XL U25884 ( .A0(n25764), .A1(n25770), .B0(n25765), .Y(n25756) );
  NAND2XL U25885 ( .A(n24584), .B(n13108), .Y(n25758) );
  INVXL U25886 ( .A(n25758), .Y(n12130) );
  CMPR22X1 U25887 ( .A(U0_U2_y2[21]), .B(U0_U2_y0[21]), .CO(n12136), .S(n12083) );
  NAND2X1 U25888 ( .A(n12136), .B(n12135), .Y(n12152) );
  OAI21X1 U25889 ( .A0(n12151), .A1(n12148), .B0(n12152), .Y(n12137) );
  CMPR22X1 U25890 ( .A(U0_U2_y2[22]), .B(U0_U2_y0[22]), .CO(n12141), .S(n12135) );
  NOR2XL U25891 ( .A(n24616), .B(n14530), .Y(n25739) );
  OAI21XL U25892 ( .A0(n12150), .A1(n12149), .B0(n12148), .Y(n12155) );
  INVXL U25893 ( .A(n12151), .Y(n12153) );
  NAND2XL U25894 ( .A(n12153), .B(n12152), .Y(n12154) );
  NOR2XL U25895 ( .A(n24617), .B(n13113), .Y(n25738) );
  INVXL U25896 ( .A(n25738), .Y(n25400) );
  NAND2XL U25897 ( .A(n12170), .B(n25400), .Y(n25725) );
  CMPR22X1 U25898 ( .A(U0_U2_y2[25]), .B(U0_U2_y0[25]), .CO(n12162), .S(n12160) );
  INVXL U25899 ( .A(n12176), .Y(n12164) );
  NOR2XL U25900 ( .A(n24620), .B(n14533), .Y(n12167) );
  INVXL U25901 ( .A(n12167), .Y(n25733) );
  NAND2XL U25902 ( .A(n24617), .B(n13113), .Y(n25737) );
  INVXL U25903 ( .A(n25737), .Y(n12169) );
  NAND2XL U25904 ( .A(n24616), .B(n14530), .Y(n25747) );
  NAND2XL U25905 ( .A(n24620), .B(n14533), .Y(n25732) );
  INVXL U25906 ( .A(n25732), .Y(n25726) );
  NAND2XL U25907 ( .A(n24619), .B(n14532), .Y(n25727) );
  INVXL U25908 ( .A(n25727), .Y(n12171) );
  ADDHX2 U25909 ( .A(U0_U2_y2[28]), .B(U0_U2_y0[28]), .CO(n12186), .S(n12183)
         );
  NOR2X4 U25910 ( .A(n12188), .B(n12187), .Y(n12210) );
  NAND2X1 U25911 ( .A(n12188), .B(n12187), .Y(n12208) );
  OR2X2 U25912 ( .A(n24644), .B(n13125), .Y(n25705) );
  NOR2XL U25913 ( .A(n24645), .B(n14547), .Y(n25703) );
  NAND2X1 U25914 ( .A(n12197), .B(n12196), .Y(n12198) );
  NAND2XL U25915 ( .A(n12201), .B(n12200), .Y(n12202) );
  XOR2X1 U25916 ( .A(n12203), .B(n12202), .Y(n14548) );
  NOR2X1 U25917 ( .A(n12234), .B(n25699), .Y(n25679) );
  ADDHX2 U25918 ( .A(U0_U2_y0[30]), .B(U0_U2_y2[30]), .CO(n12214), .S(n12187)
         );
  ADDHX2 U25919 ( .A(U0_U2_y2[31]), .B(U0_U2_y0[31]), .CO(n12216), .S(n12213)
         );
  NAND2X2 U25920 ( .A(n12214), .B(n12213), .Y(n12230) );
  CMPR22X1 U25921 ( .A(U0_U2_y2[33]), .B(U0_U2_y0[33]), .CO(n12220), .S(n12217) );
  INVXL U25922 ( .A(n12245), .Y(n12221) );
  NAND2X1 U25923 ( .A(n25328), .B(n25332), .Y(n12240) );
  INVXL U25924 ( .A(n12225), .Y(n12227) );
  NAND2XL U25925 ( .A(n24647), .B(n14548), .Y(n25720) );
  NAND2XL U25926 ( .A(n24646), .B(n13123), .Y(n25715) );
  NAND2XL U25927 ( .A(n24645), .B(n14547), .Y(n25709) );
  INVXL U25928 ( .A(n25709), .Y(n12232) );
  NAND2XL U25929 ( .A(n24644), .B(n13125), .Y(n25704) );
  INVXL U25930 ( .A(n25704), .Y(n12231) );
  INVXL U25931 ( .A(n25691), .Y(n12236) );
  INVXL U25932 ( .A(n25338), .Y(n12235) );
  INVXL U25933 ( .A(n25683), .Y(n12238) );
  NAND2XL U25934 ( .A(n24640), .B(n13131), .Y(n25327) );
  INVXL U25935 ( .A(n25327), .Y(n12237) );
  AOI21X1 U25936 ( .A0(n25328), .A1(n12238), .B0(n12237), .Y(n12239) );
  OAI21XL U25937 ( .A0(n12247), .A1(n12252), .B0(n12256), .Y(n12251) );
  CMPR22X1 U25938 ( .A(U0_U2_y2[34]), .B(U0_U2_y0[34]), .CO(n12249), .S(n12219) );
  XNOR2X2 U25939 ( .A(n12251), .B(n12250), .Y(n13166) );
  NOR2XL U25940 ( .A(n24674), .B(n13166), .Y(n25670) );
  INVXL U25941 ( .A(n25670), .Y(n25315) );
  CMPR22X1 U25942 ( .A(U0_U2_y2[35]), .B(U0_U2_y0[35]), .CO(n12261), .S(n12248) );
  NAND2XL U25943 ( .A(n25315), .B(n25311), .Y(n25665) );
  NOR2X1 U25944 ( .A(n12266), .B(n12265), .Y(n12272) );
  XOR2X2 U25945 ( .A(n12273), .B(n12268), .Y(n14570) );
  NOR2XL U25946 ( .A(n24676), .B(n14570), .Y(n25302) );
  NAND2XL U25947 ( .A(n24674), .B(n13166), .Y(n25669) );
  INVXL U25948 ( .A(n25669), .Y(n12270) );
  NAND2XL U25949 ( .A(n24675), .B(n13167), .Y(n25310) );
  INVXL U25950 ( .A(n25310), .Y(n12269) );
  NAND2XL U25951 ( .A(n24676), .B(n14570), .Y(n25303) );
  CMPR22X1 U25952 ( .A(U0_U2_y2[37]), .B(U0_U2_y0[37]), .CO(n12276), .S(n12265) );
  CMPR22X1 U25953 ( .A(U0_U2_y2[38]), .B(U0_U2_y0[38]), .CO(n12282), .S(n12275) );
  NAND2XL U25954 ( .A(n24692), .B(n14579), .Y(n25650) );
  NOR2XL U25955 ( .A(n12295), .B(U1_A_r_d0[5]), .Y(n19923) );
  NOR2XL U25956 ( .A(n19917), .B(n19923), .Y(n20279) );
  NAND2XL U25957 ( .A(n20279), .B(n12286), .Y(n12299) );
  NOR2XL U25958 ( .A(n12292), .B(U1_A_r_d0[4]), .Y(n19930) );
  NOR2XL U25959 ( .A(n12291), .B(U1_A_r_d0[3]), .Y(n20294) );
  NOR2XL U25960 ( .A(n19930), .B(n20294), .Y(n12294) );
  NAND2XL U25961 ( .A(n12288), .B(U1_A_r_d0[1]), .Y(n19946) );
  INVXL U25962 ( .A(n19946), .Y(n12289) );
  AOI21XL U25963 ( .A0(n20304), .A1(n12287), .B0(n12289), .Y(n20301) );
  NOR2XL U25964 ( .A(n12290), .B(U1_A_r_d0[2]), .Y(n19940) );
  OAI21XL U25965 ( .A0(n20301), .A1(n19940), .B0(n19941), .Y(n20292) );
  NAND2XL U25966 ( .A(n12291), .B(U1_A_r_d0[3]), .Y(n20293) );
  NAND2XL U25967 ( .A(n12292), .B(U1_A_r_d0[4]), .Y(n19931) );
  OAI21XL U25968 ( .A0(n19930), .A1(n20293), .B0(n19931), .Y(n12293) );
  AOI21XL U25969 ( .A0(n12294), .A1(n20292), .B0(n12293), .Y(n20277) );
  NAND2XL U25970 ( .A(n12295), .B(U1_A_r_d0[5]), .Y(n20283) );
  OAI21XL U25971 ( .A0(n19917), .A1(n20283), .B0(n19918), .Y(n20278) );
  NAND2XL U25972 ( .A(n12296), .B(U1_A_r_d0[7]), .Y(n19909) );
  INVXL U25973 ( .A(n19909), .Y(n12297) );
  AOI21XL U25974 ( .A0(n20278), .A1(n12286), .B0(n12297), .Y(n12298) );
  OAI21XL U25975 ( .A0(n12299), .A1(n20277), .B0(n12298), .Y(n20253) );
  NOR2XL U25976 ( .A(n19732), .B(U1_A_r_d0[9]), .Y(n19898) );
  NOR2XL U25977 ( .A(n19892), .B(n19898), .Y(n12304) );
  NOR2XL U25978 ( .A(n12301), .B(U1_A_r_d0[8]), .Y(n20264) );
  INVXL U25979 ( .A(n20264), .Y(n19902) );
  NAND2X1 U25980 ( .A(n12304), .B(n19902), .Y(n20255) );
  NOR2X1 U25981 ( .A(n20255), .B(n12307), .Y(n12309) );
  NAND2XL U25982 ( .A(n12301), .B(U1_A_r_d0[8]), .Y(n20263) );
  INVXL U25983 ( .A(n20263), .Y(n12303) );
  NAND2XL U25984 ( .A(n19732), .B(U1_A_r_d0[9]), .Y(n20265) );
  OAI21XL U25985 ( .A0(n19892), .A1(n20265), .B0(n19893), .Y(n12302) );
  AOI21X1 U25986 ( .A0(n12304), .A1(n12303), .B0(n12302), .Y(n20254) );
  NAND2XL U25987 ( .A(n19736), .B(U1_A_r_d0[11]), .Y(n19882) );
  INVXL U25988 ( .A(n19882), .Y(n20256) );
  NAND2XL U25989 ( .A(n19734), .B(U1_A_r_d0[12]), .Y(n19877) );
  INVXL U25990 ( .A(n19877), .Y(n12305) );
  AOI21XL U25991 ( .A0(n19878), .A1(n20256), .B0(n12305), .Y(n12306) );
  AOI21X1 U25992 ( .A0(n20253), .A1(n12309), .B0(n12308), .Y(n20208) );
  OR2X2 U25993 ( .A(n19751), .B(U1_A_r_d0[16]), .Y(n19854) );
  NOR2XL U25994 ( .A(n12313), .B(U1_A_r_d0[15]), .Y(n20237) );
  INVXL U25995 ( .A(n20237), .Y(n19858) );
  NAND2XL U25996 ( .A(n19854), .B(n19858), .Y(n12317) );
  OR2X2 U25997 ( .A(n12311), .B(U1_A_r_d0[13]), .Y(n20246) );
  NAND2XL U25998 ( .A(n12310), .B(n20246), .Y(n20232) );
  NOR2XL U25999 ( .A(n12317), .B(n20232), .Y(n20210) );
  INVXL U26000 ( .A(n20216), .Y(n19833) );
  NOR2XL U26001 ( .A(n19756), .B(U1_A_r_d0[17]), .Y(n20224) );
  INVXL U26002 ( .A(n20224), .Y(n19843) );
  NAND2XL U26003 ( .A(n12311), .B(U1_A_r_d0[13]), .Y(n19868) );
  INVXL U26004 ( .A(n19868), .Y(n20245) );
  NAND2XL U26005 ( .A(n19754), .B(U1_A_r_d0[14]), .Y(n19864) );
  INVXL U26006 ( .A(n19864), .Y(n12312) );
  NAND2XL U26007 ( .A(n12313), .B(U1_A_r_d0[15]), .Y(n20236) );
  INVXL U26008 ( .A(n20236), .Y(n12315) );
  NAND2X1 U26009 ( .A(n19751), .B(U1_A_r_d0[16]), .Y(n19853) );
  INVXL U26010 ( .A(n19853), .Y(n12314) );
  AOI21XL U26011 ( .A0(n19854), .A1(n12315), .B0(n12314), .Y(n12316) );
  OAI21X1 U26012 ( .A0(n12317), .A1(n20233), .B0(n12316), .Y(n20209) );
  INVXL U26013 ( .A(n20223), .Y(n12319) );
  INVXL U26014 ( .A(n19838), .Y(n12318) );
  AOI21X1 U26015 ( .A0(n19839), .A1(n12319), .B0(n12318), .Y(n20212) );
  INVXL U26016 ( .A(n20215), .Y(n12321) );
  INVXL U26017 ( .A(n19828), .Y(n12320) );
  OAI21XL U26018 ( .A0(n12323), .A1(n20212), .B0(n12322), .Y(n12324) );
  NOR2XL U26019 ( .A(n12327), .B(U1_A_r_d0[21]), .Y(n20201) );
  INVXL U26020 ( .A(n20201), .Y(n19818) );
  NOR2XL U26021 ( .A(n19773), .B(U1_A_r_d0[22]), .Y(n12326) );
  INVXL U26022 ( .A(n12326), .Y(n19814) );
  NAND2XL U26023 ( .A(n19818), .B(n19814), .Y(n20196) );
  NOR2XL U26024 ( .A(n19774), .B(U1_A_r_d0[23]), .Y(n19805) );
  NOR2XL U26025 ( .A(n20196), .B(n19805), .Y(n12331) );
  NAND2XL U26026 ( .A(n12327), .B(U1_A_r_d0[21]), .Y(n20200) );
  INVXL U26027 ( .A(n20200), .Y(n12329) );
  NAND2XL U26028 ( .A(n19773), .B(U1_A_r_d0[22]), .Y(n19813) );
  INVXL U26029 ( .A(n19813), .Y(n12328) );
  AOI21XL U26030 ( .A0(n12329), .A1(n19814), .B0(n12328), .Y(n20195) );
  NAND2XL U26031 ( .A(n19774), .B(U1_A_r_d0[23]), .Y(n19806) );
  NAND2XL U26032 ( .A(n12334), .B(U1_A_r_d0[25]), .Y(n19791) );
  INVX1 U26033 ( .A(n12335), .Y(n12336) );
  MXI2X1 U26034 ( .A(U1_pipe8[27]), .B(n12336), .S0(n5812), .Y(n4809) );
  MXI2X1 U26035 ( .A(U1_pipe14[27]), .B(n12340), .S0(n24784), .Y(n4778) );
  OAI21XL U26036 ( .A0(n12350), .A1(n12349), .B0(n12348), .Y(n12354) );
  NOR2XL U26037 ( .A(n14526), .B(n24582), .Y(n25413) );
  NOR2XL U26038 ( .A(n14525), .B(n24583), .Y(n25411) );
  NOR2XL U26039 ( .A(n25413), .B(n25411), .Y(n25406) );
  NAND2XL U26040 ( .A(n25406), .B(n12362), .Y(n12373) );
  NOR2XL U26041 ( .A(n14522), .B(n24586), .Y(n12368) );
  NOR2XL U26042 ( .A(n14521), .B(n24587), .Y(n25426) );
  NOR2XL U26043 ( .A(n12368), .B(n25426), .Y(n12370) );
  OR2X2 U26044 ( .A(n14515), .B(n24588), .Y(n25444) );
  NAND2XL U26045 ( .A(n14515), .B(n24588), .Y(n25443) );
  INVXL U26046 ( .A(n25443), .Y(n12363) );
  AOI21XL U26047 ( .A0(n12364), .A1(n25444), .B0(n12363), .Y(n25440) );
  INVX1 U26048 ( .A(n13101), .Y(n14518) );
  NOR2XL U26049 ( .A(n14518), .B(n24595), .Y(n12366) );
  NAND2XL U26050 ( .A(n14518), .B(n24595), .Y(n12365) );
  OAI21XL U26051 ( .A0(n25440), .A1(n12366), .B0(n12365), .Y(n25424) );
  NAND2XL U26052 ( .A(n14521), .B(n24587), .Y(n25425) );
  NAND2XL U26053 ( .A(n14522), .B(n24586), .Y(n12367) );
  OAI21XL U26054 ( .A0(n12368), .A1(n25425), .B0(n12367), .Y(n12369) );
  AOI21XL U26055 ( .A0(n12370), .A1(n25424), .B0(n12369), .Y(n25404) );
  NAND2XL U26056 ( .A(n14525), .B(n24583), .Y(n25419) );
  NAND2XL U26057 ( .A(n14526), .B(n24582), .Y(n25414) );
  OAI21XL U26058 ( .A0(n25413), .A1(n25419), .B0(n25414), .Y(n25405) );
  NAND2XL U26059 ( .A(n14527), .B(n24584), .Y(n25407) );
  INVXL U26060 ( .A(n25407), .Y(n12371) );
  AOI21XL U26061 ( .A0(n25405), .A1(n12362), .B0(n12371), .Y(n12372) );
  OAI21XL U26062 ( .A0(n12373), .A1(n25404), .B0(n12372), .Y(n25372) );
  NOR2XL U26063 ( .A(n14535), .B(n24616), .Y(n25387) );
  INVX1 U26064 ( .A(n13113), .Y(n14534) );
  NOR2XL U26065 ( .A(n14534), .B(n24617), .Y(n25386) );
  INVXL U26066 ( .A(n25386), .Y(n12374) );
  NAND2XL U26067 ( .A(n12377), .B(n12374), .Y(n25374) );
  NAND2XL U26068 ( .A(n14534), .B(n24617), .Y(n25385) );
  INVXL U26069 ( .A(n25385), .Y(n12376) );
  NAND2XL U26070 ( .A(n14535), .B(n24616), .Y(n25395) );
  OAI21XL U26071 ( .A0(n25389), .A1(n25395), .B0(n25390), .Y(n12375) );
  AOI21X1 U26072 ( .A0(n12377), .A1(n12376), .B0(n12375), .Y(n25373) );
  NAND2XL U26073 ( .A(n12378), .B(n24620), .Y(n25381) );
  INVXL U26074 ( .A(n25381), .Y(n25375) );
  NAND2XL U26075 ( .A(n12379), .B(n24619), .Y(n25376) );
  INVXL U26076 ( .A(n25376), .Y(n12380) );
  NOR2XL U26077 ( .A(n5852), .B(n24641), .Y(n12386) );
  INVXL U26078 ( .A(n12386), .Y(n25326) );
  NAND2X1 U26079 ( .A(n7963), .B(n25326), .Y(n12396) );
  NOR2XL U26080 ( .A(n14560), .B(n24643), .Y(n12387) );
  INVXL U26081 ( .A(n12387), .Y(n25337) );
  NOR2X2 U26082 ( .A(n12396), .B(n25324), .Y(n12397) );
  NAND2XL U26083 ( .A(n12388), .B(n24647), .Y(n25368) );
  INVXL U26084 ( .A(n25368), .Y(n25362) );
  INVXL U26085 ( .A(n25363), .Y(n12389) );
  NAND2XL U26086 ( .A(n5864), .B(n24645), .Y(n25357) );
  INVXL U26087 ( .A(n25357), .Y(n12391) );
  NAND2XL U26088 ( .A(n14555), .B(n24644), .Y(n25352) );
  INVXL U26089 ( .A(n25352), .Y(n12390) );
  AND2X2 U26090 ( .A(n5852), .B(n24641), .Y(n25325) );
  AOI21XL U26091 ( .A0(n7963), .A1(n25325), .B0(n7964), .Y(n12395) );
  CLKINVX3 U26092 ( .A(n13166), .Y(n14571) );
  NOR2XL U26093 ( .A(n14571), .B(n24674), .Y(n25309) );
  NOR2XL U26094 ( .A(n14572), .B(n24675), .Y(n12399) );
  NOR2XL U26095 ( .A(n25309), .B(n12399), .Y(n25298) );
  NAND2XL U26096 ( .A(n25298), .B(n8083), .Y(n25291) );
  NAND2XL U26097 ( .A(n14571), .B(n24674), .Y(n25308) );
  NAND2XL U26098 ( .A(n14572), .B(n24675), .Y(n12398) );
  OAI21XL U26099 ( .A0(n25308), .A1(n12399), .B0(n12398), .Y(n25299) );
  AOI21X1 U26100 ( .A0(n25299), .A1(n8083), .B0(n8082), .Y(n25290) );
  NAND2XL U26101 ( .A(n14577), .B(n24677), .Y(n12400) );
  NOR2X1 U26102 ( .A(n12404), .B(n24692), .Y(n12406) );
  NAND2XL U26103 ( .A(n12404), .B(n24692), .Y(n12405) );
  MXI2X1 U26104 ( .A(U0_pipe13[26]), .B(n12407), .S0(n5812), .Y(n4666) );
  OR2XL U26105 ( .A(U0_U1_y2[1]), .B(U0_U1_y0[1]), .Y(n12410) );
  AND2XL U26106 ( .A(U0_U1_y2[0]), .B(U0_U1_y0[0]), .Y(n12409) );
  AOI21XL U26107 ( .A0(n12410), .A1(n12409), .B0(n12408), .Y(n12417) );
  NAND2XL U26108 ( .A(n12411), .B(n12414), .Y(n12416) );
  AND2XL U26109 ( .A(U0_U1_y2[2]), .B(U0_U1_y0[2]), .Y(n12413) );
  AOI21XL U26110 ( .A0(n12414), .A1(n12413), .B0(n12412), .Y(n12415) );
  OAI21XL U26111 ( .A0(n12417), .A1(n12416), .B0(n12415), .Y(n12432) );
  OR2X2 U26112 ( .A(U0_U1_y2[5]), .B(U0_U1_y0[5]), .Y(n12423) );
  OR2X2 U26113 ( .A(U0_U1_y2[6]), .B(U0_U1_y0[6]), .Y(n12419) );
  OR2X2 U26114 ( .A(U0_U1_y2[7]), .B(U0_U1_y0[7]), .Y(n12426) );
  AOI21XL U26115 ( .A0(n12423), .A1(n12422), .B0(n12421), .Y(n12429) );
  AOI21XL U26116 ( .A0(n12426), .A1(n12425), .B0(n12424), .Y(n12427) );
  OAI21XL U26117 ( .A0(n12429), .A1(n12428), .B0(n12427), .Y(n12430) );
  AOI21XL U26118 ( .A0(n12432), .A1(n12431), .B0(n12430), .Y(n12492) );
  OR2X2 U26119 ( .A(U0_U1_y2[12]), .B(U0_U1_y0[12]), .Y(n12433) );
  OR2X2 U26120 ( .A(U0_U1_y2[9]), .B(U0_U1_y0[9]), .Y(n12439) );
  OR2X2 U26121 ( .A(U0_U1_y2[10]), .B(U0_U1_y0[10]), .Y(n12435) );
  OR2X2 U26122 ( .A(U0_U1_y2[11]), .B(U0_U1_y0[11]), .Y(n12442) );
  OAI21XL U26123 ( .A0(n12445), .A1(n12444), .B0(n12443), .Y(n12493) );
  NAND2XL U26124 ( .A(n12449), .B(U0_U1_y2[13]), .Y(n12503) );
  OAI21XL U26125 ( .A0(n12498), .A1(n12502), .B0(n12503), .Y(n12450) );
  CMPR22X1 U26126 ( .A(U0_U1_y2[14]), .B(U0_U1_y0[14]), .CO(n12455), .S(n12449) );
  NOR2XL U26127 ( .A(n12488), .B(n12482), .Y(n12511) );
  NOR2XL U26128 ( .A(n12516), .B(n12518), .Y(n12463) );
  NAND2X1 U26129 ( .A(n12511), .B(n12463), .Y(n12531) );
  OAI21XL U26130 ( .A0(n12482), .A1(n12489), .B0(n12483), .Y(n12512) );
  OAI21XL U26131 ( .A0(n12518), .A1(n12523), .B0(n12519), .Y(n12462) );
  AOI21X1 U26132 ( .A0(n12463), .A1(n12512), .B0(n12462), .Y(n12539) );
  OAI21X1 U26133 ( .A0(n12515), .A1(n12531), .B0(n12539), .Y(n12476) );
  CMPR22X1 U26134 ( .A(U0_U1_y2[18]), .B(U0_U1_y0[18]), .CO(n12465), .S(n12460) );
  INVXL U26135 ( .A(n12475), .Y(n12468) );
  NAND2XL U26136 ( .A(n12468), .B(n12473), .Y(n12469) );
  NOR2XL U26137 ( .A(n24608), .B(n22885), .Y(n22696) );
  NOR2XL U26138 ( .A(n24606), .B(n22886), .Y(n22694) );
  NOR2XL U26139 ( .A(n22696), .B(n22694), .Y(n22689) );
  OAI21XL U26140 ( .A0(n12475), .A1(n12474), .B0(n12473), .Y(n12535) );
  AOI21XL U26141 ( .A0(n12476), .A1(n12530), .B0(n12535), .Y(n12554) );
  INVXL U26142 ( .A(n12553), .Y(n12479) );
  NAND2XL U26143 ( .A(n12479), .B(n12552), .Y(n12480) );
  XOR2X1 U26144 ( .A(n12554), .B(n12480), .Y(n22887) );
  NOR2XL U26145 ( .A(n24610), .B(n22887), .Y(n12481) );
  OAI21XL U26146 ( .A0(n12515), .A1(n12488), .B0(n12489), .Y(n12486) );
  INVXL U26147 ( .A(n12482), .Y(n12484) );
  NOR2XL U26148 ( .A(n24596), .B(n22897), .Y(n12487) );
  INVXL U26149 ( .A(n12487), .Y(n22720) );
  NAND2XL U26150 ( .A(n22720), .B(n22724), .Y(n12510) );
  INVXL U26151 ( .A(n12497), .Y(n12500) );
  NAND2XL U26152 ( .A(n24596), .B(n22897), .Y(n22719) );
  INVXL U26153 ( .A(n22719), .Y(n12507) );
  AOI21XL U26154 ( .A0(n22720), .A1(n12508), .B0(n12507), .Y(n12509) );
  INVXL U26155 ( .A(n12511), .Y(n12514) );
  INVXL U26156 ( .A(n12512), .Y(n12513) );
  OAI21XL U26157 ( .A0(n12515), .A1(n12514), .B0(n12513), .Y(n12526) );
  INVXL U26158 ( .A(n12516), .Y(n12524) );
  INVXL U26159 ( .A(n12523), .Y(n12517) );
  AOI21XL U26160 ( .A0(n12526), .A1(n12524), .B0(n12517), .Y(n12522) );
  INVXL U26161 ( .A(n12518), .Y(n12520) );
  NAND2XL U26162 ( .A(n12520), .B(n12519), .Y(n12521) );
  XOR2X1 U26163 ( .A(n12522), .B(n12521), .Y(n22889) );
  NOR2XL U26164 ( .A(n24602), .B(n22889), .Y(n22708) );
  NAND2XL U26165 ( .A(n12524), .B(n12523), .Y(n12525) );
  NOR2XL U26166 ( .A(n24600), .B(n22890), .Y(n22713) );
  NOR2XL U26167 ( .A(n22708), .B(n22713), .Y(n12528) );
  OAI21XL U26168 ( .A0(n22708), .A1(n22714), .B0(n22709), .Y(n12527) );
  NAND2XL U26169 ( .A(n24606), .B(n22886), .Y(n22702) );
  NAND2XL U26170 ( .A(n24608), .B(n22885), .Y(n22697) );
  OAI21XL U26171 ( .A0(n22696), .A1(n22702), .B0(n22697), .Y(n22688) );
  NAND2XL U26172 ( .A(n24610), .B(n22887), .Y(n22690) );
  NAND2X1 U26173 ( .A(n12544), .B(n12543), .Y(n12561) );
  INVXL U26174 ( .A(n12562), .Y(n12547) );
  NAND2XL U26175 ( .A(n12549), .B(n12561), .Y(n12550) );
  XNOR2X1 U26176 ( .A(n12551), .B(n12550), .Y(n22914) );
  NOR2XL U26177 ( .A(n22914), .B(n24623), .Y(n22670) );
  OAI21XL U26178 ( .A0(n12554), .A1(n12553), .B0(n12552), .Y(n12558) );
  NOR2XL U26179 ( .A(n24621), .B(n22915), .Y(n22669) );
  INVXL U26180 ( .A(n22669), .Y(n22684) );
  NAND2XL U26181 ( .A(n12575), .B(n22684), .Y(n22659) );
  NOR2XL U26182 ( .A(n12559), .B(n12562), .Y(n12582) );
  INVXL U26183 ( .A(n12582), .Y(n12563) );
  CMPR22X1 U26184 ( .A(U0_U1_y2[24]), .B(U0_U1_y0[24]), .CO(n12565), .S(n12545) );
  NOR2X1 U26185 ( .A(n12565), .B(n12564), .Y(n12581) );
  INVXL U26186 ( .A(n12585), .Y(n12568) );
  NOR2X1 U26187 ( .A(n22659), .B(n12578), .Y(n12580) );
  INVXL U26188 ( .A(n22683), .Y(n12574) );
  NAND2XL U26189 ( .A(n22914), .B(n24623), .Y(n22678) );
  OAI21XL U26190 ( .A0(n22672), .A1(n22678), .B0(n22673), .Y(n12573) );
  NAND2XL U26191 ( .A(n22918), .B(n24631), .Y(n22665) );
  INVXL U26192 ( .A(n22665), .Y(n22660) );
  NAND2XL U26193 ( .A(n22917), .B(n24633), .Y(n22661) );
  INVXL U26194 ( .A(n22661), .Y(n12576) );
  OAI21XL U26195 ( .A0(n12585), .A1(n12584), .B0(n12583), .Y(n12586) );
  NAND2XL U26196 ( .A(n12594), .B(n12622), .Y(n12595) );
  XOR2X1 U26197 ( .A(n12596), .B(n12595), .Y(n22934) );
  NOR2XL U26198 ( .A(n22934), .B(n24652), .Y(n22636) );
  INVXL U26199 ( .A(n22636), .Y(n22643) );
  INVXL U26200 ( .A(n12623), .Y(n12599) );
  NAND2XL U26201 ( .A(n12609), .B(n12608), .Y(n12610) );
  XOR2X1 U26202 ( .A(n12611), .B(n12610), .Y(n22936) );
  NAND2XL U26203 ( .A(n22649), .B(n12612), .Y(n22632) );
  NOR2XL U26204 ( .A(n12617), .B(n22632), .Y(n14113) );
  NAND2XL U26205 ( .A(n22936), .B(n24649), .Y(n22653) );
  INVXL U26206 ( .A(n22653), .Y(n22647) );
  INVXL U26207 ( .A(n22648), .Y(n12613) );
  NAND2XL U26208 ( .A(n22934), .B(n24652), .Y(n22642) );
  INVXL U26209 ( .A(n22642), .Y(n12615) );
  INVXL U26210 ( .A(n22637), .Y(n12614) );
  AOI21XL U26211 ( .A0(n22638), .A1(n12615), .B0(n12614), .Y(n12616) );
  OAI21XL U26212 ( .A0(n12617), .A1(n22633), .B0(n12616), .Y(n14122) );
  ADDHX2 U26213 ( .A(U0_U1_y2[31]), .B(U0_U1_y0[31]), .CO(n12631), .S(n12628)
         );
  INVXL U26214 ( .A(n12640), .Y(n12632) );
  NAND2X1 U26215 ( .A(n5886), .B(n12639), .Y(n12633) );
  NOR2XL U26216 ( .A(n24661), .B(n22933), .Y(n22622) );
  INVXL U26217 ( .A(n22622), .Y(n22629) );
  NAND2X1 U26218 ( .A(n6904), .B(n22629), .Y(n14112) );
  INVXL U26219 ( .A(n22628), .Y(n12635) );
  NAND2XL U26220 ( .A(n24662), .B(n22932), .Y(n22624) );
  INVXL U26221 ( .A(n22624), .Y(n12634) );
  INVXL U26222 ( .A(n14119), .Y(n12636) );
  OAI21X1 U26223 ( .A0(n22619), .A1(n14111), .B0(n22616), .Y(n12648) );
  INVXL U26224 ( .A(n13138), .Y(n12646) );
  NAND2XL U26225 ( .A(n24666), .B(n22930), .Y(n14114) );
  MXI2X1 U26226 ( .A(U0_pipe15[20]), .B(n12649), .S0(n5812), .Y(n4616) );
  NOR2XL U26227 ( .A(U1_U1_y2[1]), .B(U1_U1_y0[1]), .Y(n12650) );
  INVXL U26228 ( .A(n12650), .Y(n12653) );
  AND2XL U26229 ( .A(U1_U1_y2[0]), .B(U1_U1_y0[0]), .Y(n12652) );
  AOI21XL U26230 ( .A0(n12653), .A1(n12652), .B0(n12651), .Y(n12661) );
  NOR2XL U26231 ( .A(U1_U1_y2[3]), .B(U1_U1_y0[3]), .Y(n12655) );
  INVXL U26232 ( .A(n12655), .Y(n12658) );
  NAND2XL U26233 ( .A(n12656), .B(n12658), .Y(n12660) );
  AOI21XL U26234 ( .A0(n12658), .A1(n7020), .B0(n12657), .Y(n12659) );
  OAI21XL U26235 ( .A0(n12661), .A1(n12660), .B0(n12659), .Y(n12678) );
  NOR2XL U26236 ( .A(U1_U1_y2[5]), .B(U1_U1_y0[5]), .Y(n12663) );
  INVXL U26237 ( .A(n12663), .Y(n12670) );
  NAND2XL U26238 ( .A(n12664), .B(n12670), .Y(n12668) );
  NOR2XL U26239 ( .A(U1_U1_y2[7]), .B(U1_U1_y0[7]), .Y(n12666) );
  INVXL U26240 ( .A(n12666), .Y(n12672) );
  NAND2XL U26241 ( .A(n12667), .B(n12672), .Y(n12674) );
  NOR2XL U26242 ( .A(n12668), .B(n12674), .Y(n12677) );
  AOI21XL U26243 ( .A0(n12670), .A1(n7021), .B0(n12669), .Y(n12675) );
  AOI21XL U26244 ( .A0(n12672), .A1(n7017), .B0(n12671), .Y(n12673) );
  OAI21XL U26245 ( .A0(n12675), .A1(n12674), .B0(n12673), .Y(n12676) );
  OR2X2 U26246 ( .A(n12689), .B(U1_U1_y0[13]), .Y(n12691) );
  NAND2XL U26247 ( .A(n12691), .B(n12679), .Y(n12831) );
  NAND2XL U26248 ( .A(n7979), .B(n12682), .Y(n12687) );
  NOR2XL U26249 ( .A(n12683), .B(n12687), .Y(n12828) );
  AOI21XL U26250 ( .A0(n12681), .A1(n7022), .B0(n12684), .Y(n12688) );
  AOI21XL U26251 ( .A0(n12682), .A1(n7013), .B0(n12685), .Y(n12686) );
  OAI21XL U26252 ( .A0(n12688), .A1(n12687), .B0(n12686), .Y(n12827) );
  AOI21X1 U26253 ( .A0(n12691), .A1(n12690), .B0(n6998), .Y(n12832) );
  NAND2XL U26254 ( .A(n12692), .B(U1_U1_y2[13]), .Y(n12837) );
  OAI21XL U26255 ( .A0(n12832), .A1(n12836), .B0(n12837), .Y(n12693) );
  CMPR22X1 U26256 ( .A(U1_U1_y2[14]), .B(U1_U1_y0[14]), .CO(n12695), .S(n12692) );
  CMPR22X1 U26257 ( .A(U1_U1_y2[17]), .B(U1_U1_y0[17]), .CO(n12701), .S(n12698) );
  CMPR22X1 U26258 ( .A(U1_U1_y2[18]), .B(U1_U1_y0[18]), .CO(n12703), .S(n12700) );
  NOR2X1 U26259 ( .A(n12703), .B(n12702), .Y(n12777) );
  INVXL U26260 ( .A(n14922), .Y(n12885) );
  OR2XL U26261 ( .A(U1_U2_y1[1]), .B(U1_U2_y0[1]), .Y(n12708) );
  AOI21XL U26262 ( .A0(n12708), .A1(n12707), .B0(n8142), .Y(n12717) );
  NOR2XL U26263 ( .A(U1_U2_y1[2]), .B(U1_U2_y0[2]), .Y(n12709) );
  INVXL U26264 ( .A(n12709), .Y(n12711) );
  NOR2XL U26265 ( .A(U1_U2_y1[3]), .B(U1_U2_y0[3]), .Y(n12710) );
  INVXL U26266 ( .A(n12710), .Y(n12714) );
  NAND2XL U26267 ( .A(n12711), .B(n12714), .Y(n12716) );
  AOI21XL U26268 ( .A0(n12714), .A1(n12713), .B0(n12712), .Y(n12715) );
  OAI21XL U26269 ( .A0(n12717), .A1(n12716), .B0(n12715), .Y(n12732) );
  OR2X2 U26270 ( .A(U1_U2_y1[7]), .B(U1_U2_y0[7]), .Y(n12726) );
  NAND2XL U26271 ( .A(n12719), .B(n12726), .Y(n12728) );
  AOI21XL U26272 ( .A0(n12723), .A1(n12722), .B0(n12721), .Y(n12729) );
  OAI21XL U26273 ( .A0(n12729), .A1(n12728), .B0(n12727), .Y(n12730) );
  AOI21XL U26274 ( .A0(n12732), .A1(n12731), .B0(n12730), .Y(n12841) );
  INVXL U26275 ( .A(U1_U2_y1[13]), .Y(n12746) );
  OR2X2 U26276 ( .A(n12746), .B(U1_U2_y0[13]), .Y(n12749) );
  OR2X2 U26277 ( .A(U1_U2_y1[12]), .B(U1_U2_y0[12]), .Y(n12733) );
  NAND2XL U26278 ( .A(n12749), .B(n12733), .Y(n12846) );
  NOR2XL U26279 ( .A(n12846), .B(n12851), .Y(n12752) );
  OR2X2 U26280 ( .A(U1_U2_y1[9]), .B(U1_U2_y0[9]), .Y(n12739) );
  OR2X2 U26281 ( .A(U1_U2_y1[10]), .B(U1_U2_y0[10]), .Y(n12735) );
  OR2X2 U26282 ( .A(U1_U2_y1[11]), .B(U1_U2_y0[11]), .Y(n12742) );
  NAND2XL U26283 ( .A(n12735), .B(n12742), .Y(n12744) );
  NOR2XL U26284 ( .A(n12736), .B(n12744), .Y(n12843) );
  NAND2XL U26285 ( .A(n12752), .B(n12843), .Y(n12754) );
  AOI21XL U26286 ( .A0(n12739), .A1(n12738), .B0(n12737), .Y(n12745) );
  AOI21XL U26287 ( .A0(n12742), .A1(n12741), .B0(n12740), .Y(n12743) );
  OAI21XL U26288 ( .A0(n12745), .A1(n12744), .B0(n12743), .Y(n12842) );
  AOI21XL U26289 ( .A0(n12749), .A1(n12748), .B0(n12747), .Y(n12847) );
  NAND2XL U26290 ( .A(n12750), .B(U1_U2_y1[13]), .Y(n12852) );
  OAI21XL U26291 ( .A0(n12847), .A1(n12851), .B0(n12852), .Y(n12751) );
  AOI21XL U26292 ( .A0(n12752), .A1(n12842), .B0(n12751), .Y(n12753) );
  CMPR22X1 U26293 ( .A(U1_U2_y1[14]), .B(U1_U2_y0[14]), .CO(n12756), .S(n12750) );
  NOR2XL U26294 ( .A(n12872), .B(n12874), .Y(n12807) );
  CMPR22X1 U26295 ( .A(U1_U2_y1[17]), .B(U1_U2_y0[17]), .CO(n12762), .S(n12759) );
  INVXL U26296 ( .A(n12790), .Y(n12776) );
  CMPR22X1 U26297 ( .A(U1_U2_y1[18]), .B(U1_U2_y0[18]), .CO(n12765), .S(n12761) );
  INVXL U26298 ( .A(n12789), .Y(n12768) );
  XNOR2X2 U26299 ( .A(n12770), .B(n12769), .Y(n19519) );
  NAND2XL U26300 ( .A(n12771), .B(n12779), .Y(n12772) );
  INVXL U26301 ( .A(n14921), .Y(n12884) );
  INVXL U26302 ( .A(n12786), .Y(n12774) );
  NAND2XL U26303 ( .A(n12774), .B(n12788), .Y(n12775) );
  NOR2XL U26304 ( .A(n17708), .B(n17706), .Y(n17701) );
  NAND2XL U26305 ( .A(n12784), .B(n12919), .Y(n12785) );
  XOR2X1 U26306 ( .A(n12921), .B(n12785), .Y(n14923) );
  INVXL U26307 ( .A(n14923), .Y(n12886) );
  NAND2XL U26308 ( .A(n12793), .B(n12927), .Y(n12794) );
  NAND2XL U26309 ( .A(n17701), .B(n12795), .Y(n12889) );
  INVXL U26310 ( .A(n12796), .Y(n12799) );
  INVXL U26311 ( .A(n12797), .Y(n12798) );
  OAI21XL U26312 ( .A0(n7827), .A1(n12799), .B0(n12798), .Y(n12821) );
  INVXL U26313 ( .A(n12800), .Y(n12819) );
  AOI21XL U26314 ( .A0(n12821), .A1(n12819), .B0(n12801), .Y(n12806) );
  NAND2XL U26315 ( .A(n12804), .B(n12803), .Y(n12805) );
  XOR2X1 U26316 ( .A(n12806), .B(n12805), .Y(n14916) );
  INVXL U26317 ( .A(n14916), .Y(n12881) );
  INVXL U26318 ( .A(n12807), .Y(n12810) );
  INVXL U26319 ( .A(n12808), .Y(n12809) );
  OAI21XL U26320 ( .A0(n12873), .A1(n12810), .B0(n12809), .Y(n12825) );
  INVXL U26321 ( .A(n12811), .Y(n12823) );
  AOI21XL U26322 ( .A0(n12825), .A1(n12823), .B0(n12812), .Y(n12817) );
  NAND2XL U26323 ( .A(n12815), .B(n12814), .Y(n12816) );
  NOR2XL U26324 ( .A(n12881), .B(n19358), .Y(n17720) );
  XNOR2X1 U26325 ( .A(n12821), .B(n12820), .Y(n14915) );
  INVXL U26326 ( .A(n14915), .Y(n12880) );
  NAND2XL U26327 ( .A(n12823), .B(n12822), .Y(n12824) );
  NOR2XL U26328 ( .A(n12880), .B(n19363), .Y(n17726) );
  NOR2XL U26329 ( .A(n17720), .B(n17726), .Y(n12883) );
  INVXL U26330 ( .A(n12846), .Y(n12849) );
  INVXL U26331 ( .A(n12851), .Y(n12853) );
  NAND2XL U26332 ( .A(n12856), .B(n12864), .Y(n12857) );
  XOR2X1 U26333 ( .A(n7827), .B(n12857), .Y(n14907) );
  INVXL U26334 ( .A(n14907), .Y(n12861) );
  INVXL U26335 ( .A(n12872), .Y(n12858) );
  NAND2XL U26336 ( .A(n12858), .B(n12871), .Y(n12859) );
  XOR2X1 U26337 ( .A(n12873), .B(n12859), .Y(n19373) );
  NAND2XL U26338 ( .A(n12861), .B(n19373), .Y(n17738) );
  INVXL U26339 ( .A(n17738), .Y(n12862) );
  AOI21XL U26340 ( .A0(n12863), .A1(n12860), .B0(n12862), .Y(n17735) );
  OAI21XL U26341 ( .A0(n7827), .A1(n12865), .B0(n12864), .Y(n12870) );
  INVXL U26342 ( .A(n12866), .Y(n12868) );
  NAND2XL U26343 ( .A(n12868), .B(n12867), .Y(n12869) );
  INVXL U26344 ( .A(n14912), .Y(n12879) );
  OAI21XL U26345 ( .A0(n12873), .A1(n12872), .B0(n12871), .Y(n12878) );
  INVXL U26346 ( .A(n12874), .Y(n12876) );
  NOR2XL U26347 ( .A(n12879), .B(n19369), .Y(n17732) );
  NAND2XL U26348 ( .A(n12879), .B(n19369), .Y(n17733) );
  OAI21XL U26349 ( .A0(n17735), .A1(n17732), .B0(n17733), .Y(n17719) );
  NAND2XL U26350 ( .A(n12880), .B(n19363), .Y(n17727) );
  NAND2XL U26351 ( .A(n12881), .B(n19358), .Y(n17721) );
  OAI21XL U26352 ( .A0(n17720), .A1(n17727), .B0(n17721), .Y(n12882) );
  AOI21XL U26353 ( .A0(n12883), .A1(n17719), .B0(n12882), .Y(n17699) );
  NAND2XL U26354 ( .A(n12884), .B(n19518), .Y(n17714) );
  NAND2XL U26355 ( .A(n12885), .B(n19519), .Y(n17709) );
  OAI21XL U26356 ( .A0(n17708), .A1(n17714), .B0(n17709), .Y(n17700) );
  NAND2XL U26357 ( .A(n12886), .B(n19520), .Y(n17702) );
  INVXL U26358 ( .A(n12948), .Y(n12909) );
  INVXL U26359 ( .A(n12949), .Y(n12912) );
  NOR2X1 U26360 ( .A(n12965), .B(n19321), .Y(n17684) );
  XNOR2X1 U26361 ( .A(n7830), .B(n12916), .Y(n14933) );
  INVXL U26362 ( .A(n14933), .Y(n12964) );
  NAND2XL U26363 ( .A(n12917), .B(n12948), .Y(n12918) );
  NOR2XL U26364 ( .A(n12964), .B(n19326), .Y(n17682) );
  NOR2XL U26365 ( .A(n17684), .B(n17682), .Y(n12968) );
  OAI21XL U26366 ( .A0(n12921), .A1(n12920), .B0(n12919), .Y(n12926) );
  OAI21XL U26367 ( .A0(n12929), .A1(n12928), .B0(n12927), .Y(n12934) );
  INVXL U26368 ( .A(n12930), .Y(n12932) );
  NAND2XL U26369 ( .A(n12932), .B(n12931), .Y(n12933) );
  NOR2XL U26370 ( .A(n12963), .B(n19330), .Y(n17681) );
  INVXL U26371 ( .A(n17681), .Y(n12935) );
  NAND2XL U26372 ( .A(n12968), .B(n12935), .Y(n17668) );
  ADDHX2 U26373 ( .A(U1_U1_y2[24]), .B(U1_U1_y0[24]), .CO(n12941), .S(n12897)
         );
  INVXL U26374 ( .A(n12978), .Y(n12944) );
  NOR2X2 U26375 ( .A(n12951), .B(n12950), .Y(n12992) );
  OAI21X1 U26376 ( .A0(n12962), .A1(n12992), .B0(n12995), .Y(n12956) );
  CMPR22X1 U26377 ( .A(U1_U2_y1[25]), .B(U1_U2_y0[25]), .CO(n12953), .S(n12950) );
  INVXL U26378 ( .A(n12996), .Y(n12954) );
  OR2X2 U26379 ( .A(n12970), .B(n19532), .Y(n17671) );
  XOR2X2 U26380 ( .A(n12959), .B(n12958), .Y(n14940) );
  INVXL U26381 ( .A(n14940), .Y(n12969) );
  OR2X2 U26382 ( .A(n12969), .B(n19311), .Y(n17676) );
  NAND2XL U26383 ( .A(n12964), .B(n19326), .Y(n17690) );
  NAND2XL U26384 ( .A(n12965), .B(n19321), .Y(n17685) );
  OAI21XL U26385 ( .A0(n17684), .A1(n17690), .B0(n17685), .Y(n12966) );
  NAND2XL U26386 ( .A(n12969), .B(n19311), .Y(n17675) );
  INVXL U26387 ( .A(n17675), .Y(n17669) );
  NAND2XL U26388 ( .A(n12970), .B(n19532), .Y(n17670) );
  INVXL U26389 ( .A(n17670), .Y(n12971) );
  AOI21XL U26390 ( .A0(n17671), .A1(n17669), .B0(n12971), .Y(n12972) );
  CMPR22X1 U26391 ( .A(U1_U1_y2[27]), .B(U1_U1_y0[27]), .CO(n12985), .S(n12982) );
  NAND2X1 U26392 ( .A(n12990), .B(n13059), .Y(n12991) );
  OAI21X1 U26393 ( .A0(n12996), .A1(n12995), .B0(n12994), .Y(n12997) );
  CMPR22X1 U26394 ( .A(U1_U2_y1[29]), .B(U1_U2_y0[29]), .CO(n13007), .S(n13004) );
  INVXL U26395 ( .A(n13044), .Y(n13008) );
  NAND2XL U26396 ( .A(n13007), .B(n13006), .Y(n13042) );
  NOR2XL U26397 ( .A(n5862), .B(n19544), .Y(n17648) );
  INVXL U26398 ( .A(n17648), .Y(n13015) );
  INVXL U26399 ( .A(n13020), .Y(n13022) );
  XNOR2X2 U26400 ( .A(n13024), .B(n13023), .Y(n19542) );
  INVXL U26401 ( .A(n13026), .Y(n13028) );
  NAND2XL U26402 ( .A(n13025), .B(n13034), .Y(n17643) );
  NAND2XL U26403 ( .A(n5869), .B(n19542), .Y(n17658) );
  INVXL U26404 ( .A(n17658), .Y(n13036) );
  NAND2XL U26405 ( .A(n5862), .B(n19544), .Y(n17647) );
  INVXL U26406 ( .A(n17647), .Y(n13038) );
  ADDHX2 U26407 ( .A(U1_U2_y1[31]), .B(U1_U2_y0[31]), .CO(n13053), .S(n13049)
         );
  INVXL U26408 ( .A(n13074), .Y(n13054) );
  INVXL U26409 ( .A(n13081), .Y(n13068) );
  CMPR22X1 U26410 ( .A(U1_U2_y1[32]), .B(U1_U2_y0[32]), .CO(n13076), .S(n13052) );
  INVXL U26411 ( .A(n13564), .Y(n13087) );
  INVXL U26412 ( .A(n13577), .Y(n13085) );
  OR2X2 U26413 ( .A(n19553), .B(n5856), .Y(n17628) );
  INVXL U26414 ( .A(n13568), .Y(n13090) );
  NAND2X1 U26415 ( .A(n13090), .B(n13566), .Y(n13091) );
  NOR2X1 U26416 ( .A(n13093), .B(n13092), .Y(n13581) );
  INVXL U26417 ( .A(n13581), .Y(n13094) );
  NAND2XL U26418 ( .A(n13093), .B(n13092), .Y(n13579) );
  NAND2XL U26419 ( .A(n19259), .B(n5853), .Y(n14501) );
  MXI2X1 U26420 ( .A(U1_pipe11[20]), .B(n13096), .S0(n24784), .Y(n4886) );
  NOR2XL U26421 ( .A(n22885), .B(n13107), .Y(n22395) );
  NOR2XL U26422 ( .A(n22886), .B(n13106), .Y(n22393) );
  NOR2XL U26423 ( .A(n22395), .B(n22393), .Y(n22388) );
  NAND2XL U26424 ( .A(n22388), .B(n13097), .Y(n13111) );
  NOR2XL U26425 ( .A(n22889), .B(n13103), .Y(n22409) );
  NOR2XL U26426 ( .A(n22890), .B(n13102), .Y(n22408) );
  NOR2XL U26427 ( .A(n22409), .B(n22408), .Y(n13105) );
  NAND2XL U26428 ( .A(n22892), .B(n13099), .Y(n22097) );
  INVXL U26429 ( .A(n22097), .Y(n13100) );
  AOI21XL U26430 ( .A0(n22421), .A1(n5768), .B0(n13100), .Y(n22418) );
  NOR2XL U26431 ( .A(n22897), .B(n13101), .Y(n22091) );
  OAI21XL U26432 ( .A0(n22418), .A1(n22091), .B0(n22092), .Y(n22406) );
  NAND2XL U26433 ( .A(n22890), .B(n13102), .Y(n22407) );
  NAND2XL U26434 ( .A(n22889), .B(n13103), .Y(n22410) );
  OAI21XL U26435 ( .A0(n22409), .A1(n22407), .B0(n22410), .Y(n13104) );
  AOI21XL U26436 ( .A0(n13105), .A1(n22406), .B0(n13104), .Y(n22386) );
  NAND2XL U26437 ( .A(n22886), .B(n13106), .Y(n22401) );
  NAND2XL U26438 ( .A(n22885), .B(n13107), .Y(n22396) );
  OAI21XL U26439 ( .A0(n22395), .A1(n22401), .B0(n22396), .Y(n22387) );
  NAND2XL U26440 ( .A(n22887), .B(n13108), .Y(n22389) );
  INVXL U26441 ( .A(n22389), .Y(n13109) );
  AOI21XL U26442 ( .A0(n22387), .A1(n13097), .B0(n13109), .Y(n13110) );
  OAI21XL U26443 ( .A0(n13111), .A1(n22386), .B0(n13110), .Y(n22361) );
  NOR2XL U26444 ( .A(n22914), .B(n14530), .Y(n22050) );
  NOR2XL U26445 ( .A(n22915), .B(n13113), .Y(n22373) );
  INVXL U26446 ( .A(n22373), .Y(n22054) );
  NAND2XL U26447 ( .A(n13117), .B(n22054), .Y(n22363) );
  OR2X2 U26448 ( .A(n22917), .B(n14532), .Y(n22030) );
  NAND2X1 U26449 ( .A(n22030), .B(n22365), .Y(n13120) );
  NAND2XL U26450 ( .A(n22915), .B(n13113), .Y(n22372) );
  INVXL U26451 ( .A(n22372), .Y(n13116) );
  NAND2XL U26452 ( .A(n22914), .B(n14530), .Y(n22374) );
  NAND2XL U26453 ( .A(n22913), .B(n13114), .Y(n22045) );
  INVXL U26454 ( .A(n22034), .Y(n22364) );
  NAND2XL U26455 ( .A(n22917), .B(n14532), .Y(n22029) );
  INVXL U26456 ( .A(n22029), .Y(n13118) );
  NOR2XL U26457 ( .A(n22934), .B(n14547), .Y(n22341) );
  INVXL U26458 ( .A(n22341), .Y(n22347) );
  NAND2XL U26459 ( .A(n22353), .B(n13122), .Y(n22337) );
  NAND2XL U26460 ( .A(n22936), .B(n14548), .Y(n22357) );
  NAND2XL U26461 ( .A(n22935), .B(n13123), .Y(n22352) );
  INVXL U26462 ( .A(n22352), .Y(n13124) );
  NAND2XL U26463 ( .A(n22934), .B(n14547), .Y(n22346) );
  INVXL U26464 ( .A(n22346), .Y(n13127) );
  INVXL U26465 ( .A(n22342), .Y(n13126) );
  NAND2XL U26466 ( .A(n22930), .B(n13131), .Y(n21984) );
  INVXL U26467 ( .A(n21984), .Y(n13132) );
  OAI21X1 U26468 ( .A0(n13141), .A1(n13147), .B0(n13151), .Y(n13146) );
  CMPR22X1 U26469 ( .A(U0_U1_y2[34]), .B(U0_U1_y0[34]), .CO(n13143), .S(n12644) );
  NOR2XL U26470 ( .A(n22957), .B(n13166), .Y(n22310) );
  INVXL U26471 ( .A(n22310), .Y(n21974) );
  NAND2XL U26472 ( .A(n13155), .B(n13159), .Y(n13158) );
  NAND2XL U26473 ( .A(n21974), .B(n6987), .Y(n22305) );
  INVXL U26474 ( .A(n22309), .Y(n13169) );
  NAND2XL U26475 ( .A(n22958), .B(n13167), .Y(n21969) );
  INVXL U26476 ( .A(n21969), .Y(n13168) );
  NAND2XL U26477 ( .A(n22959), .B(n14570), .Y(n21962) );
  CMPR22X1 U26478 ( .A(U0_U1_y2[37]), .B(U0_U1_y0[37]), .CO(n13176), .S(n13162) );
  CMPR22X1 U26479 ( .A(U0_U1_y2[38]), .B(U0_U1_y0[38]), .CO(n13183), .S(n13175) );
  INVXL U26480 ( .A(n21948), .Y(n13185) );
  NAND2XL U26481 ( .A(n13192), .B(n22295), .Y(n13193) );
  MXI2X1 U26482 ( .A(U0_pipe5[26]), .B(n13194), .S0(n5812), .Y(n4492) );
  CMPR22X1 U26483 ( .A(U0_U0_y1[16]), .B(U0_U0_y0[16]), .CO(n13249), .S(n13246) );
  CMPR22X1 U26484 ( .A(U0_U0_y1[17]), .B(U0_U0_y0[17]), .CO(n13251), .S(n13248) );
  OR2XL U26485 ( .A(U0_U0_y1[1]), .B(U0_U0_y0[1]), .Y(n13196) );
  AOI21XL U26486 ( .A0(n13196), .A1(n7958), .B0(n13195), .Y(n13203) );
  NAND2XL U26487 ( .A(n13197), .B(n13200), .Y(n13202) );
  AOI21XL U26488 ( .A0(n13200), .A1(n13199), .B0(n13198), .Y(n13201) );
  OAI21XL U26489 ( .A0(n13203), .A1(n13202), .B0(n13201), .Y(n13219) );
  OR2X2 U26490 ( .A(U0_U0_y1[5]), .B(U0_U0_y0[5]), .Y(n13210) );
  NAND2XL U26491 ( .A(n13204), .B(n13210), .Y(n13207) );
  OR2X2 U26492 ( .A(U0_U0_y1[7]), .B(U0_U0_y0[7]), .Y(n13213) );
  NAND2XL U26493 ( .A(n13206), .B(n13213), .Y(n13215) );
  NOR2XL U26494 ( .A(n13207), .B(n13215), .Y(n13218) );
  AOI21XL U26495 ( .A0(n13210), .A1(n13209), .B0(n13208), .Y(n13216) );
  AOI21XL U26496 ( .A0(n13213), .A1(n13212), .B0(n13211), .Y(n13214) );
  OAI21XL U26497 ( .A0(n13216), .A1(n13215), .B0(n13214), .Y(n13217) );
  AOI21XL U26498 ( .A0(n13219), .A1(n13218), .B0(n13217), .Y(n13332) );
  NOR2XL U26499 ( .A(U0_U0_y1[12]), .B(U0_U0_y0[12]), .Y(n13220) );
  INVXL U26500 ( .A(n13220), .Y(n13221) );
  CMPR22X1 U26501 ( .A(U0_U0_y1[14]), .B(U0_U0_y0[14]), .CO(n13245), .S(n13239) );
  NOR2X1 U26502 ( .A(n13337), .B(n13342), .Y(n13241) );
  OAI21XL U26503 ( .A0(n13234), .A1(n13233), .B0(n13232), .Y(n13333) );
  AOI21X1 U26504 ( .A0(n13238), .A1(n13237), .B0(n13236), .Y(n13338) );
  NAND2XL U26505 ( .A(n13239), .B(U0_U0_y1[13]), .Y(n13343) );
  OAI21XL U26506 ( .A0(n13338), .A1(n13342), .B0(n13343), .Y(n13240) );
  NOR2X2 U26507 ( .A(n13266), .B(n13265), .Y(n13421) );
  NOR2X2 U26508 ( .A(n13268), .B(n13267), .Y(n13416) );
  ADDHX2 U26509 ( .A(U0_U0_y0[28]), .B(U0_U0_y1[28]), .CO(n13270), .S(n13267)
         );
  CMPR22X1 U26510 ( .A(U0_U0_y1[29]), .B(U0_U0_y0[29]), .CO(n13272), .S(n13269) );
  NOR2X2 U26511 ( .A(n13272), .B(n13271), .Y(n13405) );
  ADDHX2 U26512 ( .A(U0_U0_y1[31]), .B(U0_U0_y0[31]), .CO(n13276), .S(n13273)
         );
  NOR2X2 U26513 ( .A(n13446), .B(n13442), .Y(n13431) );
  ADDHX2 U26514 ( .A(U0_U0_y1[32]), .B(U0_U0_y0[32]), .CO(n13278), .S(n13275)
         );
  NOR2X2 U26515 ( .A(n13278), .B(n13277), .Y(n13437) );
  NOR2X1 U26516 ( .A(n13437), .B(n13432), .Y(n13282) );
  NAND2X1 U26517 ( .A(n13431), .B(n13282), .Y(n13468) );
  CMPR22X1 U26518 ( .A(U0_U0_y1[34]), .B(U0_U0_y0[34]), .CO(n13284), .S(n13279) );
  NAND2XL U26519 ( .A(n13264), .B(n13263), .Y(n13385) );
  NAND2XL U26520 ( .A(n13272), .B(n13271), .Y(n13406) );
  OAI21XL U26521 ( .A0(n13432), .A1(n13438), .B0(n13433), .Y(n13281) );
  NOR2X1 U26522 ( .A(n13290), .B(n13289), .Y(n13477) );
  CMPR22X1 U26523 ( .A(U0_U0_y1[37]), .B(U0_U0_y0[37]), .CO(n13293), .S(n13289) );
  CMPR22X1 U26524 ( .A(U0_U0_y1[38]), .B(U0_U0_y0[38]), .CO(n13296), .S(n13292) );
  INVXL U26525 ( .A(n13304), .Y(n13306) );
  NAND2XL U26526 ( .A(n13310), .B(n13309), .Y(n13311) );
  NOR2XL U26527 ( .A(n14065), .B(U2_A_r_d[5]), .Y(n24545) );
  NAND2XL U26528 ( .A(n13315), .B(n13373), .Y(n13316) );
  XOR2X1 U26529 ( .A(n13375), .B(n13316), .Y(n14025) );
  OR2X2 U26530 ( .A(n14067), .B(U2_A_r_d[7]), .Y(n24541) );
  INVXL U26531 ( .A(n13318), .Y(n13319) );
  OAI21XL U26532 ( .A0(n5903), .A1(n13320), .B0(n13319), .Y(n13331) );
  INVXL U26533 ( .A(n13328), .Y(n13322) );
  AOI21X1 U26534 ( .A0(n13331), .A1(n13329), .B0(n13322), .Y(n13327) );
  NAND2XL U26535 ( .A(n13329), .B(n13328), .Y(n13330) );
  XNOR2X1 U26536 ( .A(n13331), .B(n13330), .Y(n14021) );
  NOR2XL U26537 ( .A(n14062), .B(U2_A_r_d[3]), .Y(n24565) );
  INVX1 U26538 ( .A(n14016), .Y(n24581) );
  NOR2XL U26539 ( .A(n24581), .B(U2_A_r_d[0]), .Y(n24578) );
  NAND2XL U26540 ( .A(n13347), .B(n13352), .Y(n13348) );
  XOR2X1 U26541 ( .A(n5903), .B(n13348), .Y(n14018) );
  AND2XL U26542 ( .A(n14057), .B(U2_A_r_d[1]), .Y(n13349) );
  AOI21XL U26543 ( .A0(n13351), .A1(n13350), .B0(n13349), .Y(n24574) );
  OAI21XL U26544 ( .A0(n5903), .A1(n13353), .B0(n13352), .Y(n13358) );
  INVXL U26545 ( .A(n13354), .Y(n13356) );
  XNOR2X1 U26546 ( .A(n13358), .B(n13357), .Y(n14020) );
  NOR2XL U26547 ( .A(n14061), .B(U2_A_r_d[2]), .Y(n24571) );
  OAI21XL U26548 ( .A0(n24574), .A1(n24571), .B0(n24572), .Y(n24558) );
  NAND2XL U26549 ( .A(n14062), .B(U2_A_r_d[3]), .Y(n24566) );
  NAND2XL U26550 ( .A(n13359), .B(U2_A_r_d[4]), .Y(n24560) );
  OAI21XL U26551 ( .A0(n24559), .A1(n24566), .B0(n24560), .Y(n13360) );
  AOI21XL U26552 ( .A0(n13361), .A1(n24558), .B0(n13360), .Y(n24537) );
  AOI21XL U26553 ( .A0(n24538), .A1(n24541), .B0(n13362), .Y(n13363) );
  INVXL U26554 ( .A(n13366), .Y(n13368) );
  NOR2XL U26555 ( .A(n14076), .B(U2_A_r_d[10]), .Y(n13394) );
  NOR2XL U26556 ( .A(n5877), .B(U2_A_r_d[9]), .Y(n24519) );
  OAI21XL U26557 ( .A0(n13375), .A1(n13374), .B0(n13373), .Y(n13380) );
  INVXL U26558 ( .A(n13376), .Y(n13378) );
  INVX1 U26559 ( .A(n14030), .Y(n14075) );
  NOR2XL U26560 ( .A(n14075), .B(U2_A_r_d[8]), .Y(n24518) );
  INVXL U26561 ( .A(n24518), .Y(n13381) );
  NAND2XL U26562 ( .A(n13397), .B(n13381), .Y(n24505) );
  OR2X2 U26563 ( .A(n13398), .B(U2_A_r_d[12]), .Y(n13399) );
  OR2X2 U26564 ( .A(n5876), .B(U2_A_r_d[11]), .Y(n24507) );
  NAND2XL U26565 ( .A(n14075), .B(U2_A_r_d[8]), .Y(n24517) );
  INVXL U26566 ( .A(n24517), .Y(n13396) );
  NAND2XL U26567 ( .A(n5877), .B(U2_A_r_d[9]), .Y(n24520) );
  NAND2XL U26568 ( .A(n14076), .B(U2_A_r_d[10]), .Y(n13393) );
  OAI21XL U26569 ( .A0(n13394), .A1(n24520), .B0(n13393), .Y(n13395) );
  INVXL U26570 ( .A(n13405), .Y(n13407) );
  INVXL U26571 ( .A(n13408), .Y(n13455) );
  XOR2X2 U26572 ( .A(n13413), .B(n13412), .Y(n14042) );
  INVX1 U26573 ( .A(n14042), .Y(n14091) );
  NOR2XL U26574 ( .A(n14091), .B(U2_A_r_d[15]), .Y(n24482) );
  INVXL U26575 ( .A(n24482), .Y(n13414) );
  OAI21X1 U26576 ( .A0(n13425), .A1(n13421), .B0(n13422), .Y(n13420) );
  INVXL U26577 ( .A(n13416), .Y(n13418) );
  NAND2XL U26578 ( .A(n13423), .B(n13422), .Y(n13424) );
  INVX1 U26579 ( .A(n14040), .Y(n14088) );
  OR2X2 U26580 ( .A(n14088), .B(U2_A_r_d[13]), .Y(n24493) );
  NAND2XL U26581 ( .A(n13451), .B(n24493), .Y(n24477) );
  NOR2XL U26582 ( .A(n13457), .B(n24477), .Y(n24451) );
  INVXL U26583 ( .A(n13432), .Y(n13434) );
  NAND2X1 U26584 ( .A(n13434), .B(n13433), .Y(n13435) );
  XNOR2X4 U26585 ( .A(n13436), .B(n13435), .Y(n14053) );
  INVXL U26586 ( .A(n13437), .Y(n13439) );
  OR2X2 U26587 ( .A(n14103), .B(U2_A_r_d[19]), .Y(n24455) );
  NAND2X1 U26588 ( .A(n8078), .B(n24455), .Y(n13462) );
  INVXL U26589 ( .A(n13442), .Y(n13444) );
  NOR2XL U26590 ( .A(n14099), .B(U2_A_r_d[17]), .Y(n13449) );
  INVXL U26591 ( .A(n13449), .Y(n24467) );
  NAND2XL U26592 ( .A(n14091), .B(U2_A_r_d[15]), .Y(n24481) );
  INVXL U26593 ( .A(n24481), .Y(n13454) );
  AND2X1 U26594 ( .A(n13452), .B(U2_A_r_d[16]), .Y(n13453) );
  AND2X2 U26595 ( .A(n14099), .B(U2_A_r_d[17]), .Y(n24466) );
  AND2X2 U26596 ( .A(n14103), .B(U2_A_r_d[19]), .Y(n24454) );
  AND2X2 U26597 ( .A(n14133), .B(U2_A_r_d[20]), .Y(n13460) );
  OAI21X1 U26598 ( .A0(n24449), .A1(n13466), .B0(n13465), .Y(n24421) );
  NAND2X1 U26599 ( .A(n13472), .B(n13471), .Y(n13473) );
  INVX1 U26600 ( .A(n22448), .Y(n13486) );
  NOR2XL U26601 ( .A(n13486), .B(U2_A_r_d[21]), .Y(n24440) );
  INVX1 U26602 ( .A(n22452), .Y(n14150) );
  NOR2XL U26603 ( .A(n14150), .B(U2_A_r_d[23]), .Y(n13482) );
  INVXL U26604 ( .A(n13482), .Y(n13489) );
  NAND2XL U26605 ( .A(n24430), .B(n13489), .Y(n24423) );
  NAND2X1 U26606 ( .A(n13291), .B(n13483), .Y(n13484) );
  INVX2 U26607 ( .A(n22453), .Y(n14153) );
  NOR2XL U26608 ( .A(n14153), .B(U2_A_r_d[24]), .Y(n13491) );
  NOR2XL U26609 ( .A(n24423), .B(n13491), .Y(n13493) );
  NAND2XL U26610 ( .A(n14147), .B(U2_A_r_d[22]), .Y(n13487) );
  NAND2XL U26611 ( .A(n14153), .B(U2_A_r_d[24]), .Y(n13490) );
  NOR2XL U26612 ( .A(n14158), .B(U2_A_r_d[25]), .Y(n24416) );
  NAND2XL U26613 ( .A(n14158), .B(U2_A_r_d[25]), .Y(n24417) );
  MXI2X1 U26614 ( .A(U0_pipe2[26]), .B(n13499), .S0(n22853), .Y(n4377) );
  NOR2XL U26615 ( .A(n24953), .B(n24951), .Y(n24945) );
  OR2X2 U26616 ( .A(n14025), .B(U2_A_r_d[7]), .Y(n24947) );
  NAND2XL U26617 ( .A(n24945), .B(n24947), .Y(n13505) );
  NOR2XL U26618 ( .A(n14056), .B(U2_A_r_d[4]), .Y(n24965) );
  NOR2XL U26619 ( .A(n14021), .B(U2_A_r_d[3]), .Y(n24971) );
  NOR2XL U26620 ( .A(n24965), .B(n24971), .Y(n13502) );
  NAND2XL U26621 ( .A(n14018), .B(U2_A_r_d[1]), .Y(n24577) );
  INVXL U26622 ( .A(n24577), .Y(n13500) );
  AOI21XL U26623 ( .A0(n24983), .A1(n5778), .B0(n13500), .Y(n24980) );
  NOR2XL U26624 ( .A(n14020), .B(U2_A_r_d[2]), .Y(n24977) );
  OAI21XL U26625 ( .A0(n24980), .A1(n24977), .B0(n24978), .Y(n24964) );
  NAND2XL U26626 ( .A(n14021), .B(U2_A_r_d[3]), .Y(n24972) );
  NAND2XL U26627 ( .A(n14056), .B(U2_A_r_d[4]), .Y(n24966) );
  OAI21XL U26628 ( .A0(n24965), .A1(n24972), .B0(n24966), .Y(n13501) );
  AOI21XL U26629 ( .A0(n13502), .A1(n24964), .B0(n13501), .Y(n24943) );
  NAND2XL U26630 ( .A(n14024), .B(U2_A_r_d[5]), .Y(n24959) );
  OAI21XL U26631 ( .A0(n24953), .A1(n24959), .B0(n24954), .Y(n24944) );
  AOI21XL U26632 ( .A0(n24944), .A1(n24947), .B0(n13503), .Y(n13504) );
  NOR2X1 U26633 ( .A(n14031), .B(U2_A_r_d[10]), .Y(n24523) );
  NOR2XL U26634 ( .A(n14071), .B(U2_A_r_d[9]), .Y(n24529) );
  NAND2XL U26635 ( .A(n13510), .B(n24533), .Y(n24921) );
  NAND2XL U26636 ( .A(n14030), .B(U2_A_r_d[8]), .Y(n24929) );
  INVXL U26637 ( .A(n24929), .Y(n13509) );
  NAND2XL U26638 ( .A(n14071), .B(U2_A_r_d[9]), .Y(n24931) );
  NAND2XL U26639 ( .A(n14031), .B(U2_A_r_d[10]), .Y(n24524) );
  OAI21XL U26640 ( .A0(n24523), .A1(n24931), .B0(n24524), .Y(n13508) );
  INVXL U26641 ( .A(n24513), .Y(n24922) );
  INVXL U26642 ( .A(n24508), .Y(n13511) );
  OR2X2 U26643 ( .A(n14086), .B(U2_A_r_d[16]), .Y(n24484) );
  NOR2XL U26644 ( .A(n14042), .B(U2_A_r_d[15]), .Y(n24904) );
  OR2X2 U26645 ( .A(n14040), .B(U2_A_r_d[13]), .Y(n24912) );
  NAND2XL U26646 ( .A(n24495), .B(n24912), .Y(n24899) );
  NOR2X1 U26647 ( .A(n13518), .B(n24899), .Y(n13997) );
  NOR2XL U26648 ( .A(n14102), .B(U2_A_r_d[19]), .Y(n14002) );
  NOR2XL U26649 ( .A(n14047), .B(U2_A_r_d[17]), .Y(n24891) );
  NAND2XL U26650 ( .A(n14040), .B(U2_A_r_d[13]), .Y(n24499) );
  INVXL U26651 ( .A(n24499), .Y(n24911) );
  INVXL U26652 ( .A(n24494), .Y(n13514) );
  AOI21XL U26653 ( .A0(n24495), .A1(n24911), .B0(n13514), .Y(n24900) );
  NAND2XL U26654 ( .A(n14042), .B(U2_A_r_d[15]), .Y(n24903) );
  INVXL U26655 ( .A(n24903), .Y(n13516) );
  NAND2XL U26656 ( .A(n14086), .B(U2_A_r_d[16]), .Y(n24483) );
  INVXL U26657 ( .A(n24483), .Y(n13515) );
  AOI21XL U26658 ( .A0(n24484), .A1(n13516), .B0(n13515), .Y(n13517) );
  NAND2X1 U26659 ( .A(n14047), .B(U2_A_r_d[17]), .Y(n24890) );
  NAND2XL U26660 ( .A(n14048), .B(U2_A_r_d[18]), .Y(n24468) );
  INVXL U26661 ( .A(n24468), .Y(n13519) );
  NAND2XL U26662 ( .A(n14102), .B(U2_A_r_d[19]), .Y(n24460) );
  INVXL U26663 ( .A(n24460), .Y(n13522) );
  NAND2XL U26664 ( .A(n14053), .B(U2_A_r_d[20]), .Y(n14003) );
  INVXL U26665 ( .A(n14003), .Y(n13521) );
  AOI21X1 U26666 ( .A0(n6995), .A1(n13522), .B0(n13521), .Y(n13523) );
  NAND2XL U26667 ( .A(n24445), .B(n13527), .Y(n24875) );
  NAND2X1 U26668 ( .A(n22448), .B(U2_A_r_d[21]), .Y(n24879) );
  INVXL U26669 ( .A(n24879), .Y(n13529) );
  NAND2XL U26670 ( .A(n22449), .B(U2_A_r_d[22]), .Y(n24441) );
  INVXL U26671 ( .A(n24441), .Y(n13528) );
  AOI21XL U26672 ( .A0(n13529), .A1(n13527), .B0(n13528), .Y(n24874) );
  NOR2X1 U26673 ( .A(n22453), .B(U2_A_r_d[24]), .Y(n24424) );
  OR2X2 U26674 ( .A(n22454), .B(U2_A_r_d[25]), .Y(n24866) );
  NOR2XL U26675 ( .A(n22456), .B(n29010), .Y(n24861) );
  INVXL U26676 ( .A(n24861), .Y(n13531) );
  MXI2X1 U26677 ( .A(U0_pipe0[26]), .B(n13533), .S0(n5812), .Y(n4286) );
  NOR2XL U26678 ( .A(n19519), .B(n14922), .Y(n17412) );
  NOR2XL U26679 ( .A(n17412), .B(n17410), .Y(n17405) );
  NAND2XL U26680 ( .A(n17405), .B(n13534), .Y(n13544) );
  NOR2XL U26681 ( .A(n19373), .B(n14907), .Y(n17436) );
  INVXL U26682 ( .A(n17436), .Y(n17442) );
  NAND2XL U26683 ( .A(n13535), .B(n17442), .Y(n13539) );
  NAND2XL U26684 ( .A(n19373), .B(n14907), .Y(n17441) );
  INVXL U26685 ( .A(n17441), .Y(n13537) );
  NAND2XL U26686 ( .A(n19369), .B(n14912), .Y(n17437) );
  INVXL U26687 ( .A(n17437), .Y(n13536) );
  AOI21XL U26688 ( .A0(n13535), .A1(n13537), .B0(n13536), .Y(n13538) );
  NOR2XL U26689 ( .A(n19358), .B(n14916), .Y(n17424) );
  NOR2XL U26690 ( .A(n19363), .B(n14915), .Y(n17430) );
  NOR2XL U26691 ( .A(n17424), .B(n17430), .Y(n13541) );
  NAND2XL U26692 ( .A(n19363), .B(n14915), .Y(n17431) );
  NAND2XL U26693 ( .A(n19358), .B(n14916), .Y(n17425) );
  OAI21XL U26694 ( .A0(n17424), .A1(n17431), .B0(n17425), .Y(n13540) );
  AOI21XL U26695 ( .A0(n17423), .A1(n13541), .B0(n13540), .Y(n17403) );
  NAND2XL U26696 ( .A(n19518), .B(n14921), .Y(n17418) );
  NAND2XL U26697 ( .A(n19519), .B(n14922), .Y(n17413) );
  OAI21XL U26698 ( .A0(n17412), .A1(n17418), .B0(n17413), .Y(n17404) );
  NAND2XL U26699 ( .A(n19520), .B(n14923), .Y(n17406) );
  INVXL U26700 ( .A(n17406), .Y(n13542) );
  AOI21XL U26701 ( .A0(n17404), .A1(n13534), .B0(n13542), .Y(n13543) );
  NOR2XL U26702 ( .A(n14933), .B(n19326), .Y(n17386) );
  NOR2XL U26703 ( .A(n17388), .B(n17386), .Y(n13548) );
  NOR2XL U26704 ( .A(n19330), .B(n14932), .Y(n17385) );
  INVXL U26705 ( .A(n17385), .Y(n17400) );
  NAND2XL U26706 ( .A(n13548), .B(n17400), .Y(n17374) );
  OR2X2 U26707 ( .A(n14941), .B(n19532), .Y(n17377) );
  NAND2XL U26708 ( .A(n17377), .B(n13545), .Y(n13551) );
  NAND2XL U26709 ( .A(n19330), .B(n14932), .Y(n17399) );
  INVXL U26710 ( .A(n17399), .Y(n13547) );
  NAND2XL U26711 ( .A(n14933), .B(n19326), .Y(n17394) );
  OAI21XL U26712 ( .A0(n17388), .A1(n17394), .B0(n17389), .Y(n13546) );
  NAND2XL U26713 ( .A(n14940), .B(n19311), .Y(n17381) );
  INVXL U26714 ( .A(n17381), .Y(n17375) );
  NAND2XL U26715 ( .A(n14941), .B(n19532), .Y(n17376) );
  INVXL U26716 ( .A(n17376), .Y(n13549) );
  AOI21XL U26717 ( .A0(n17377), .A1(n17375), .B0(n13549), .Y(n13550) );
  OAI21XL U26718 ( .A0(n17373), .A1(n13551), .B0(n13550), .Y(n13552) );
  NOR2X1 U26719 ( .A(n19553), .B(n14959), .Y(n17328) );
  INVXL U26720 ( .A(n17328), .Y(n17335) );
  NAND2XL U26721 ( .A(n17364), .B(n13554), .Y(n17349) );
  NOR2X1 U26722 ( .A(n13557), .B(n17349), .Y(n17323) );
  NAND2XL U26723 ( .A(n14950), .B(n19541), .Y(n17368) );
  INVXL U26724 ( .A(n17368), .Y(n17362) );
  NAND2XL U26725 ( .A(n14951), .B(n19542), .Y(n17363) );
  INVXL U26726 ( .A(n17363), .Y(n13555) );
  NAND2XL U26727 ( .A(n14954), .B(n19282), .Y(n17354) );
  INVXL U26728 ( .A(n17354), .Y(n13556) );
  NAND2XL U26729 ( .A(n19272), .B(n14955), .Y(n17344) );
  INVXL U26730 ( .A(n17344), .Y(n13559) );
  INVXL U26731 ( .A(n17340), .Y(n13558) );
  AOI21X1 U26732 ( .A0(n17341), .A1(n13559), .B0(n13558), .Y(n17325) );
  NAND2XL U26733 ( .A(n19259), .B(n14960), .Y(n17329) );
  INVXL U26734 ( .A(n17329), .Y(n13560) );
  INVXL U26735 ( .A(n13598), .Y(n13572) );
  INVXL U26736 ( .A(n13602), .Y(n13571) );
  CMPR22X1 U26737 ( .A(U1_U2_y1[34]), .B(U1_U2_y0[34]), .CO(n13575), .S(n13088) );
  NOR2X1 U26738 ( .A(n13577), .B(n13581), .Y(n13584) );
  CMPR22X1 U26739 ( .A(U1_U1_y2[34]), .B(U1_U1_y0[34]), .CO(n13587), .S(n13092) );
  NOR2XL U26740 ( .A(n19557), .B(n14962), .Y(n17312) );
  INVXL U26741 ( .A(n17312), .Y(n17318) );
  CMPR22X1 U26742 ( .A(U1_U1_y2[35]), .B(U1_U1_y0[35]), .CO(n13597), .S(n13586) );
  CMPR22X1 U26743 ( .A(U1_U1_y2[36]), .B(U1_U1_y0[36]), .CO(n13611), .S(n13596) );
  NOR2X1 U26744 ( .A(n13611), .B(n13610), .Y(n13626) );
  NAND2X1 U26745 ( .A(n13612), .B(n13625), .Y(n13613) );
  CMPR22X1 U26746 ( .A(U1_U2_y1[36]), .B(U1_U2_y0[36]), .CO(n13618), .S(n13605) );
  NAND2XL U26747 ( .A(n19557), .B(n14962), .Y(n17317) );
  INVXL U26748 ( .A(n17317), .Y(n13622) );
  NAND2XL U26749 ( .A(n14963), .B(n19248), .Y(n17313) );
  INVXL U26750 ( .A(n17313), .Y(n13621) );
  CMPR22X1 U26751 ( .A(U1_U1_y2[37]), .B(U1_U1_y0[37]), .CO(n13630), .S(n13610) );
  CMPR22X1 U26752 ( .A(U1_U2_y1[37]), .B(U1_U2_y0[37]), .CO(n13636), .S(n13617) );
  CMPR22X1 U26753 ( .A(U1_U1_y2[38]), .B(U1_U1_y0[38]), .CO(n13641), .S(n13629) );
  CMPR22X1 U26754 ( .A(U1_U2_y1[38]), .B(U1_U2_y0[38]), .CO(n13648), .S(n13635) );
  NOR2X1 U26755 ( .A(n13648), .B(n13647), .Y(n13659) );
  NAND2X1 U26756 ( .A(n13649), .B(n13658), .Y(n13650) );
  OR2X2 U26757 ( .A(n14972), .B(n19233), .Y(n17297) );
  NAND2XL U26758 ( .A(n14972), .B(n19233), .Y(n17296) );
  XOR2X1 U26759 ( .A(n13656), .B(n13655), .Y(n13657) );
  XOR2X1 U26760 ( .A(n13662), .B(n13661), .Y(n13663) );
  NOR2XL U26761 ( .A(n19197), .B(n19203), .Y(n19476) );
  NAND2XL U26762 ( .A(n19476), .B(n13664), .Y(n13679) );
  NOR2XL U26763 ( .A(n19210), .B(n19491), .Y(n13673) );
  NAND2XL U26764 ( .A(n13667), .B(U1_A_r_d0[1]), .Y(n19227) );
  INVXL U26765 ( .A(n19227), .Y(n13668) );
  AOI21XL U26766 ( .A0(n19501), .A1(n13666), .B0(n13668), .Y(n19498) );
  OAI21XL U26767 ( .A0(n19498), .A1(n19221), .B0(n19222), .Y(n19489) );
  NAND2XL U26768 ( .A(n13671), .B(U1_A_r_d0[4]), .Y(n19211) );
  AOI21XL U26769 ( .A0(n13673), .A1(n19489), .B0(n13672), .Y(n19474) );
  NAND2XL U26770 ( .A(n13674), .B(U1_A_r_d0[5]), .Y(n19480) );
  NAND2XL U26771 ( .A(n13675), .B(U1_A_r_d0[6]), .Y(n19198) );
  OAI21XL U26772 ( .A0(n19197), .A1(n19480), .B0(n19198), .Y(n19475) );
  NAND2XL U26773 ( .A(n13676), .B(U1_A_r_d0[7]), .Y(n19189) );
  INVXL U26774 ( .A(n19189), .Y(n13677) );
  AOI21XL U26775 ( .A0(n19475), .A1(n13664), .B0(n13677), .Y(n13678) );
  OAI21XL U26776 ( .A0(n13679), .A1(n19474), .B0(n13678), .Y(n19450) );
  NOR2XL U26777 ( .A(n13682), .B(U1_A_r_d0[9]), .Y(n19178) );
  NOR2XL U26778 ( .A(n19172), .B(n19178), .Y(n13686) );
  NOR2XL U26779 ( .A(n13681), .B(U1_A_r_d0[8]), .Y(n19461) );
  INVXL U26780 ( .A(n19461), .Y(n19182) );
  NAND2XL U26781 ( .A(n13686), .B(n19182), .Y(n19452) );
  NAND2XL U26782 ( .A(n13681), .B(U1_A_r_d0[8]), .Y(n19460) );
  INVXL U26783 ( .A(n19460), .Y(n13685) );
  NAND2XL U26784 ( .A(n13682), .B(U1_A_r_d0[9]), .Y(n19462) );
  NAND2XL U26785 ( .A(n13683), .B(U1_A_r_d0[10]), .Y(n19173) );
  NAND2XL U26786 ( .A(n13687), .B(U1_A_r_d0[11]), .Y(n19162) );
  INVXL U26787 ( .A(n19162), .Y(n19453) );
  INVXL U26788 ( .A(n19157), .Y(n13688) );
  AOI21XL U26789 ( .A0(n19158), .A1(n19453), .B0(n13688), .Y(n13689) );
  NOR2XL U26790 ( .A(n13694), .B(U1_A_r_d0[15]), .Y(n19436) );
  INVXL U26791 ( .A(n19436), .Y(n19138) );
  OR2X2 U26792 ( .A(n13691), .B(U1_A_r_d0[13]), .Y(n19444) );
  NOR2X1 U26793 ( .A(n13697), .B(n19431), .Y(n19409) );
  OR2X2 U26794 ( .A(n13699), .B(U1_A_r_d0[18]), .Y(n19118) );
  NAND2XL U26795 ( .A(n13691), .B(U1_A_r_d0[13]), .Y(n19148) );
  INVXL U26796 ( .A(n19148), .Y(n19443) );
  NAND2XL U26797 ( .A(n13692), .B(U1_A_r_d0[14]), .Y(n19144) );
  INVXL U26798 ( .A(n19144), .Y(n13693) );
  INVXL U26799 ( .A(n19435), .Y(n13695) );
  OAI21X1 U26800 ( .A0(n13697), .A1(n19432), .B0(n13696), .Y(n19408) );
  NAND2X1 U26801 ( .A(n13698), .B(U1_A_r_d0[17]), .Y(n19422) );
  INVXL U26802 ( .A(n19422), .Y(n13701) );
  NAND2XL U26803 ( .A(n13699), .B(U1_A_r_d0[18]), .Y(n19119) );
  INVXL U26804 ( .A(n19119), .Y(n13700) );
  INVXL U26805 ( .A(n19414), .Y(n13704) );
  NAND2XL U26806 ( .A(n7696), .B(U1_A_r_d0[20]), .Y(n19108) );
  INVXL U26807 ( .A(n19108), .Y(n13703) );
  NOR2XL U26808 ( .A(n13709), .B(U1_A_r_d0[21]), .Y(n19399) );
  INVXL U26809 ( .A(n19399), .Y(n19098) );
  OR2X2 U26810 ( .A(n13710), .B(U1_A_r_d0[22]), .Y(n19094) );
  NAND2XL U26811 ( .A(n19098), .B(n19094), .Y(n19394) );
  NAND2X1 U26812 ( .A(n13709), .B(U1_A_r_d0[21]), .Y(n19398) );
  INVXL U26813 ( .A(n19398), .Y(n13712) );
  INVXL U26814 ( .A(n19093), .Y(n13711) );
  AOI21X1 U26815 ( .A0(n13712), .A1(n19094), .B0(n13711), .Y(n19393) );
  NAND2XL U26816 ( .A(n13713), .B(U1_A_r_d0[23]), .Y(n19086) );
  OR2X2 U26817 ( .A(n13717), .B(U1_A_r_d0[25]), .Y(n14895) );
  NAND2XL U26818 ( .A(n13717), .B(U1_A_r_d0[25]), .Y(n14893) );
  XNOR2X1 U26819 ( .A(n14896), .B(n19069), .Y(n13718) );
  INVXL U26820 ( .A(n13722), .Y(n13725) );
  INVXL U26821 ( .A(n13723), .Y(n13724) );
  OAI21XL U26822 ( .A0(n17200), .A1(n13726), .B0(n17198), .Y(n13729) );
  MXI2X1 U26823 ( .A(U1_pipe14[20]), .B(n13730), .S0(n5812), .Y(n4771) );
  NOR2XL U26824 ( .A(U1_U2_y2[1]), .B(U1_U2_y0[1]), .Y(n13731) );
  INVXL U26825 ( .A(n13731), .Y(n13734) );
  AND2XL U26826 ( .A(U1_U2_y2[0]), .B(U1_U2_y0[0]), .Y(n13733) );
  NOR2XL U26827 ( .A(U1_U2_y2[2]), .B(U1_U2_y0[2]), .Y(n13735) );
  INVXL U26828 ( .A(n13735), .Y(n13737) );
  NAND2XL U26829 ( .A(n13737), .B(n13739), .Y(n13741) );
  OAI21XL U26830 ( .A0(n13742), .A1(n13741), .B0(n13740), .Y(n13758) );
  OR2X1 U26831 ( .A(U1_U2_y2[6]), .B(U1_U2_y0[6]), .Y(n13746) );
  AOI21XL U26832 ( .A0(n13752), .A1(n13751), .B0(n13750), .Y(n13753) );
  OAI21XL U26833 ( .A0(n13755), .A1(n13754), .B0(n13753), .Y(n13756) );
  AOI21XL U26834 ( .A0(n13758), .A1(n13757), .B0(n13756), .Y(n13817) );
  OR2X2 U26835 ( .A(U1_U2_y2[12]), .B(U1_U2_y0[12]), .Y(n13759) );
  AOI21XL U26836 ( .A0(n13762), .A1(n7957), .B0(n13767), .Y(n13768) );
  OAI21XL U26837 ( .A0(n13770), .A1(n13769), .B0(n13768), .Y(n13818) );
  AOI21XL U26838 ( .A0(n13773), .A1(n13772), .B0(n7971), .Y(n13823) );
  NAND2XL U26839 ( .A(n13774), .B(U1_U2_y2[13]), .Y(n13827) );
  CMPR22X1 U26840 ( .A(U1_U2_y2[14]), .B(U1_U2_y0[14]), .CO(n13776), .S(n13774) );
  CMPR22X1 U26841 ( .A(U1_U2_y2[16]), .B(U1_U2_y0[16]), .CO(n13780), .S(n13777) );
  OAI21XL U26842 ( .A0(n13791), .A1(n13792), .B0(n13794), .Y(n13788) );
  CMPR22X1 U26843 ( .A(U1_U2_y2[19]), .B(U1_U2_y0[19]), .CO(n13786), .S(n13783) );
  INVXL U26844 ( .A(n13795), .Y(n13787) );
  INVXL U26845 ( .A(n13792), .Y(n13789) );
  NAND2XL U26846 ( .A(n13789), .B(n13794), .Y(n13790) );
  NOR2XL U26847 ( .A(n14921), .B(n14901), .Y(n17138) );
  NOR2X1 U26848 ( .A(n17140), .B(n17138), .Y(n17133) );
  CMPR22X1 U26849 ( .A(U1_U2_y2[20]), .B(U1_U2_y0[20]), .CO(n13798), .S(n13785) );
  NAND2XL U26850 ( .A(n13799), .B(n13862), .Y(n13800) );
  XOR2X1 U26851 ( .A(n13864), .B(n13800), .Y(n14902) );
  NAND2XL U26852 ( .A(n17133), .B(n13801), .Y(n13846) );
  INVXL U26853 ( .A(n13802), .Y(n13805) );
  INVXL U26854 ( .A(n13803), .Y(n13804) );
  OAI21XL U26855 ( .A0(n7046), .A1(n13805), .B0(n13804), .Y(n13816) );
  INVXL U26856 ( .A(n13806), .Y(n13814) );
  INVXL U26857 ( .A(n13813), .Y(n13807) );
  AOI21XL U26858 ( .A0(n13816), .A1(n13814), .B0(n13807), .Y(n13812) );
  NAND2XL U26859 ( .A(n13810), .B(n13809), .Y(n13811) );
  NOR2XL U26860 ( .A(n14916), .B(n19951), .Y(n16912) );
  NAND2XL U26861 ( .A(n13814), .B(n13813), .Y(n13815) );
  NOR2XL U26862 ( .A(n14915), .B(n14904), .Y(n17153) );
  NOR2XL U26863 ( .A(n16912), .B(n17153), .Y(n13843) );
  INVXL U26864 ( .A(n13836), .Y(n13831) );
  NAND2XL U26865 ( .A(n13831), .B(n13835), .Y(n13832) );
  XOR2X1 U26866 ( .A(n7046), .B(n13832), .Y(n19952) );
  NAND2XL U26867 ( .A(n14907), .B(n19952), .Y(n16928) );
  INVXL U26868 ( .A(n16928), .Y(n13834) );
  OAI21XL U26869 ( .A0(n7046), .A1(n13836), .B0(n13835), .Y(n13841) );
  INVXL U26870 ( .A(n13837), .Y(n13839) );
  NOR2XL U26871 ( .A(n14912), .B(n14911), .Y(n16922) );
  NAND2XL U26872 ( .A(n14912), .B(n14911), .Y(n16923) );
  OAI21XL U26873 ( .A0(n17160), .A1(n16922), .B0(n16923), .Y(n17151) );
  NAND2XL U26874 ( .A(n14915), .B(n14904), .Y(n17152) );
  NAND2XL U26875 ( .A(n14916), .B(n19951), .Y(n16913) );
  OAI21XL U26876 ( .A0(n16912), .A1(n17152), .B0(n16913), .Y(n13842) );
  AOI21XL U26877 ( .A0(n13843), .A1(n17151), .B0(n13842), .Y(n17131) );
  NAND2XL U26878 ( .A(n14921), .B(n14901), .Y(n17146) );
  NAND2XL U26879 ( .A(n14922), .B(n14900), .Y(n17141) );
  OAI21XL U26880 ( .A0(n17140), .A1(n17146), .B0(n17141), .Y(n17132) );
  NAND2XL U26881 ( .A(n14923), .B(n14902), .Y(n17134) );
  INVXL U26882 ( .A(n17134), .Y(n13844) );
  AOI21XL U26883 ( .A0(n17132), .A1(n13801), .B0(n13844), .Y(n13845) );
  ADDHX2 U26884 ( .A(U1_U2_y0[21]), .B(U1_U2_y2[21]), .CO(n13850), .S(n13797)
         );
  NOR2X1 U26885 ( .A(n14935), .B(n14926), .Y(n16875) );
  NOR2XL U26886 ( .A(n14933), .B(n19974), .Y(n16881) );
  NOR2XL U26887 ( .A(n16875), .B(n16881), .Y(n13884) );
  OAI21XL U26888 ( .A0(n13864), .A1(n13863), .B0(n13862), .Y(n13869) );
  NOR2XL U26889 ( .A(n14932), .B(n14927), .Y(n17118) );
  INVXL U26890 ( .A(n17118), .Y(n16885) );
  NAND2XL U26891 ( .A(n13884), .B(n16885), .Y(n17109) );
  CMPR22X1 U26892 ( .A(U1_U2_y2[24]), .B(U1_U2_y0[24]), .CO(n13875), .S(n13856) );
  NOR2X2 U26893 ( .A(n13875), .B(n13874), .Y(n13890) );
  CMPR22X1 U26894 ( .A(U1_U2_y2[25]), .B(U1_U2_y0[25]), .CO(n13876), .S(n13874) );
  INVXL U26895 ( .A(n13894), .Y(n13877) );
  NAND2XL U26896 ( .A(n14933), .B(n19974), .Y(n17119) );
  NAND2XL U26897 ( .A(n14935), .B(n14926), .Y(n16876) );
  OAI21XL U26898 ( .A0(n16875), .A1(n17119), .B0(n16876), .Y(n13882) );
  NAND2XL U26899 ( .A(n14940), .B(n14930), .Y(n16865) );
  INVXL U26900 ( .A(n16865), .Y(n17110) );
  NAND2XL U26901 ( .A(n14941), .B(n14929), .Y(n16861) );
  INVXL U26902 ( .A(n16861), .Y(n13885) );
  NAND2X1 U26903 ( .A(n6941), .B(n17093), .Y(n13945) );
  INVXL U26904 ( .A(n13909), .Y(n13911) );
  INVXL U26905 ( .A(n13913), .Y(n13915) );
  INVXL U26906 ( .A(n13953), .Y(n13932) );
  NAND2XL U26907 ( .A(n14951), .B(n19994), .Y(n17098) );
  NAND2XL U26908 ( .A(n14953), .B(n14945), .Y(n17092) );
  INVXL U26909 ( .A(n17092), .Y(n13943) );
  NAND2X1 U26910 ( .A(n14954), .B(n19993), .Y(n17088) );
  INVXL U26911 ( .A(n17088), .Y(n13942) );
  AOI21X1 U26912 ( .A0(n6941), .A1(n13943), .B0(n13942), .Y(n13944) );
  NAND2X1 U26913 ( .A(n14959), .B(n19996), .Y(n16818) );
  INVXL U26914 ( .A(n16818), .Y(n13947) );
  NAND2XL U26915 ( .A(n14960), .B(n14948), .Y(n14012) );
  INVXL U26916 ( .A(n14012), .Y(n13946) );
  CMPR22X1 U26917 ( .A(U1_U2_y2[34]), .B(U1_U2_y0[34]), .CO(n13957), .S(n13930) );
  NAND2X1 U26918 ( .A(n5879), .B(n13961), .Y(n13958) );
  NOR2XL U26919 ( .A(n14962), .B(n20050), .Y(n17064) );
  CMPR22X1 U26920 ( .A(U1_U2_y2[36]), .B(U1_U2_y0[36]), .CO(n13972), .S(n13964) );
  NAND2XL U26921 ( .A(n14963), .B(n20047), .Y(n16801) );
  INVXL U26922 ( .A(n16801), .Y(n13974) );
  CMPR22X1 U26923 ( .A(U1_U2_y2[37]), .B(U1_U2_y0[37]), .CO(n13979), .S(n13971) );
  INVX1 U26924 ( .A(n13980), .Y(n13981) );
  CMPR22X1 U26925 ( .A(U1_U2_y2[38]), .B(U1_U2_y0[38]), .CO(n13985), .S(n13978) );
  NAND2XL U26926 ( .A(n14972), .B(n20028), .Y(n17051) );
  INVXL U26927 ( .A(n17051), .Y(n13988) );
  INVXL U26928 ( .A(n17050), .Y(n13994) );
  INVXL U26929 ( .A(n13998), .Y(n14001) );
  INVXL U26930 ( .A(n13999), .Y(n14000) );
  AOI21X1 U26931 ( .A0(n24897), .A1(n14001), .B0(n14000), .Y(n24888) );
  XNOR2X1 U26932 ( .A(n14004), .B(n24456), .Y(n14005) );
  MXI2X1 U26933 ( .A(U0_pipe0[20]), .B(n14005), .S0(n5812), .Y(n4292) );
  XNOR2X1 U26934 ( .A(n14013), .B(n16814), .Y(n14014) );
  MXI2X1 U26935 ( .A(U1_pipe5[20]), .B(n14014), .S0(n5812), .Y(n4917) );
  NAND2XL U26936 ( .A(n22551), .B(n14015), .Y(n14028) );
  NOR2XL U26937 ( .A(n14056), .B(U2_A_i_d[4]), .Y(n22570) );
  NOR2XL U26938 ( .A(n14021), .B(U2_A_i_d[3]), .Y(n22576) );
  NOR2XL U26939 ( .A(n22570), .B(n22576), .Y(n14023) );
  NAND2XL U26940 ( .A(n14018), .B(U2_A_i_d[1]), .Y(n22588) );
  INVXL U26941 ( .A(n22588), .Y(n14019) );
  AOI21XL U26942 ( .A0(n22589), .A1(n14017), .B0(n14019), .Y(n22585) );
  NOR2XL U26943 ( .A(n14020), .B(U2_A_i_d[2]), .Y(n22582) );
  OAI21XL U26944 ( .A0(n22585), .A1(n22582), .B0(n22583), .Y(n22569) );
  NAND2XL U26945 ( .A(n14056), .B(U2_A_i_d[4]), .Y(n22571) );
  OAI21XL U26946 ( .A0(n22570), .A1(n22577), .B0(n22571), .Y(n14022) );
  AOI21XL U26947 ( .A0(n14023), .A1(n22569), .B0(n14022), .Y(n22549) );
  NAND2XL U26948 ( .A(n14024), .B(U2_A_i_d[5]), .Y(n22564) );
  OAI21XL U26949 ( .A0(n22558), .A1(n22564), .B0(n22559), .Y(n22550) );
  NAND2XL U26950 ( .A(n14025), .B(U2_A_i_d[7]), .Y(n22552) );
  INVXL U26951 ( .A(n22552), .Y(n14026) );
  AOI21XL U26952 ( .A0(n22550), .A1(n14015), .B0(n14026), .Y(n14027) );
  OAI21XL U26953 ( .A0(n14028), .A1(n22549), .B0(n14027), .Y(n22521) );
  NOR2XL U26954 ( .A(n14071), .B(U2_A_i_d[9]), .Y(n22533) );
  NOR2XL U26955 ( .A(n14030), .B(U2_A_i_d[8]), .Y(n22532) );
  INVXL U26956 ( .A(n22532), .Y(n22546) );
  NAND2XL U26957 ( .A(n14034), .B(n22546), .Y(n22523) );
  NOR2XL U26958 ( .A(n22523), .B(n14037), .Y(n14039) );
  NAND2XL U26959 ( .A(n14030), .B(U2_A_i_d[8]), .Y(n22545) );
  INVXL U26960 ( .A(n22545), .Y(n14033) );
  NAND2XL U26961 ( .A(n14071), .B(U2_A_i_d[9]), .Y(n22540) );
  OAI21XL U26962 ( .A0(n22535), .A1(n22540), .B0(n22536), .Y(n14032) );
  NAND2XL U26963 ( .A(n14074), .B(U2_A_i_d[11]), .Y(n22529) );
  INVXL U26964 ( .A(n22529), .Y(n22524) );
  NAND2XL U26965 ( .A(n14073), .B(U2_A_i_d[12]), .Y(n22525) );
  INVXL U26966 ( .A(n22525), .Y(n14035) );
  OR2X2 U26967 ( .A(n14086), .B(U2_A_i_d[16]), .Y(n22506) );
  NOR2XL U26968 ( .A(n14042), .B(U2_A_i_d[15]), .Y(n22504) );
  INVXL U26969 ( .A(n22504), .Y(n22510) );
  OR2X2 U26970 ( .A(n14040), .B(U2_A_i_d[13]), .Y(n22519) );
  NAND2XL U26971 ( .A(n22515), .B(n22519), .Y(n22500) );
  NOR2X1 U26972 ( .A(n14046), .B(n22500), .Y(n22434) );
  NAND2XL U26973 ( .A(n14040), .B(U2_A_i_d[13]), .Y(n22518) );
  INVXL U26974 ( .A(n22514), .Y(n14041) );
  AOI21X1 U26975 ( .A0(n22515), .A1(n22513), .B0(n14041), .Y(n22501) );
  NAND2XL U26976 ( .A(n14042), .B(U2_A_i_d[15]), .Y(n22509) );
  INVXL U26977 ( .A(n22509), .Y(n14044) );
  NAND2XL U26978 ( .A(n14086), .B(U2_A_i_d[16]), .Y(n22505) );
  INVXL U26979 ( .A(n22505), .Y(n14043) );
  OR2X2 U26980 ( .A(n14048), .B(U2_A_i_d[18]), .Y(n22494) );
  INVXL U26981 ( .A(n22433), .Y(n14052) );
  NAND2XL U26982 ( .A(n14047), .B(U2_A_i_d[17]), .Y(n22497) );
  INVXL U26983 ( .A(n22497), .Y(n14050) );
  NAND2XL U26984 ( .A(n14048), .B(U2_A_i_d[18]), .Y(n22493) );
  INVXL U26985 ( .A(n22493), .Y(n14049) );
  INVXL U26986 ( .A(n22439), .Y(n14051) );
  NOR2XL U26987 ( .A(n14102), .B(U2_A_i_d[19]), .Y(n22432) );
  NAND2XL U26988 ( .A(n14102), .B(U2_A_i_d[19]), .Y(n22488) );
  NAND2XL U26989 ( .A(n14053), .B(U2_A_i_d[20]), .Y(n22435) );
  NOR2XL U26990 ( .A(n14065), .B(U2_A_i_d[5]), .Y(n22846) );
  NOR2X1 U26991 ( .A(n22848), .B(n22846), .Y(n22840) );
  OR2X2 U26992 ( .A(n14067), .B(U2_A_i_d[7]), .Y(n22842) );
  NOR2XL U26993 ( .A(n13359), .B(U2_A_i_d[4]), .Y(n22861) );
  NOR2XL U26994 ( .A(n14062), .B(U2_A_i_d[3]), .Y(n22867) );
  NOR2XL U26995 ( .A(n22861), .B(n22867), .Y(n14064) );
  NOR2XL U26996 ( .A(n24581), .B(U2_A_i_d[0]), .Y(n22880) );
  AND2XL U26997 ( .A(n14057), .B(U2_A_i_d[1]), .Y(n14058) );
  AOI21XL U26998 ( .A0(n14060), .A1(n14059), .B0(n14058), .Y(n22876) );
  NOR2XL U26999 ( .A(n14061), .B(U2_A_i_d[2]), .Y(n22873) );
  OAI21XL U27000 ( .A0(n22876), .A1(n22873), .B0(n22874), .Y(n22860) );
  NAND2XL U27001 ( .A(n14062), .B(U2_A_i_d[3]), .Y(n22868) );
  NAND2XL U27002 ( .A(n13359), .B(U2_A_i_d[4]), .Y(n22862) );
  OAI21XL U27003 ( .A0(n22861), .A1(n22868), .B0(n22862), .Y(n14063) );
  AOI21XL U27004 ( .A0(n14064), .A1(n22860), .B0(n14063), .Y(n22838) );
  AOI21XL U27005 ( .A0(n22839), .A1(n22842), .B0(n14068), .Y(n14069) );
  OAI21XL U27006 ( .A0(n14070), .A1(n22838), .B0(n14069), .Y(n22807) );
  NOR2XL U27007 ( .A(n5877), .B(U2_A_i_d[9]), .Y(n22822) );
  NOR2XL U27008 ( .A(n14075), .B(U2_A_i_d[8]), .Y(n22821) );
  INVXL U27009 ( .A(n22821), .Y(n14072) );
  NAND2XL U27010 ( .A(n14081), .B(n14072), .Y(n22809) );
  OR2X2 U27011 ( .A(n5876), .B(U2_A_i_d[11]), .Y(n22811) );
  NAND2XL U27012 ( .A(n14075), .B(U2_A_i_d[8]), .Y(n22820) );
  INVXL U27013 ( .A(n22820), .Y(n14080) );
  NAND2XL U27014 ( .A(n5877), .B(U2_A_i_d[9]), .Y(n22823) );
  NAND2XL U27015 ( .A(n14076), .B(U2_A_i_d[10]), .Y(n14077) );
  OAI21XL U27016 ( .A0(n14078), .A1(n22823), .B0(n14077), .Y(n14079) );
  AND2X2 U27017 ( .A(n5876), .B(U2_A_i_d[11]), .Y(n22810) );
  NOR2XL U27018 ( .A(n14091), .B(U2_A_i_d[15]), .Y(n22788) );
  INVXL U27019 ( .A(n22788), .Y(n14087) );
  NAND2XL U27020 ( .A(n14094), .B(n14087), .Y(n14096) );
  OR2X2 U27021 ( .A(n14088), .B(U2_A_i_d[13]), .Y(n22798) );
  NAND2XL U27022 ( .A(n14090), .B(n22798), .Y(n22783) );
  NOR2XL U27023 ( .A(n14096), .B(n22783), .Y(n14132) );
  AND2X2 U27024 ( .A(n14088), .B(U2_A_i_d[13]), .Y(n22797) );
  NAND2XL U27025 ( .A(n14091), .B(U2_A_i_d[15]), .Y(n22787) );
  INVXL U27026 ( .A(n22787), .Y(n14093) );
  AND2X2 U27027 ( .A(n13452), .B(U2_A_i_d[16]), .Y(n14092) );
  AOI21XL U27028 ( .A0(n14094), .A1(n14093), .B0(n14092), .Y(n14095) );
  OAI21XL U27029 ( .A0(n14096), .A1(n22784), .B0(n14095), .Y(n14141) );
  AND2X2 U27030 ( .A(n14099), .B(U2_A_i_d[17]), .Y(n22774) );
  OR2X2 U27031 ( .A(n14103), .B(U2_A_i_d[19]), .Y(n14130) );
  AND2X2 U27032 ( .A(n14103), .B(U2_A_i_d[19]), .Y(n14135) );
  MXI2X1 U27033 ( .A(U1_pipe15[26]), .B(n14110), .S0(n5812), .Y(n4805) );
  NOR2X1 U27034 ( .A(n14120), .B(n14112), .Y(n14123) );
  INVXL U27035 ( .A(n22616), .Y(n14116) );
  INVXL U27036 ( .A(n14114), .Y(n14115) );
  OAI21XL U27037 ( .A0(n14120), .A1(n14119), .B0(n14118), .Y(n14121) );
  NOR2XL U27038 ( .A(n24679), .B(n22957), .Y(n22608) );
  INVXL U27039 ( .A(n22608), .Y(n22613) );
  NAND2XL U27040 ( .A(n22613), .B(n14124), .Y(n22601) );
  INVXL U27041 ( .A(n22612), .Y(n14126) );
  NAND2XL U27042 ( .A(n22958), .B(n24680), .Y(n22609) );
  INVXL U27043 ( .A(n22609), .Y(n14125) );
  NAND2XL U27044 ( .A(n22959), .B(n24684), .Y(n22603) );
  NAND2X1 U27045 ( .A(n22960), .B(n24687), .Y(n22596) );
  OR2X2 U27046 ( .A(n22968), .B(n24693), .Y(n22594) );
  NAND2XL U27047 ( .A(n22968), .B(n24693), .Y(n22593) );
  INVXL U27048 ( .A(n22593), .Y(n14128) );
  NAND2X1 U27049 ( .A(n14136), .B(n14130), .Y(n14138) );
  AND2X2 U27050 ( .A(n14133), .B(U2_A_i_d[20]), .Y(n14134) );
  AOI21X1 U27051 ( .A0(n14136), .A1(n14135), .B0(n14134), .Y(n14137) );
  OAI21X1 U27052 ( .A0(n14144), .A1(n14143), .B0(n14142), .Y(n22744) );
  NOR2XL U27053 ( .A(n14146), .B(U2_A_i_d[21]), .Y(n22760) );
  INVX1 U27054 ( .A(n22449), .Y(n14147) );
  NOR2X1 U27055 ( .A(n14147), .B(U2_A_i_d[22]), .Y(n14149) );
  NOR2XL U27056 ( .A(n22760), .B(n14149), .Y(n22751) );
  NOR2XL U27057 ( .A(n14150), .B(U2_A_i_d[23]), .Y(n14145) );
  INVXL U27058 ( .A(n14145), .Y(n14152) );
  NAND2XL U27059 ( .A(n22751), .B(n14152), .Y(n22746) );
  NOR2XL U27060 ( .A(n14153), .B(U2_A_i_d[24]), .Y(n14155) );
  NOR2XL U27061 ( .A(n22746), .B(n14155), .Y(n14157) );
  NAND2XL U27062 ( .A(n14147), .B(U2_A_i_d[22]), .Y(n14148) );
  OAI21XL U27063 ( .A0(n22759), .A1(n14149), .B0(n14148), .Y(n22752) );
  AND2X1 U27064 ( .A(n14150), .B(U2_A_i_d[23]), .Y(n14151) );
  AOI21X1 U27065 ( .A0(n22752), .A1(n14152), .B0(n14151), .Y(n22745) );
  NAND2XL U27066 ( .A(n14153), .B(U2_A_i_d[24]), .Y(n14154) );
  NOR2XL U27067 ( .A(n14158), .B(U2_A_i_d[25]), .Y(n22738) );
  NAND2XL U27068 ( .A(n14158), .B(U2_A_i_d[25]), .Y(n22739) );
  OAI21X1 U27069 ( .A0(n22742), .A1(n22738), .B0(n22739), .Y(n22735) );
  MXI2X1 U27070 ( .A(U0_pipe10[26]), .B(n14159), .S0(n5812), .Y(n4551) );
  INVXL U27071 ( .A(U0_U0_y2[13]), .Y(n14170) );
  INVXL U27072 ( .A(n14160), .Y(n14172) );
  NAND2XL U27073 ( .A(n14172), .B(n14161), .Y(n14312) );
  OR2X2 U27074 ( .A(U0_U0_y2[9]), .B(U0_U0_y0[9]), .Y(n14175) );
  OR2X2 U27075 ( .A(U0_U0_y2[11]), .B(U0_U0_y0[11]), .Y(n14167) );
  OAI21XL U27076 ( .A0(n14169), .A1(n14177), .B0(n14168), .Y(n14308) );
  AOI21XL U27077 ( .A0(n14172), .A1(n14171), .B0(n8049), .Y(n14313) );
  NAND2XL U27078 ( .A(n14173), .B(U0_U0_y2[13]), .Y(n14318) );
  OAI21XL U27079 ( .A0(n14313), .A1(n14317), .B0(n14318), .Y(n14174) );
  AOI21XL U27080 ( .A0(n14179), .A1(n14308), .B0(n14174), .Y(n14208) );
  NAND2XL U27081 ( .A(n14179), .B(n14309), .Y(n14206) );
  AND2XL U27082 ( .A(U0_U0_y2[0]), .B(U0_U0_y0[0]), .Y(n14181) );
  OR2X2 U27083 ( .A(U0_U0_y2[3]), .B(U0_U0_y0[3]), .Y(n14186) );
  AOI21XL U27084 ( .A0(n14186), .A1(n14185), .B0(n14184), .Y(n14187) );
  OAI21XL U27085 ( .A0(n14189), .A1(n14188), .B0(n14187), .Y(n14205) );
  OR2X2 U27086 ( .A(U0_U0_y2[4]), .B(U0_U0_y0[4]), .Y(n14190) );
  OR2X2 U27087 ( .A(U0_U0_y2[5]), .B(U0_U0_y0[5]), .Y(n14196) );
  OR2X2 U27088 ( .A(U0_U0_y2[7]), .B(U0_U0_y0[7]), .Y(n14199) );
  OAI21XL U27089 ( .A0(n14202), .A1(n14201), .B0(n14200), .Y(n14203) );
  AOI21XL U27090 ( .A0(n14205), .A1(n14204), .B0(n14203), .Y(n14307) );
  OR2X2 U27091 ( .A(n14206), .B(n14307), .Y(n14207) );
  AND2X4 U27092 ( .A(n14208), .B(n14207), .Y(n14330) );
  NOR2XL U27093 ( .A(n14329), .B(n14331), .Y(n14292) );
  NAND2X1 U27094 ( .A(n14292), .B(n14217), .Y(n14276) );
  CMPR22X1 U27095 ( .A(U0_U0_y2[18]), .B(U0_U0_y0[18]), .CO(n14219), .S(n14215) );
  NOR2X2 U27096 ( .A(n14221), .B(n14220), .Y(n14277) );
  ADDHX2 U27097 ( .A(U0_U0_y0[20]), .B(U0_U0_y2[20]), .CO(n14223), .S(n14220)
         );
  NAND2XL U27098 ( .A(n14212), .B(n14211), .Y(n14332) );
  NAND2X2 U27099 ( .A(n14223), .B(n14222), .Y(n14358) );
  ADDHX2 U27100 ( .A(U0_U0_y2[22]), .B(U0_U0_y0[22]), .CO(n14228), .S(n14224)
         );
  CMPR22X1 U27101 ( .A(U0_U0_y2[23]), .B(U0_U0_y0[23]), .CO(n14230), .S(n14227) );
  NOR2X1 U27102 ( .A(n14349), .B(n14351), .Y(n14368) );
  NOR2X2 U27103 ( .A(n14232), .B(n14231), .Y(n14375) );
  NOR2X2 U27104 ( .A(n14234), .B(n14233), .Y(n14370) );
  NOR2X2 U27105 ( .A(n14375), .B(n14370), .Y(n14236) );
  NAND2X1 U27106 ( .A(n14368), .B(n14236), .Y(n14394) );
  CMPR22X1 U27107 ( .A(U0_U0_y2[26]), .B(U0_U0_y0[26]), .CO(n14238), .S(n14233) );
  NOR2X1 U27108 ( .A(n14238), .B(n14237), .Y(n14416) );
  NOR2X1 U27109 ( .A(n14416), .B(n14410), .Y(n14396) );
  NOR2X2 U27110 ( .A(n14242), .B(n14241), .Y(n14403) );
  ADDHX2 U27111 ( .A(U0_U0_y2[29]), .B(U0_U0_y0[29]), .CO(n14244), .S(n14241)
         );
  NOR2X4 U27112 ( .A(n14403), .B(n14397), .Y(n14246) );
  ADDHX2 U27113 ( .A(U0_U0_y2[30]), .B(U0_U0_y0[30]), .CO(n14249), .S(n14243)
         );
  ADDHX2 U27114 ( .A(U0_U0_y2[33]), .B(U0_U0_y0[33]), .CO(n14255), .S(n14252)
         );
  NAND2X1 U27115 ( .A(n14228), .B(n14227), .Y(n14355) );
  NAND2X2 U27116 ( .A(n14232), .B(n14231), .Y(n14376) );
  NAND2XL U27117 ( .A(n14234), .B(n14233), .Y(n14371) );
  OAI21X1 U27118 ( .A0(n14370), .A1(n14376), .B0(n14371), .Y(n14235) );
  AOI21X2 U27119 ( .A0(n14367), .A1(n14236), .B0(n14235), .Y(n14393) );
  NAND2X1 U27120 ( .A(n14238), .B(n14237), .Y(n14417) );
  OAI21X1 U27121 ( .A0(n14397), .A1(n14404), .B0(n14398), .Y(n14245) );
  AOI21X2 U27122 ( .A0(n14246), .A1(n14395), .B0(n14245), .Y(n14247) );
  NAND2X1 U27123 ( .A(n14253), .B(n14252), .Y(n14430) );
  CMPR22X1 U27124 ( .A(U0_U0_y2[37]), .B(U0_U0_y0[37]), .CO(n14268), .S(n14264) );
  CMPR22X1 U27125 ( .A(U0_U0_y2[38]), .B(U0_U0_y0[38]), .CO(n14271), .S(n14267) );
  INVXL U27126 ( .A(n14277), .Y(n14279) );
  NOR2XL U27127 ( .A(n21748), .B(U2_A_r_d[6]), .Y(n14344) );
  INVXL U27128 ( .A(n14282), .Y(n14284) );
  NAND2XL U27129 ( .A(n14284), .B(n14283), .Y(n14285) );
  XOR2X1 U27130 ( .A(n14286), .B(n14285), .Y(n25256) );
  NOR2XL U27131 ( .A(n21747), .B(U2_A_r_d[5]), .Y(n25247) );
  AOI21XL U27132 ( .A0(n14289), .A1(n14288), .B0(n14287), .Y(n14360) );
  NAND2XL U27133 ( .A(n14290), .B(n14358), .Y(n14291) );
  XOR2X1 U27134 ( .A(n14360), .B(n14291), .Y(n25243) );
  OR2X2 U27135 ( .A(n21751), .B(U2_A_r_d[7]), .Y(n14346) );
  NAND2XL U27136 ( .A(n25241), .B(n14346), .Y(n14348) );
  INVXL U27137 ( .A(n14292), .Y(n14295) );
  INVXL U27138 ( .A(n14293), .Y(n14294) );
  OAI21XL U27139 ( .A0(n14330), .A1(n14295), .B0(n14294), .Y(n14306) );
  INVXL U27140 ( .A(n14296), .Y(n14304) );
  INVXL U27141 ( .A(n14303), .Y(n14297) );
  AOI21XL U27142 ( .A0(n14306), .A1(n14304), .B0(n14297), .Y(n14302) );
  INVXL U27143 ( .A(n14298), .Y(n14300) );
  NOR2XL U27144 ( .A(n14338), .B(U2_A_r_d[4]), .Y(n14340) );
  NAND2XL U27145 ( .A(n14304), .B(n14303), .Y(n14305) );
  XNOR2X1 U27146 ( .A(n14306), .B(n14305), .Y(n25269) );
  NOR2XL U27147 ( .A(n21742), .B(U2_A_r_d[3]), .Y(n25262) );
  NOR2XL U27148 ( .A(n14340), .B(n25262), .Y(n14342) );
  INVXL U27149 ( .A(n14307), .Y(n14310) );
  AOI21XL U27150 ( .A0(n14310), .A1(n14309), .B0(n14308), .Y(n14311) );
  INVXL U27151 ( .A(n14311), .Y(n14316) );
  AOI21XL U27152 ( .A0(n14316), .A1(n14315), .B0(n14314), .Y(n14321) );
  INVXL U27153 ( .A(n14317), .Y(n14319) );
  NOR2XL U27154 ( .A(n25285), .B(U2_A_r_d[0]), .Y(n25282) );
  INVXL U27155 ( .A(n25282), .Y(n14327) );
  NOR2XL U27156 ( .A(n21735), .B(U2_A_r_d[1]), .Y(n14324) );
  INVXL U27157 ( .A(n14324), .Y(n14326) );
  AOI21XL U27158 ( .A0(n14327), .A1(n14326), .B0(n14325), .Y(n25277) );
  OAI21XL U27159 ( .A0(n14330), .A1(n14329), .B0(n14328), .Y(n14335) );
  INVXL U27160 ( .A(n14331), .Y(n14333) );
  NOR2XL U27161 ( .A(n21739), .B(U2_A_r_d[2]), .Y(n14337) );
  OAI21XL U27162 ( .A0(n25277), .A1(n14337), .B0(n14336), .Y(n25260) );
  NAND2XL U27163 ( .A(n21742), .B(U2_A_r_d[3]), .Y(n25261) );
  NAND2XL U27164 ( .A(n14338), .B(U2_A_r_d[4]), .Y(n14339) );
  OAI21XL U27165 ( .A0(n14340), .A1(n25261), .B0(n14339), .Y(n14341) );
  AOI21XL U27166 ( .A0(n14342), .A1(n25260), .B0(n14341), .Y(n25239) );
  NAND2XL U27167 ( .A(n21747), .B(U2_A_r_d[5]), .Y(n25248) );
  NAND2XL U27168 ( .A(n21748), .B(U2_A_r_d[6]), .Y(n14343) );
  OAI21XL U27169 ( .A0(n14344), .A1(n25248), .B0(n14343), .Y(n25240) );
  INVXL U27170 ( .A(n14351), .Y(n14353) );
  NOR2XL U27171 ( .A(n5871), .B(U2_A_r_d[10]), .Y(n14382) );
  XNOR2X1 U27172 ( .A(n14369), .B(n14357), .Y(n25231) );
  NOR2XL U27173 ( .A(n14380), .B(U2_A_r_d[9]), .Y(n25222) );
  NOR2XL U27174 ( .A(n21758), .B(U2_A_r_d[8]), .Y(n25221) );
  INVXL U27175 ( .A(n25221), .Y(n14366) );
  NAND2XL U27176 ( .A(n14385), .B(n14366), .Y(n25209) );
  INVXL U27177 ( .A(n14370), .Y(n14372) );
  INVX1 U27178 ( .A(n25212), .Y(n21764) );
  NOR2XL U27179 ( .A(n21764), .B(U2_A_r_d[12]), .Y(n14374) );
  INVXL U27180 ( .A(n14374), .Y(n14388) );
  INVXL U27181 ( .A(n14375), .Y(n14377) );
  NAND2XL U27182 ( .A(n14377), .B(n14376), .Y(n14378) );
  INVXL U27183 ( .A(n25216), .Y(n14386) );
  OR2XL U27184 ( .A(n14386), .B(U2_A_r_d[11]), .Y(n25211) );
  NAND2XL U27185 ( .A(n14388), .B(n25211), .Y(n14390) );
  NOR2XL U27186 ( .A(n25209), .B(n14390), .Y(n14392) );
  NAND2XL U27187 ( .A(n21758), .B(U2_A_r_d[8]), .Y(n25220) );
  INVXL U27188 ( .A(n25220), .Y(n14384) );
  NAND2XL U27189 ( .A(n14380), .B(U2_A_r_d[9]), .Y(n25223) );
  NAND2XL U27190 ( .A(n5871), .B(U2_A_r_d[10]), .Y(n14381) );
  OAI21XL U27191 ( .A0(n14382), .A1(n25223), .B0(n14381), .Y(n14383) );
  AOI21XL U27192 ( .A0(n14388), .A1(n25210), .B0(n14387), .Y(n14389) );
  OAI21X2 U27193 ( .A0(n14421), .A1(n14394), .B0(n14393), .Y(n14409) );
  INVX1 U27194 ( .A(n14397), .Y(n14399) );
  NAND2XL U27195 ( .A(n14399), .B(n14398), .Y(n14400) );
  XNOR2X2 U27196 ( .A(n14401), .B(n14400), .Y(n25189) );
  NOR2XL U27197 ( .A(n14445), .B(U2_A_r_d[16]), .Y(n14402) );
  INVXL U27198 ( .A(n14402), .Y(n14448) );
  NAND2XL U27199 ( .A(n14405), .B(n14404), .Y(n14406) );
  NOR2XL U27200 ( .A(n14444), .B(U2_A_r_d[15]), .Y(n25187) );
  INVXL U27201 ( .A(n25187), .Y(n14408) );
  NAND2XL U27202 ( .A(n14448), .B(n14408), .Y(n14450) );
  INVXL U27203 ( .A(n14410), .Y(n14412) );
  XNOR2X2 U27204 ( .A(n14414), .B(n14413), .Y(n25199) );
  NOR2XL U27205 ( .A(n21774), .B(U2_A_r_d[14]), .Y(n14415) );
  INVXL U27206 ( .A(n14415), .Y(n14443) );
  INVXL U27207 ( .A(n14416), .Y(n14418) );
  NAND2XL U27208 ( .A(n14418), .B(n14417), .Y(n14419) );
  INVXL U27209 ( .A(n25203), .Y(n14441) );
  OR2X2 U27210 ( .A(n14441), .B(U2_A_r_d[13]), .Y(n25198) );
  NAND2XL U27211 ( .A(n14443), .B(n25198), .Y(n25182) );
  NOR2XL U27212 ( .A(n14450), .B(n25182), .Y(n25157) );
  INVXL U27213 ( .A(n14425), .Y(n14427) );
  NAND2X1 U27214 ( .A(n14431), .B(n14430), .Y(n14432) );
  INVX1 U27215 ( .A(n25166), .Y(n14453) );
  OR2X2 U27216 ( .A(n14453), .B(U2_A_r_d[19]), .Y(n25161) );
  NAND2X1 U27217 ( .A(n14455), .B(n25161), .Y(n14457) );
  OR2X2 U27218 ( .A(n21781), .B(U2_A_r_d[18]), .Y(n14452) );
  XOR2X2 U27219 ( .A(n14464), .B(n14440), .Y(n25178) );
  OR2X2 U27220 ( .A(n5863), .B(U2_A_r_d[17]), .Y(n25172) );
  NAND2XL U27221 ( .A(n14452), .B(n25172), .Y(n25159) );
  NOR2XL U27222 ( .A(n14457), .B(n25159), .Y(n14459) );
  NAND2XL U27223 ( .A(n25157), .B(n14459), .Y(n14461) );
  AOI21XL U27224 ( .A0(n14443), .A1(n25197), .B0(n14442), .Y(n25183) );
  NAND2XL U27225 ( .A(n14444), .B(U2_A_r_d[15]), .Y(n25186) );
  INVXL U27226 ( .A(n25186), .Y(n14447) );
  AOI21XL U27227 ( .A0(n14448), .A1(n14447), .B0(n14446), .Y(n14449) );
  OAI21XL U27228 ( .A0(n14450), .A1(n25183), .B0(n14449), .Y(n25156) );
  AND2X2 U27229 ( .A(n5863), .B(U2_A_r_d[17]), .Y(n25171) );
  AND2X2 U27230 ( .A(n21781), .B(U2_A_r_d[18]), .Y(n14451) );
  AOI21X1 U27231 ( .A0(n14452), .A1(n25171), .B0(n14451), .Y(n25158) );
  OAI21XL U27232 ( .A0(n14457), .A1(n25158), .B0(n14456), .Y(n14458) );
  AOI21X1 U27233 ( .A0(n25156), .A1(n14459), .B0(n14458), .Y(n14460) );
  OAI21X1 U27234 ( .A0(n25155), .A1(n14461), .B0(n14460), .Y(n25129) );
  XNOR2X2 U27235 ( .A(n14469), .B(n14468), .Y(n25151) );
  NOR2XL U27236 ( .A(n21794), .B(U2_A_r_d[21]), .Y(n25146) );
  NAND2XL U27237 ( .A(n14260), .B(n14470), .Y(n14471) );
  NOR2XL U27238 ( .A(n14482), .B(U2_A_r_d[22]), .Y(n14483) );
  NOR2XL U27239 ( .A(n25146), .B(n14483), .Y(n25137) );
  NOR2XL U27240 ( .A(n14484), .B(U2_A_r_d[23]), .Y(n14478) );
  INVXL U27241 ( .A(n14478), .Y(n14486) );
  NAND2XL U27242 ( .A(n25137), .B(n14486), .Y(n25131) );
  XNOR2X2 U27243 ( .A(n14481), .B(n14480), .Y(n25132) );
  INVX1 U27244 ( .A(n25132), .Y(n21800) );
  NOR2XL U27245 ( .A(n21800), .B(U2_A_r_d[24]), .Y(n14488) );
  NOR2XL U27246 ( .A(n25131), .B(n14488), .Y(n14490) );
  NAND2XL U27247 ( .A(n21794), .B(U2_A_r_d[21]), .Y(n25145) );
  NAND2XL U27248 ( .A(n21800), .B(U2_A_r_d[24]), .Y(n14487) );
  OAI21XL U27249 ( .A0(n25130), .A1(n14488), .B0(n14487), .Y(n14489) );
  NOR2XL U27250 ( .A(n21805), .B(U2_A_r_d[25]), .Y(n14497) );
  NAND2XL U27251 ( .A(n21805), .B(U2_A_r_d[25]), .Y(n14496) );
  OAI21X1 U27252 ( .A0(n25127), .A1(n14497), .B0(n14496), .Y(n25122) );
  INVXL U27253 ( .A(n14962), .Y(n14507) );
  NOR2XL U27254 ( .A(n19557), .B(n14507), .Y(n17621) );
  NAND2XL U27255 ( .A(n5861), .B(n19248), .Y(n14508) );
  NAND2XL U27256 ( .A(n14510), .B(n19237), .Y(n14511) );
  NOR2XL U27257 ( .A(n14525), .B(n22886), .Y(n22065) );
  NOR2XL U27258 ( .A(n22067), .B(n22065), .Y(n22060) );
  NAND2XL U27259 ( .A(n22060), .B(n14514), .Y(n14529) );
  NOR2XL U27260 ( .A(n14522), .B(n22889), .Y(n22081) );
  NOR2XL U27261 ( .A(n22081), .B(n22080), .Y(n14524) );
  NOR2XL U27262 ( .A(n25449), .B(n22727), .Y(n22098) );
  AOI21XL U27263 ( .A0(n14517), .A1(n5767), .B0(n14516), .Y(n22094) );
  OAI21XL U27264 ( .A0(n22094), .A1(n14520), .B0(n14519), .Y(n22078) );
  NAND2XL U27265 ( .A(n14521), .B(n22890), .Y(n22079) );
  NAND2XL U27266 ( .A(n14522), .B(n22889), .Y(n22082) );
  AOI21XL U27267 ( .A0(n14524), .A1(n22078), .B0(n14523), .Y(n22058) );
  NAND2XL U27268 ( .A(n14526), .B(n22885), .Y(n22068) );
  NOR2X1 U27269 ( .A(n14536), .B(n22913), .Y(n14538) );
  NOR2XL U27270 ( .A(n14535), .B(n22914), .Y(n22040) );
  NOR2XL U27271 ( .A(n14534), .B(n22915), .Y(n22039) );
  INVXL U27272 ( .A(n22039), .Y(n14531) );
  NOR2X1 U27273 ( .A(n22026), .B(n14544), .Y(n14546) );
  NAND2XL U27274 ( .A(n14534), .B(n22915), .Y(n22038) );
  INVXL U27275 ( .A(n22038), .Y(n14540) );
  NAND2XL U27276 ( .A(n14535), .B(n22914), .Y(n22041) );
  NAND2XL U27277 ( .A(n14536), .B(n22913), .Y(n14537) );
  OAI21XL U27278 ( .A0(n14538), .A1(n22041), .B0(n14537), .Y(n14539) );
  OR2X2 U27279 ( .A(n14553), .B(n22935), .Y(n22016) );
  NAND2XL U27280 ( .A(n22016), .B(n14549), .Y(n22000) );
  OR2X2 U27281 ( .A(n14564), .B(n22930), .Y(n14566) );
  NOR2XL U27282 ( .A(n5852), .B(n22931), .Y(n14551) );
  INVXL U27283 ( .A(n14551), .Y(n21983) );
  NAND2X1 U27284 ( .A(n14566), .B(n21983), .Y(n14568) );
  OR2X2 U27285 ( .A(n14562), .B(n22932), .Y(n14563) );
  NAND2X1 U27286 ( .A(n14563), .B(n14552), .Y(n21981) );
  NOR2X1 U27287 ( .A(n14568), .B(n21981), .Y(n14569) );
  NAND2XL U27288 ( .A(n12388), .B(n22936), .Y(n22020) );
  INVXL U27289 ( .A(n22020), .Y(n22014) );
  NAND2XL U27290 ( .A(n14553), .B(n22935), .Y(n22015) );
  INVXL U27291 ( .A(n22015), .Y(n14554) );
  AOI21X1 U27292 ( .A0(n22016), .A1(n22014), .B0(n14554), .Y(n22001) );
  NAND2XL U27293 ( .A(n5864), .B(n22934), .Y(n22009) );
  INVXL U27294 ( .A(n22009), .Y(n14557) );
  INVXL U27295 ( .A(n22005), .Y(n14556) );
  AOI21X1 U27296 ( .A0(n14563), .A1(n14561), .B0(n8105), .Y(n21980) );
  AND2X2 U27297 ( .A(n5852), .B(n22931), .Y(n21982) );
  AOI21XL U27298 ( .A0(n14566), .A1(n21982), .B0(n14565), .Y(n14567) );
  NOR2XL U27299 ( .A(n14571), .B(n22957), .Y(n21968) );
  NOR2XL U27300 ( .A(n21968), .B(n14574), .Y(n21957) );
  INVX1 U27301 ( .A(n14570), .Y(n14575) );
  NAND2XL U27302 ( .A(n21957), .B(n14576), .Y(n21954) );
  NAND2XL U27303 ( .A(n14571), .B(n22957), .Y(n21967) );
  NAND2XL U27304 ( .A(n14572), .B(n22958), .Y(n14573) );
  OAI21XL U27305 ( .A0(n21967), .A1(n14574), .B0(n14573), .Y(n21958) );
  NAND2XL U27306 ( .A(n14577), .B(n22960), .Y(n14578) );
  MXI2X1 U27307 ( .A(U0_pipe7[27]), .B(n14583), .S0(n5812), .Y(n4435) );
  CMPR22X1 U27308 ( .A(U1_U1_y1[16]), .B(U1_U1_y0[16]), .CO(n14639), .S(n14636) );
  CMPR22X1 U27309 ( .A(U1_U1_y1[17]), .B(U1_U1_y0[17]), .CO(n14641), .S(n14638) );
  OR2XL U27310 ( .A(U1_U1_y1[1]), .B(U1_U1_y0[1]), .Y(n14586) );
  AND2XL U27311 ( .A(U1_U1_y1[0]), .B(U1_U1_y0[0]), .Y(n14585) );
  AOI21XL U27312 ( .A0(n14586), .A1(n14585), .B0(n14584), .Y(n14595) );
  NAND2XL U27313 ( .A(n14589), .B(n14592), .Y(n14594) );
  OAI21XL U27314 ( .A0(n14595), .A1(n14594), .B0(n14593), .Y(n14612) );
  OR2X2 U27315 ( .A(U1_U1_y1[7]), .B(U1_U1_y0[7]), .Y(n14606) );
  OAI21XL U27316 ( .A0(n14609), .A1(n14608), .B0(n14607), .Y(n14610) );
  AOI21XL U27317 ( .A0(n14612), .A1(n14611), .B0(n14610), .Y(n14716) );
  INVXL U27318 ( .A(U1_U1_y1[13]), .Y(n14627) );
  OR2X2 U27319 ( .A(n14627), .B(U1_U1_y0[13]), .Y(n14630) );
  OR2X2 U27320 ( .A(U1_U1_y1[12]), .B(U1_U1_y0[12]), .Y(n14613) );
  NAND2XL U27321 ( .A(n14630), .B(n14613), .Y(n14721) );
  CMPR22X1 U27322 ( .A(U1_U1_y1[14]), .B(U1_U1_y0[14]), .CO(n14635), .S(n14631) );
  OR2X2 U27323 ( .A(U1_U1_y1[9]), .B(U1_U1_y0[9]), .Y(n14620) );
  OR2X2 U27324 ( .A(U1_U1_y1[11]), .B(U1_U1_y0[11]), .Y(n14623) );
  NAND2XL U27325 ( .A(n14616), .B(n14623), .Y(n14625) );
  AOI21XL U27326 ( .A0(n14620), .A1(n14619), .B0(n14618), .Y(n14626) );
  AOI21XL U27327 ( .A0(n14623), .A1(n14622), .B0(n14621), .Y(n14624) );
  OAI21XL U27328 ( .A0(n14626), .A1(n14625), .B0(n14624), .Y(n14717) );
  AOI21XL U27329 ( .A0(n14630), .A1(n14629), .B0(n14628), .Y(n14722) );
  NAND2XL U27330 ( .A(n14631), .B(U1_U1_y1[13]), .Y(n14727) );
  OAI21XL U27331 ( .A0(n14722), .A1(n14726), .B0(n14727), .Y(n14632) );
  CMPR22X1 U27332 ( .A(U1_U1_y1[33]), .B(U1_U1_y0[33]), .CO(n14673), .S(n14670) );
  CMPR22X1 U27333 ( .A(U1_U1_y1[34]), .B(U1_U1_y0[34]), .CO(n14676), .S(n14672) );
  OR2X2 U27334 ( .A(n14678), .B(n14677), .Y(n14845) );
  NOR2X1 U27335 ( .A(n14680), .B(n14679), .Y(n14846) );
  CMPR22X1 U27336 ( .A(U1_U1_y1[37]), .B(U1_U1_y0[37]), .CO(n14683), .S(n14679) );
  CMPR22X1 U27337 ( .A(U1_U1_y1[38]), .B(U1_U1_y0[38]), .CO(n14686), .S(n14682) );
  INVXL U27338 ( .A(n14702), .Y(n14700) );
  OAI21XL U27339 ( .A0(n14700), .A1(n14696), .B0(n14697), .Y(n14695) );
  INVXL U27340 ( .A(n14692), .Y(n14694) );
  NAND2XL U27341 ( .A(n14698), .B(n14697), .Y(n14699) );
  INVXL U27342 ( .A(n19965), .Y(n14754) );
  INVXL U27343 ( .A(n14767), .Y(n14704) );
  INVXL U27344 ( .A(n19969), .Y(n14755) );
  INVXL U27345 ( .A(n14706), .Y(n14709) );
  INVXL U27346 ( .A(n14707), .Y(n14708) );
  AOI21XL U27347 ( .A0(n14715), .A1(n7034), .B0(n7359), .Y(n14712) );
  INVXL U27348 ( .A(n19962), .Y(n14749) );
  NOR2XL U27349 ( .A(n14749), .B(n19358), .Y(n14751) );
  NAND2XL U27350 ( .A(n7034), .B(n14713), .Y(n14714) );
  INVXL U27351 ( .A(n19960), .Y(n14748) );
  NOR2XL U27352 ( .A(n14748), .B(n19363), .Y(n19357) );
  NOR2XL U27353 ( .A(n14751), .B(n19357), .Y(n14753) );
  INVXL U27354 ( .A(n14721), .Y(n14724) );
  INVXL U27355 ( .A(n14722), .Y(n14723) );
  INVXL U27356 ( .A(n14726), .Y(n14728) );
  INVXL U27357 ( .A(n14739), .Y(n14731) );
  NAND2XL U27358 ( .A(n14731), .B(n14738), .Y(n14732) );
  INVXL U27359 ( .A(n19954), .Y(n14734) );
  NOR2XL U27360 ( .A(n14734), .B(n19373), .Y(n14733) );
  INVXL U27361 ( .A(n14733), .Y(n14736) );
  AOI21XL U27362 ( .A0(n14737), .A1(n14736), .B0(n14735), .Y(n19370) );
  OAI21XL U27363 ( .A0(n14740), .A1(n14739), .B0(n14738), .Y(n14744) );
  INVXL U27364 ( .A(n19956), .Y(n14745) );
  NOR2XL U27365 ( .A(n14745), .B(n19369), .Y(n14747) );
  OAI21XL U27366 ( .A0(n19370), .A1(n14747), .B0(n14746), .Y(n19355) );
  NAND2XL U27367 ( .A(n14748), .B(n19363), .Y(n19356) );
  NAND2XL U27368 ( .A(n14749), .B(n19358), .Y(n14750) );
  OAI21XL U27369 ( .A0(n14751), .A1(n19356), .B0(n14750), .Y(n14752) );
  AOI21XL U27370 ( .A0(n14753), .A1(n19355), .B0(n14752), .Y(n19334) );
  NAND2XL U27371 ( .A(n14754), .B(n19518), .Y(n19350) );
  AOI21XL U27372 ( .A0(n19335), .A1(n19338), .B0(n14756), .Y(n14757) );
  INVXL U27373 ( .A(n14760), .Y(n14762) );
  NOR2XL U27374 ( .A(n14785), .B(n19321), .Y(n14787) );
  INVXL U27375 ( .A(n19978), .Y(n14784) );
  NOR2XL U27376 ( .A(n14784), .B(n19326), .Y(n19317) );
  NOR2XL U27377 ( .A(n14787), .B(n19317), .Y(n14790) );
  INVXL U27378 ( .A(n19316), .Y(n14773) );
  OR2X2 U27379 ( .A(n14791), .B(n19532), .Y(n19306) );
  NAND2XL U27380 ( .A(n14781), .B(n14780), .Y(n14782) );
  NAND2XL U27381 ( .A(n14783), .B(n19330), .Y(n19315) );
  INVXL U27382 ( .A(n19315), .Y(n14789) );
  NAND2XL U27383 ( .A(n14784), .B(n19326), .Y(n19318) );
  NAND2XL U27384 ( .A(n14785), .B(n19321), .Y(n14786) );
  OAI21XL U27385 ( .A0(n14787), .A1(n19318), .B0(n14786), .Y(n14788) );
  NAND2XL U27386 ( .A(n14791), .B(n19532), .Y(n19305) );
  INVXL U27387 ( .A(n14794), .Y(n14796) );
  OR2X2 U27388 ( .A(n19553), .B(n14835), .Y(n19263) );
  INVXL U27389 ( .A(n14801), .Y(n14803) );
  INVXL U27390 ( .A(n20001), .Y(n14825) );
  NAND2XL U27391 ( .A(n19293), .B(n14824), .Y(n19276) );
  NAND2XL U27392 ( .A(n14825), .B(n19541), .Y(n19297) );
  INVXL U27393 ( .A(n19297), .Y(n19291) );
  INVXL U27394 ( .A(n19292), .Y(n14827) );
  INVXL U27395 ( .A(n19286), .Y(n14829) );
  AOI21XL U27396 ( .A0(n14830), .A1(n14829), .B0(n8144), .Y(n14831) );
  INVXL U27397 ( .A(n20033), .Y(n14856) );
  NAND2XL U27398 ( .A(n14852), .B(n19248), .Y(n14853) );
  NAND2XL U27399 ( .A(n14856), .B(n19237), .Y(n14857) );
  NAND2XL U27400 ( .A(n14863), .B(n19233), .Y(n14864) );
  NOR2XL U27401 ( .A(n19965), .B(n14901), .Y(n20426) );
  NOR2XL U27402 ( .A(n20428), .B(n20426), .Y(n20421) );
  NAND2XL U27403 ( .A(n20421), .B(n14865), .Y(n14872) );
  NOR2XL U27404 ( .A(n19962), .B(n19951), .Y(n20443) );
  NOR2XL U27405 ( .A(n19960), .B(n14904), .Y(n20442) );
  NOR2XL U27406 ( .A(n20443), .B(n20442), .Y(n14869) );
  NAND2XL U27407 ( .A(n19954), .B(n19952), .Y(n20175) );
  INVXL U27408 ( .A(n20175), .Y(n14867) );
  AOI21XL U27409 ( .A0(n20455), .A1(n14866), .B0(n14867), .Y(n20452) );
  NOR2XL U27410 ( .A(n19956), .B(n14911), .Y(n20169) );
  NAND2XL U27411 ( .A(n19956), .B(n14911), .Y(n20170) );
  OAI21XL U27412 ( .A0(n20452), .A1(n20169), .B0(n20170), .Y(n20440) );
  NAND2XL U27413 ( .A(n19960), .B(n14904), .Y(n20441) );
  NAND2XL U27414 ( .A(n19962), .B(n19951), .Y(n20444) );
  AOI21XL U27415 ( .A0(n14869), .A1(n20440), .B0(n14868), .Y(n20419) );
  NAND2XL U27416 ( .A(n19965), .B(n14901), .Y(n20434) );
  NAND2XL U27417 ( .A(n19967), .B(n14900), .Y(n20429) );
  NAND2XL U27418 ( .A(n19969), .B(n14902), .Y(n20422) );
  INVXL U27419 ( .A(n20422), .Y(n14870) );
  NOR2XL U27420 ( .A(n19978), .B(n19974), .Y(n20403) );
  NOR2X1 U27421 ( .A(n20405), .B(n20403), .Y(n14877) );
  NOR2XL U27422 ( .A(n19976), .B(n14927), .Y(n20402) );
  INVXL U27423 ( .A(n20402), .Y(n20132) );
  NAND2XL U27424 ( .A(n14877), .B(n20132), .Y(n20390) );
  INVX1 U27425 ( .A(n14873), .Y(n20393) );
  NAND2X1 U27426 ( .A(n20393), .B(n14874), .Y(n14880) );
  NAND2XL U27427 ( .A(n19976), .B(n14927), .Y(n20401) );
  INVXL U27428 ( .A(n20401), .Y(n14876) );
  NAND2XL U27429 ( .A(n19978), .B(n19974), .Y(n20411) );
  NAND2XL U27430 ( .A(n19979), .B(n14926), .Y(n20406) );
  OAI21XL U27431 ( .A0(n20405), .A1(n20411), .B0(n20406), .Y(n14875) );
  NAND2XL U27432 ( .A(n19984), .B(n14930), .Y(n20397) );
  INVXL U27433 ( .A(n20397), .Y(n20391) );
  NAND2XL U27434 ( .A(n19986), .B(n14929), .Y(n20392) );
  INVXL U27435 ( .A(n20392), .Y(n14878) );
  AOI21X1 U27436 ( .A0(n20393), .A1(n20391), .B0(n14878), .Y(n14879) );
  OAI21X1 U27437 ( .A0(n20389), .A1(n14880), .B0(n14879), .Y(n14881) );
  INVX2 U27438 ( .A(n20320), .Y(n20386) );
  OR2X2 U27439 ( .A(n20001), .B(n14946), .Y(n20384) );
  NAND2XL U27440 ( .A(n20001), .B(n14946), .Y(n20383) );
  NAND2XL U27441 ( .A(n20003), .B(n19994), .Y(n20378) );
  INVXL U27442 ( .A(n20378), .Y(n14883) );
  INVXL U27443 ( .A(n20372), .Y(n14885) );
  NAND2XL U27444 ( .A(n20007), .B(n19993), .Y(n20368) );
  INVXL U27445 ( .A(n20368), .Y(n14884) );
  INVXL U27446 ( .A(n20309), .Y(n14889) );
  NAND2X1 U27447 ( .A(n20013), .B(n19996), .Y(n20311) );
  NAND2XL U27448 ( .A(n20015), .B(n14948), .Y(n20312) );
  INVXL U27449 ( .A(n14893), .Y(n14894) );
  NAND2X1 U27450 ( .A(n14897), .B(n29007), .Y(n19385) );
  NOR2XL U27451 ( .A(n19966), .B(n14921), .Y(n16896) );
  NOR2XL U27452 ( .A(n16898), .B(n16896), .Y(n16891) );
  NAND2XL U27453 ( .A(n16891), .B(n14903), .Y(n14925) );
  NOR2XL U27454 ( .A(n5883), .B(n14916), .Y(n14918) );
  NOR2XL U27455 ( .A(n19961), .B(n14915), .Y(n16911) );
  NOR2XL U27456 ( .A(n14918), .B(n16911), .Y(n14920) );
  INVXL U27457 ( .A(n19952), .Y(n14908) );
  AOI21XL U27458 ( .A0(n14910), .A1(n14906), .B0(n14909), .Y(n16925) );
  NOR2XL U27459 ( .A(n19957), .B(n14912), .Y(n14914) );
  NAND2XL U27460 ( .A(n19957), .B(n14912), .Y(n14913) );
  OAI21XL U27461 ( .A0(n16925), .A1(n14914), .B0(n14913), .Y(n16909) );
  NAND2XL U27462 ( .A(n19961), .B(n14915), .Y(n16910) );
  NAND2XL U27463 ( .A(n5883), .B(n14916), .Y(n14917) );
  OAI21XL U27464 ( .A0(n14918), .A1(n16910), .B0(n14917), .Y(n14919) );
  NAND2XL U27465 ( .A(n19966), .B(n14921), .Y(n16904) );
  NAND2XL U27466 ( .A(n19968), .B(n14922), .Y(n16899) );
  NAND2XL U27467 ( .A(n19970), .B(n14923), .Y(n16892) );
  NOR2XL U27468 ( .A(n19980), .B(n14935), .Y(n14937) );
  NOR2XL U27469 ( .A(n19977), .B(n14932), .Y(n16870) );
  INVXL U27470 ( .A(n16870), .Y(n14928) );
  NOR2XL U27471 ( .A(n19985), .B(n14940), .Y(n14931) );
  INVXL U27472 ( .A(n14931), .Y(n16860) );
  NAND2XL U27473 ( .A(n19977), .B(n14932), .Y(n16869) );
  INVXL U27474 ( .A(n16869), .Y(n14938) );
  NAND2XL U27475 ( .A(n14934), .B(n14933), .Y(n16872) );
  NAND2XL U27476 ( .A(n19980), .B(n14935), .Y(n14936) );
  NAND2XL U27477 ( .A(n16849), .B(n14947), .Y(n16834) );
  OR2X2 U27478 ( .A(n20014), .B(n14959), .Y(n16813) );
  NOR2XL U27479 ( .A(n20020), .B(n14968), .Y(n14970) );
  NAND2XL U27480 ( .A(n20016), .B(n14962), .Y(n16799) );
  NAND2XL U27481 ( .A(n5850), .B(n14963), .Y(n14964) );
  NAND2XL U27482 ( .A(n20020), .B(n14968), .Y(n14969) );
  MXI2X1 U27483 ( .A(U1_pipe7[27]), .B(n14973), .S0(n5812), .Y(n4980) );
  MXI2X1 U27484 ( .A(U1_pipe2[26]), .B(n14975), .S0(n5812), .Y(n5038) );
  OAI222X4 U27485 ( .A0(n14979), .A1(n28674), .B0(n14978), .B1(n28704), .C0(
        n28680), .C1(n14977), .Y(T1_rom_addr[4]) );
  OAI222X4 U27486 ( .A0(n14979), .A1(n28679), .B0(n14978), .B1(n28703), .C0(
        n28673), .C1(n14977), .Y(T1_rom_addr[5]) );
  AOI21XL U27487 ( .A0(Q0_addr[0]), .A1(n5826), .B0(n27081), .Y(n14983) );
  NAND3BX2 U27488 ( .AN(n28322), .B(n14981), .C(n14980), .Y(n27088) );
  OAI211X4 U27489 ( .A0(n28752), .A1(n7140), .B0(n14983), .C0(n14982), .Y(
        A3_addr[0]) );
  AOI21XL U27490 ( .A0(n5826), .A1(Q0_addr[1]), .B0(n27073), .Y(n14985) );
  OAI211X4 U27491 ( .A0(n7140), .A1(n28753), .B0(n14985), .C0(n14984), .Y(
        A3_addr[1]) );
  AOI21XL U27492 ( .A0(n27162), .A1(Q0_addr[2]), .B0(n27084), .Y(n14987) );
  OAI211X4 U27493 ( .A0(n7140), .A1(n28755), .B0(n14987), .C0(n14986), .Y(
        A3_addr[2]) );
  AOI21XL U27494 ( .A0(n5826), .A1(Q0_addr[3]), .B0(n14988), .Y(n14990) );
  OAI211X4 U27495 ( .A0(n7140), .A1(n28756), .B0(n14990), .C0(n14989), .Y(
        A3_addr[3]) );
  OAI32X4 U27496 ( .A0(n7305), .A1(n28677), .A2(n28672), .B0(n14993), .B1(
        n11633), .Y(n16569) );
  OAI21XL U27497 ( .A0(n6885), .A1(BOPA[27]), .B0(n15002), .Y(n3715) );
  AOI21XL U27498 ( .A0(n5826), .A1(Q0_addr[4]), .B0(n27078), .Y(n15005) );
  OAI211X4 U27499 ( .A0(n7140), .A1(n28754), .B0(n15005), .C0(n15004), .Y(
        A3_addr[4]) );
  OAI21XL U27500 ( .A0(n5910), .A1(BOPA[33]), .B0(n15008), .Y(n3743) );
  OAI21XL U27501 ( .A0(n5910), .A1(BOPA[35]), .B0(n15012), .Y(n3751) );
  OAI21XL U27502 ( .A0(n5907), .A1(BOPA[34]), .B0(n15016), .Y(n3747) );
  OAI21XL U27503 ( .A0(n6886), .A1(BOPA[32]), .B0(n15019), .Y(n3739) );
  OAI21XL U27504 ( .A0(n6883), .A1(BOPA[26]), .B0(n15022), .Y(n3711) );
  AOI21XL U27505 ( .A0(n27162), .A1(Q0_addr[5]), .B0(n15028), .Y(n15030) );
  OAI211X4 U27506 ( .A0(n7140), .A1(n28757), .B0(n15030), .C0(n15029), .Y(
        A3_addr[5]) );
  OAI211X4 U27507 ( .A0(n7140), .A1(n28919), .B0(n15033), .C0(n15032), .Y(
        A3_addr[6]) );
  OAI21XL U27508 ( .A0(n6886), .A1(BOPA[28]), .B0(n15037), .Y(n3719) );
  AOI21XL U27509 ( .A0(n5826), .A1(Q0_addr[7]), .B0(n15038), .Y(n15040) );
  OAI211X4 U27510 ( .A0(n7140), .A1(n28920), .B0(n15040), .C0(n15039), .Y(
        A3_addr[7]) );
  NAND2X1 U27511 ( .A(n28672), .B(n28678), .Y(n15129) );
  CLKINVX3 U27512 ( .A(n15129), .Y(n15969) );
  OAI21XL U27513 ( .A0(n5905), .A1(AOPB[51]), .B0(n15044), .Y(n3404) );
  OAI21XL U27514 ( .A0(n5905), .A1(AOPB[50]), .B0(n15048), .Y(n3400) );
  OAI21XL U27515 ( .A0(n5917), .A1(AOPB[49]), .B0(n15051), .Y(n3392) );
  OAI21XL U27516 ( .A0(n5917), .A1(AOPB[48]), .B0(n15055), .Y(n3388) );
  OAI21XL U27517 ( .A0(n16378), .A1(n5836), .B0(n5915), .Y(n15056) );
  OAI2BB2XL U27518 ( .B0(n5915), .B1(AOPB[47]), .A0N(n15058), .A1N(n15057), 
        .Y(n3384) );
  OAI21XL U27519 ( .A0(n5836), .A1(n16382), .B0(n15061), .Y(n15062) );
  OAI21XL U27520 ( .A0(R7_valid), .A1(AOPB[46]), .B0(n15062), .Y(n3380) );
  OAI21XL U27521 ( .A0(n5912), .A1(AOPB[45]), .B0(n15065), .Y(n3376) );
  OAI21XL U27522 ( .A0(n5917), .A1(AOPB[44]), .B0(n15068), .Y(n3372) );
  OAI21XL U27523 ( .A0(n6881), .A1(AOPB[43]), .B0(n15072), .Y(n3368) );
  OAI21XL U27524 ( .A0(n5917), .A1(AOPB[42]), .B0(n15075), .Y(n3364) );
  OAI21XL U27525 ( .A0(n6885), .A1(AOPB[41]), .B0(n15078), .Y(n3360) );
  OAI21XL U27526 ( .A0(n5917), .A1(AOPB[40]), .B0(n15081), .Y(n3356) );
  OAI21XL U27527 ( .A0(n16410), .A1(n5836), .B0(n5800), .Y(n15082) );
  OAI2BB2XL U27528 ( .B0(n5915), .B1(AOPB[39]), .A0N(n15084), .A1N(n15083), 
        .Y(n3348) );
  OAI21XL U27529 ( .A0(n16414), .A1(n15129), .B0(R7_valid), .Y(n15085) );
  OAI2BB2XL U27530 ( .B0(n5909), .B1(AOPB[38]), .A0N(n15087), .A1N(n15086), 
        .Y(n3344) );
  OAI21XL U27531 ( .A0(n16419), .A1(n15129), .B0(n6880), .Y(n15088) );
  OAI2BB2XL U27532 ( .B0(n5915), .B1(AOPB[37]), .A0N(n15090), .A1N(n15089), 
        .Y(n3340) );
  OAI21XL U27533 ( .A0(n6881), .A1(AOPB[36]), .B0(n15094), .Y(n3336) );
  OAI21XL U27534 ( .A0(n16427), .A1(n15129), .B0(n5907), .Y(n15095) );
  OAI2BB2XL U27535 ( .B0(n5909), .B1(AOPB[35]), .A0N(n15097), .A1N(n15096), 
        .Y(n3332) );
  OAI21XL U27536 ( .A0(n5908), .A1(AOPB[34]), .B0(n15100), .Y(n3328) );
  OAI21XL U27537 ( .A0(n6885), .A1(AOPB[33]), .B0(n15103), .Y(n3324) );
  OAI21XL U27538 ( .A0(n5836), .A1(n16439), .B0(n15106), .Y(n15107) );
  OAI21XL U27539 ( .A0(n5917), .A1(AOPB[32]), .B0(n15107), .Y(n3320) );
  OAI21XL U27540 ( .A0(n6881), .A1(AOPB[31]), .B0(n15111), .Y(n3316) );
  OAI21XL U27541 ( .A0(n16447), .A1(n5836), .B0(R7_valid), .Y(n15112) );
  OAI2BB2XL U27542 ( .B0(n5909), .B1(AOPB[30]), .A0N(n15114), .A1N(n15113), 
        .Y(n3312) );
  OAI21XL U27543 ( .A0(n16451), .A1(n15129), .B0(R7_valid), .Y(n15115) );
  OAI2BB2XL U27544 ( .B0(n5915), .B1(AOPB[29]), .A0N(n15117), .A1N(n15116), 
        .Y(n3304) );
  OAI21XL U27545 ( .A0(n5908), .A1(AOPB[28]), .B0(n15120), .Y(n3300) );
  OAI21XL U27546 ( .A0(n5910), .A1(AOPB[27]), .B0(n15124), .Y(n3296) );
  OAI21XL U27547 ( .A0(n6885), .A1(AOPB[26]), .B0(n15128), .Y(n3292) );
  OAI21XL U27548 ( .A0(n16468), .A1(n15129), .B0(n5908), .Y(n15130) );
  OAI21XL U27549 ( .A0(n16473), .A1(n5836), .B0(n5905), .Y(n15133) );
  OAI21XL U27550 ( .A0(n5906), .A1(AOPB[23]), .B0(n15139), .Y(n3280) );
  OAI21XL U27551 ( .A0(n5917), .A1(AOPB[22]), .B0(n15142), .Y(n3276) );
  OAI21XL U27552 ( .A0(R7_valid), .A1(AOPB[21]), .B0(n15146), .Y(n3272) );
  OAI21XL U27553 ( .A0(n5910), .A1(AOPB[20]), .B0(n15150), .Y(n3268) );
  OAI21XL U27554 ( .A0(n5910), .A1(AOPB[19]), .B0(n15153), .Y(n3260) );
  OAI21XL U27555 ( .A0(n5906), .A1(AOPB[18]), .B0(n15156), .Y(n3256) );
  OAI21XL U27556 ( .A0(n5836), .A1(n16504), .B0(n15159), .Y(n15160) );
  OAI21XL U27557 ( .A0(n6885), .A1(AOPB[17]), .B0(n15160), .Y(n3252) );
  OAI21XL U27558 ( .A0(n5905), .A1(AOPB[16]), .B0(n15163), .Y(n3248) );
  OAI21XL U27559 ( .A0(R7_valid), .A1(AOPB[15]), .B0(n15167), .Y(n3244) );
  OAI21XL U27560 ( .A0(n5910), .A1(AOPB[14]), .B0(n15170), .Y(n3240) );
  OAI21XL U27561 ( .A0(n6885), .A1(AOPB[13]), .B0(n15174), .Y(n3236) );
  OAI21XL U27562 ( .A0(n5912), .A1(AOPB[12]), .B0(n15178), .Y(n3232) );
  OAI21XL U27563 ( .A0(n6884), .A1(AOPB[11]), .B0(n15182), .Y(n3228) );
  OAI21XL U27564 ( .A0(n5912), .A1(AOPB[10]), .B0(n15186), .Y(n3224) );
  OAI21XL U27565 ( .A0(n6884), .A1(AOPB[9]), .B0(n15190), .Y(n3424) );
  OAI21XL U27566 ( .A0(n5905), .A1(AOPB[8]), .B0(n15193), .Y(n3420) );
  OAI21XL U27567 ( .A0(n5908), .A1(AOPB[7]), .B0(n15196), .Y(n3416) );
  OAI21XL U27568 ( .A0(n5912), .A1(AOPB[6]), .B0(n15199), .Y(n3412) );
  OAI21XL U27569 ( .A0(n6883), .A1(AOPB[5]), .B0(n15202), .Y(n3408) );
  OAI21XL U27570 ( .A0(n5913), .A1(AOPB[4]), .B0(n15205), .Y(n3396) );
  OAI21XL U27571 ( .A0(n5908), .A1(AOPB[3]), .B0(n15209), .Y(n3352) );
  OAI21XL U27572 ( .A0(n5907), .A1(AOPB[2]), .B0(n15213), .Y(n3308) );
  OAI21XL U27573 ( .A0(n15218), .A1(n16567), .B0(n15217), .Y(n15219) );
  OAI21XL U27574 ( .A0(n6884), .A1(AOPB[1]), .B0(n15219), .Y(n3264) );
  OAI21XL U27575 ( .A0(n5917), .A1(AOPB[0]), .B0(n15222), .Y(n3220) );
  OAI21XL U27576 ( .A0(n5906), .A1(BOPA[51]), .B0(n15225), .Y(n3823) );
  OAI21XL U27577 ( .A0(n6883), .A1(BOPA[25]), .B0(n15228), .Y(n3707) );
  NAND3XL U27578 ( .A(n7305), .B(cnt[9]), .C(n6880), .Y(n5696) );
  OAI21XL U27579 ( .A0(n5906), .A1(BOPA[50]), .B0(n15232), .Y(n3819) );
  OAI21XL U27580 ( .A0(R7_valid), .A1(BOPA[24]), .B0(n15235), .Y(n3703) );
  OAI21XL U27581 ( .A0(n6880), .A1(BOPA[49]), .B0(n15238), .Y(n3811) );
  OAI21XL U27582 ( .A0(n5908), .A1(BOPA[23]), .B0(n15242), .Y(n3699) );
  OAI21XL U27583 ( .A0(n5912), .A1(BOPA[48]), .B0(n15245), .Y(n3807) );
  OAI21XL U27584 ( .A0(n6880), .A1(BOPA[22]), .B0(n15249), .Y(n3695) );
  OAI21XL U27585 ( .A0(n5917), .A1(BOPA[47]), .B0(n15253), .Y(n3803) );
  OAI21XL U27586 ( .A0(n6883), .A1(BOPA[21]), .B0(n15257), .Y(n3691) );
  OAI21XL U27587 ( .A0(n5908), .A1(BOPA[46]), .B0(n15261), .Y(n3799) );
  OAI21XL U27588 ( .A0(n5907), .A1(BOPA[20]), .B0(n15265), .Y(n3687) );
  OAI21XL U27589 ( .A0(n5908), .A1(BOPA[45]), .B0(n15269), .Y(n3795) );
  OAI21XL U27590 ( .A0(n5907), .A1(BOPA[19]), .B0(n15273), .Y(n3679) );
  OAI21XL U27591 ( .A0(n5912), .A1(BOPA[44]), .B0(n15277), .Y(n3791) );
  OAI21XL U27592 ( .A0(n5913), .A1(BOPA[18]), .B0(n15280), .Y(n3675) );
  OAI21XL U27593 ( .A0(n6884), .A1(BOPA[43]), .B0(n15283), .Y(n3787) );
  OAI21XL U27594 ( .A0(n5907), .A1(BOPA[17]), .B0(n15287), .Y(n3671) );
  OAI21XL U27595 ( .A0(n6884), .A1(BOPA[42]), .B0(n15291), .Y(n3783) );
  OAI21XL U27596 ( .A0(n5906), .A1(BOPA[16]), .B0(n15295), .Y(n3667) );
  OAI21XL U27597 ( .A0(n5910), .A1(BOPA[41]), .B0(n15298), .Y(n3779) );
  OAI21XL U27598 ( .A0(n5912), .A1(BOPA[15]), .B0(n15302), .Y(n3663) );
  OAI21XL U27599 ( .A0(n5908), .A1(BOPA[40]), .B0(n15305), .Y(n3775) );
  OAI21XL U27600 ( .A0(n5906), .A1(BOPA[14]), .B0(n15309), .Y(n3659) );
  OAI21XL U27601 ( .A0(n5908), .A1(BOPA[39]), .B0(n15313), .Y(n3767) );
  OAI21XL U27602 ( .A0(n6883), .A1(BOPA[13]), .B0(n15317), .Y(n3655) );
  OAI21XL U27603 ( .A0(n5908), .A1(BOPA[38]), .B0(n15321), .Y(n3763) );
  OAI21XL U27604 ( .A0(n5908), .A1(BOPA[12]), .B0(n15325), .Y(n3651) );
  OAI21XL U27605 ( .A0(n6881), .A1(BOPA[37]), .B0(n15329), .Y(n3759) );
  OAI21XL U27606 ( .A0(n5910), .A1(BOPA[11]), .B0(n15333), .Y(n3647) );
  OAI21XL U27607 ( .A0(n5907), .A1(BOPA[36]), .B0(n15336), .Y(n3755) );
  OAI21XL U27608 ( .A0(n5907), .A1(BOPA[10]), .B0(n15340), .Y(n3643) );
  OAI21XL U27609 ( .A0(n6880), .A1(BOPA[9]), .B0(n15344), .Y(n3843) );
  OAI21XL U27610 ( .A0(n5907), .A1(BOPA[8]), .B0(n15348), .Y(n3839) );
  OAI21XL U27611 ( .A0(n5917), .A1(BOPA[7]), .B0(n15353), .Y(n3835) );
  OAI21XL U27612 ( .A0(n5908), .A1(BOPA[6]), .B0(n15357), .Y(n3831) );
  OAI21XL U27613 ( .A0(n5915), .A1(BOPA[31]), .B0(n15360), .Y(n3735) );
  OAI21XL U27614 ( .A0(n5909), .A1(BOPA[5]), .B0(n15364), .Y(n3827) );
  OAI21XL U27615 ( .A0(n5910), .A1(BOPA[30]), .B0(n15367), .Y(n3731) );
  OAI21XL U27616 ( .A0(n5910), .A1(BOPA[4]), .B0(n15370), .Y(n3815) );
  OAI21XL U27617 ( .A0(n5912), .A1(BOPA[29]), .B0(n15374), .Y(n3723) );
  OAI21XL U27618 ( .A0(n5907), .A1(BOPA[3]), .B0(n15377), .Y(n3771) );
  OAI21XL U27619 ( .A0(n5910), .A1(BOPA[2]), .B0(n15381), .Y(n3727) );
  OAI21XL U27620 ( .A0(n6881), .A1(BOPA[1]), .B0(n15384), .Y(n3683) );
  OAI21XL U27621 ( .A0(n6881), .A1(BOPA[0]), .B0(n15388), .Y(n3639) );
  NAND2X1 U27622 ( .A(n28671), .B(D_sel_reg_4__0_), .Y(n16163) );
  NOR2X1 U27623 ( .A(D_sel_reg_4__0_), .B(n28671), .Y(n15431) );
  OAI21XL U27624 ( .A0(n5910), .A1(BOPD[51]), .B0(n15391), .Y(n3822) );
  OAI21XL U27625 ( .A0(n5907), .A1(BOPD[50]), .B0(n15395), .Y(n3818) );
  OAI21XL U27626 ( .A0(n6884), .A1(BOPD[49]), .B0(n15399), .Y(n3810) );
  OAI21XL U27627 ( .A0(n6884), .A1(BOPD[48]), .B0(n15403), .Y(n3806) );
  OAI21XL U27628 ( .A0(n5908), .A1(BOPD[47]), .B0(n15406), .Y(n3802) );
  OAI21XL U27629 ( .A0(n5908), .A1(BOPD[46]), .B0(n15410), .Y(n3798) );
  OAI21XL U27630 ( .A0(n5912), .A1(BOPD[45]), .B0(n15413), .Y(n3794) );
  OAI21XL U27631 ( .A0(n5905), .A1(BOPD[44]), .B0(n15417), .Y(n3790) );
  OAI21XL U27632 ( .A0(n5913), .A1(BOPD[43]), .B0(n15420), .Y(n3786) );
  OAI21XL U27633 ( .A0(n6883), .A1(BOPD[42]), .B0(n15424), .Y(n3782) );
  AOI21XL U27634 ( .A0(B6_q[41]), .A1(n16161), .B0(n28985), .Y(n15425) );
  OAI21XL U27635 ( .A0(n5907), .A1(BOPD[41]), .B0(n15427), .Y(n3778) );
  AOI21XL U27636 ( .A0(B4_q[40]), .A1(n5933), .B0(n28985), .Y(n15428) );
  OAI21XL U27637 ( .A0(n5912), .A1(BOPD[40]), .B0(n15430), .Y(n3774) );
  OAI21XL U27638 ( .A0(n6882), .A1(BOPD[39]), .B0(n15435), .Y(n3766) );
  OAI21XL U27639 ( .A0(n5906), .A1(BOPD[38]), .B0(n15439), .Y(n3762) );
  OAI21XL U27640 ( .A0(n6882), .A1(BOPD[37]), .B0(n15443), .Y(n3758) );
  OAI21XL U27641 ( .A0(n5913), .A1(BOPD[36]), .B0(n15447), .Y(n3754) );
  OAI21XL U27642 ( .A0(n5913), .A1(BOPD[35]), .B0(n15451), .Y(n3750) );
  OAI21XL U27643 ( .A0(n6882), .A1(BOPD[34]), .B0(n15454), .Y(n3746) );
  OAI21XL U27644 ( .A0(n5912), .A1(BOPD[33]), .B0(n15457), .Y(n3742) );
  OAI21XL U27645 ( .A0(n5917), .A1(BOPD[32]), .B0(n15460), .Y(n3738) );
  OAI21XL U27646 ( .A0(n6885), .A1(BOPD[31]), .B0(n15463), .Y(n3734) );
  OAI21XL U27647 ( .A0(n5905), .A1(BOPD[30]), .B0(n15466), .Y(n3730) );
  OAI21XL U27648 ( .A0(n5905), .A1(BOPD[29]), .B0(n15470), .Y(n3722) );
  OAI21XL U27649 ( .A0(n5907), .A1(BOPD[28]), .B0(n15473), .Y(n3718) );
  OAI21XL U27650 ( .A0(n5913), .A1(BOPD[27]), .B0(n15477), .Y(n3714) );
  OAI21XL U27651 ( .A0(n6881), .A1(BOPD[26]), .B0(n15481), .Y(n3710) );
  OAI21XL U27652 ( .A0(R7_valid), .A1(BOPD[25]), .B0(n15485), .Y(n3706) );
  OAI21XL U27653 ( .A0(n5906), .A1(BOPD[24]), .B0(n15488), .Y(n3702) );
  OAI21XL U27654 ( .A0(n5913), .A1(BOPD[23]), .B0(n15492), .Y(n3698) );
  OAI21XL U27655 ( .A0(n6884), .A1(BOPD[22]), .B0(n15496), .Y(n3694) );
  OAI21XL U27656 ( .A0(n5907), .A1(BOPD[21]), .B0(n15500), .Y(n3690) );
  OAI21XL U27657 ( .A0(R7_valid), .A1(BOPD[20]), .B0(n15504), .Y(n3686) );
  OAI21XL U27658 ( .A0(n5917), .A1(BOPD[19]), .B0(n15508), .Y(n3678) );
  OAI21XL U27659 ( .A0(n5910), .A1(BOPD[18]), .B0(n15511), .Y(n3674) );
  OAI21XL U27660 ( .A0(n5905), .A1(BOPD[17]), .B0(n15515), .Y(n3670) );
  OAI21XL U27661 ( .A0(n6880), .A1(BOPD[16]), .B0(n15519), .Y(n3666) );
  OAI21XL U27662 ( .A0(n6881), .A1(BOPD[15]), .B0(n15523), .Y(n3662) );
  OAI21XL U27663 ( .A0(n5905), .A1(BOPD[14]), .B0(n15527), .Y(n3658) );
  OAI21XL U27664 ( .A0(n6885), .A1(BOPD[13]), .B0(n15530), .Y(n3654) );
  OAI21XL U27665 ( .A0(n6885), .A1(BOPD[12]), .B0(n15534), .Y(n3650) );
  OAI21XL U27666 ( .A0(n5906), .A1(BOPD[11]), .B0(n15538), .Y(n3646) );
  OAI21XL U27667 ( .A0(R7_valid), .A1(BOPD[10]), .B0(n15542), .Y(n3642) );
  OAI21XL U27668 ( .A0(n5917), .A1(BOPD[9]), .B0(n15546), .Y(n3842) );
  OAI21XL U27669 ( .A0(n6882), .A1(BOPD[8]), .B0(n15549), .Y(n3838) );
  OAI21XL U27670 ( .A0(R7_valid), .A1(BOPD[7]), .B0(n15552), .Y(n3834) );
  OAI21XL U27671 ( .A0(n5910), .A1(BOPD[6]), .B0(n15556), .Y(n3830) );
  OAI21XL U27672 ( .A0(n6882), .A1(BOPD[5]), .B0(n15561), .Y(n3826) );
  OAI21XL U27673 ( .A0(n6884), .A1(BOPD[4]), .B0(n15564), .Y(n3814) );
  OAI21XL U27674 ( .A0(n6882), .A1(BOPD[3]), .B0(n15567), .Y(n3770) );
  OAI21XL U27675 ( .A0(n6886), .A1(BOPD[2]), .B0(n15571), .Y(n3726) );
  OAI21XL U27676 ( .A0(n5907), .A1(BOPD[1]), .B0(n15575), .Y(n3682) );
  OAI21XL U27677 ( .A0(n5917), .A1(BOPD[0]), .B0(n15579), .Y(n3638) );
  CLKINVX3 U27678 ( .A(n16245), .Y(n16277) );
  OAI21XL U27679 ( .A0(n5906), .A1(BOPC[51]), .B0(n15582), .Y(n3821) );
  OAI21XL U27680 ( .A0(n5910), .A1(BOPC[50]), .B0(n15586), .Y(n3817) );
  OAI21XL U27681 ( .A0(n6885), .A1(BOPC[49]), .B0(n15589), .Y(n3809) );
  OAI21XL U27682 ( .A0(n6881), .A1(BOPC[48]), .B0(n15592), .Y(n3805) );
  OAI21XL U27683 ( .A0(n5910), .A1(BOPC[47]), .B0(n15596), .Y(n3801) );
  OAI21XL U27684 ( .A0(n5908), .A1(BOPC[46]), .B0(n15600), .Y(n3797) );
  OAI21XL U27685 ( .A0(n6881), .A1(BOPC[45]), .B0(n15603), .Y(n3793) );
  OAI21XL U27686 ( .A0(n5917), .A1(BOPC[44]), .B0(n15607), .Y(n3789) );
  OAI21XL U27687 ( .A0(n6885), .A1(BOPC[43]), .B0(n15611), .Y(n3785) );
  OAI21XL U27688 ( .A0(n5907), .A1(BOPC[42]), .B0(n15615), .Y(n3781) );
  OAI21XL U27689 ( .A0(R7_valid), .A1(BOPC[41]), .B0(n15618), .Y(n3777) );
  OAI21XL U27690 ( .A0(n5905), .A1(BOPC[40]), .B0(n15621), .Y(n3773) );
  OAI21XL U27691 ( .A0(n5905), .A1(BOPC[39]), .B0(n15624), .Y(n3765) );
  OAI21XL U27692 ( .A0(n6885), .A1(BOPC[38]), .B0(n15628), .Y(n3761) );
  OAI21XL U27693 ( .A0(n5912), .A1(BOPC[37]), .B0(n15632), .Y(n3757) );
  INVX1 U27694 ( .A(R7_valid), .Y(n16564) );
  OAI21XL U27695 ( .A0(n5907), .A1(BOPC[36]), .B0(n15636), .Y(n3753) );
  OAI21XL U27696 ( .A0(n6884), .A1(BOPC[35]), .B0(n15640), .Y(n3749) );
  OAI21XL U27697 ( .A0(n5908), .A1(BOPC[34]), .B0(n15644), .Y(n3745) );
  OAI21XL U27698 ( .A0(n6886), .A1(BOPC[33]), .B0(n15647), .Y(n3741) );
  INVX1 U27699 ( .A(R7_valid), .Y(n16487) );
  OAI21XL U27700 ( .A0(n5905), .A1(BOPC[32]), .B0(n15651), .Y(n3737) );
  OAI21XL U27701 ( .A0(n5910), .A1(BOPC[31]), .B0(n15654), .Y(n3733) );
  OAI21XL U27702 ( .A0(n5917), .A1(BOPC[30]), .B0(n15657), .Y(n3729) );
  OAI21XL U27703 ( .A0(n5910), .A1(BOPC[29]), .B0(n15661), .Y(n3721) );
  OAI21XL U27704 ( .A0(n5910), .A1(BOPC[28]), .B0(n15665), .Y(n3717) );
  OAI21XL U27705 ( .A0(n5905), .A1(BOPC[27]), .B0(n15669), .Y(n3713) );
  OAI21XL U27706 ( .A0(n6881), .A1(BOPC[26]), .B0(n15672), .Y(n3709) );
  OAI21XL U27707 ( .A0(n5908), .A1(BOPC[25]), .B0(n15675), .Y(n3705) );
  OAI21XL U27708 ( .A0(n5907), .A1(BOPC[24]), .B0(n15678), .Y(n3701) );
  OAI21XL U27709 ( .A0(n5905), .A1(BOPC[23]), .B0(n15682), .Y(n3697) );
  OAI21XL U27710 ( .A0(n5908), .A1(BOPC[22]), .B0(n15686), .Y(n3693) );
  OAI21XL U27711 ( .A0(n5917), .A1(BOPC[21]), .B0(n15691), .Y(n3689) );
  OAI21XL U27712 ( .A0(n5908), .A1(BOPC[20]), .B0(n15694), .Y(n3685) );
  OAI21XL U27713 ( .A0(n6881), .A1(BOPC[19]), .B0(n15698), .Y(n3677) );
  OAI21XL U27714 ( .A0(n6884), .A1(BOPC[18]), .B0(n15702), .Y(n3673) );
  OAI21XL U27715 ( .A0(n5908), .A1(BOPC[17]), .B0(n15706), .Y(n3669) );
  OAI21XL U27716 ( .A0(n5905), .A1(BOPC[16]), .B0(n15710), .Y(n3665) );
  OAI21XL U27717 ( .A0(n6881), .A1(BOPC[15]), .B0(n15714), .Y(n3661) );
  OAI21XL U27718 ( .A0(n5905), .A1(BOPC[14]), .B0(n15718), .Y(n3657) );
  OAI21XL U27719 ( .A0(n5908), .A1(BOPC[13]), .B0(n15722), .Y(n3653) );
  OAI21XL U27720 ( .A0(n6881), .A1(BOPC[12]), .B0(n15726), .Y(n3649) );
  OAI21XL U27721 ( .A0(n5912), .A1(BOPC[11]), .B0(n15730), .Y(n3645) );
  OAI21XL U27722 ( .A0(n5907), .A1(BOPC[10]), .B0(n15734), .Y(n3641) );
  OAI21XL U27723 ( .A0(n6881), .A1(BOPC[9]), .B0(n15738), .Y(n3841) );
  OAI21XL U27724 ( .A0(n5910), .A1(BOPC[8]), .B0(n15742), .Y(n3837) );
  OAI21XL U27725 ( .A0(n6884), .A1(BOPC[7]), .B0(n15746), .Y(n3833) );
  OAI21XL U27726 ( .A0(R7_valid), .A1(BOPC[6]), .B0(n15751), .Y(n3829) );
  OAI21XL U27727 ( .A0(n5910), .A1(BOPC[5]), .B0(n15755), .Y(n3825) );
  OAI21XL U27728 ( .A0(n5908), .A1(BOPC[4]), .B0(n15759), .Y(n3813) );
  OAI21XL U27729 ( .A0(n5910), .A1(BOPC[3]), .B0(n15762), .Y(n3769) );
  OAI21XL U27730 ( .A0(n5907), .A1(BOPC[2]), .B0(n15766), .Y(n3725) );
  OAI21XL U27731 ( .A0(n5910), .A1(BOPC[1]), .B0(n15769), .Y(n3681) );
  OAI21XL U27732 ( .A0(n5800), .A1(BOPC[0]), .B0(n15772), .Y(n3637) );
  OAI21XL U27733 ( .A0(n5913), .A1(BOPB[51]), .B0(n15776), .Y(n3820) );
  OAI21XL U27734 ( .A0(n5912), .A1(BOPB[50]), .B0(n15780), .Y(n3816) );
  OAI21XL U27735 ( .A0(n5905), .A1(BOPB[49]), .B0(n15784), .Y(n3808) );
  OAI21XL U27736 ( .A0(n5910), .A1(BOPB[48]), .B0(n15788), .Y(n3804) );
  OAI21XL U27737 ( .A0(n5905), .A1(BOPB[47]), .B0(n15792), .Y(n3800) );
  OAI21XL U27738 ( .A0(R7_valid), .A1(BOPB[46]), .B0(n15796), .Y(n3796) );
  OAI21XL U27739 ( .A0(n5910), .A1(BOPB[45]), .B0(n15800), .Y(n3792) );
  OAI21XL U27740 ( .A0(n5917), .A1(BOPB[44]), .B0(n15804), .Y(n3788) );
  OAI21XL U27741 ( .A0(n5905), .A1(BOPB[43]), .B0(n15808), .Y(n3784) );
  OAI21XL U27742 ( .A0(n5917), .A1(BOPB[42]), .B0(n15812), .Y(n3780) );
  OAI21XL U27743 ( .A0(n5905), .A1(BOPB[41]), .B0(n15816), .Y(n3776) );
  OAI21XL U27744 ( .A0(n5917), .A1(BOPB[40]), .B0(n15820), .Y(n3772) );
  OAI21XL U27745 ( .A0(n5907), .A1(BOPB[39]), .B0(n15824), .Y(n3764) );
  OAI21XL U27746 ( .A0(n5913), .A1(BOPB[38]), .B0(n15828), .Y(n3760) );
  OAI21XL U27747 ( .A0(n6883), .A1(BOPB[37]), .B0(n15832), .Y(n3756) );
  OAI21XL U27748 ( .A0(n5910), .A1(BOPB[36]), .B0(n15836), .Y(n3752) );
  OAI21XL U27749 ( .A0(n5906), .A1(BOPB[35]), .B0(n15840), .Y(n3748) );
  OAI21XL U27750 ( .A0(n6881), .A1(BOPB[34]), .B0(n15844), .Y(n3744) );
  OAI21XL U27751 ( .A0(n5906), .A1(BOPB[33]), .B0(n15848), .Y(n3740) );
  OAI21XL U27752 ( .A0(n5912), .A1(BOPB[32]), .B0(n15852), .Y(n3736) );
  OAI21XL U27753 ( .A0(n6880), .A1(BOPB[31]), .B0(n15856), .Y(n3732) );
  OAI21XL U27754 ( .A0(n5913), .A1(BOPB[30]), .B0(n15860), .Y(n3728) );
  OAI21XL U27755 ( .A0(n5906), .A1(BOPB[29]), .B0(n15864), .Y(n3720) );
  OAI21XL U27756 ( .A0(n5908), .A1(BOPB[28]), .B0(n15868), .Y(n3716) );
  OAI21XL U27757 ( .A0(n6886), .A1(BOPB[27]), .B0(n15872), .Y(n3712) );
  OAI21XL U27758 ( .A0(n6886), .A1(BOPB[26]), .B0(n15876), .Y(n3708) );
  OAI21XL U27759 ( .A0(n5912), .A1(BOPB[25]), .B0(n15880), .Y(n3704) );
  OAI21XL U27760 ( .A0(n6881), .A1(BOPB[24]), .B0(n15884), .Y(n3700) );
  OAI21XL U27761 ( .A0(n5906), .A1(BOPB[23]), .B0(n15888), .Y(n3696) );
  OAI21XL U27762 ( .A0(n6886), .A1(BOPB[22]), .B0(n15892), .Y(n3692) );
  OAI21XL U27763 ( .A0(n5905), .A1(BOPB[21]), .B0(n15896), .Y(n3688) );
  OAI21XL U27764 ( .A0(n6881), .A1(BOPB[20]), .B0(n15900), .Y(n3684) );
  OAI21XL U27765 ( .A0(n5912), .A1(BOPB[19]), .B0(n15904), .Y(n3676) );
  OAI21XL U27766 ( .A0(n5906), .A1(BOPB[18]), .B0(n15908), .Y(n3672) );
  OAI21XL U27767 ( .A0(n6886), .A1(BOPB[17]), .B0(n15912), .Y(n3668) );
  OAI21XL U27768 ( .A0(n6882), .A1(BOPB[16]), .B0(n15916), .Y(n3664) );
  OAI21XL U27769 ( .A0(n5913), .A1(BOPB[15]), .B0(n15920), .Y(n3660) );
  OAI21XL U27770 ( .A0(n6882), .A1(BOPB[14]), .B0(n15924), .Y(n3656) );
  OAI21XL U27771 ( .A0(n5913), .A1(BOPB[13]), .B0(n15928), .Y(n3652) );
  OAI21XL U27772 ( .A0(n5913), .A1(BOPB[12]), .B0(n15932), .Y(n3648) );
  OAI21XL U27773 ( .A0(n5910), .A1(BOPB[11]), .B0(n15936), .Y(n3644) );
  OAI21XL U27774 ( .A0(n6882), .A1(BOPB[10]), .B0(n15940), .Y(n3640) );
  OAI21XL U27775 ( .A0(n5907), .A1(BOPB[9]), .B0(n15944), .Y(n3840) );
  OAI21XL U27776 ( .A0(n6886), .A1(BOPB[8]), .B0(n15949), .Y(n3836) );
  OAI21XL U27777 ( .A0(n5915), .A1(BOPB[7]), .B0(n15953), .Y(n3832) );
  OAI21XL U27778 ( .A0(n6881), .A1(BOPB[6]), .B0(n15957), .Y(n3828) );
  OAI21XL U27779 ( .A0(n5800), .A1(BOPB[5]), .B0(n15962), .Y(n3824) );
  OAI21XL U27780 ( .A0(n5905), .A1(BOPB[4]), .B0(n15968), .Y(n3812) );
  OAI21XL U27781 ( .A0(n5800), .A1(BOPB[3]), .B0(n15973), .Y(n3768) );
  OAI21XL U27782 ( .A0(n5905), .A1(BOPB[2]), .B0(n15977), .Y(n3724) );
  OAI21XL U27783 ( .A0(n6882), .A1(BOPB[1]), .B0(n15981), .Y(n3680) );
  OAI21XL U27784 ( .A0(n6882), .A1(BOPB[0]), .B0(n15986), .Y(n3636) );
  OAI21XL U27785 ( .A0(n16361), .A1(n16154), .B0(n5906), .Y(n15987) );
  OAI21XL U27786 ( .A0(n5800), .A1(AOPD[50]), .B0(n15992), .Y(n3402) );
  OAI21XL U27787 ( .A0(n5907), .A1(AOPD[49]), .B0(n15996), .Y(n3394) );
  OAI21XL U27788 ( .A0(n6882), .A1(AOPD[48]), .B0(n15999), .Y(n3390) );
  OAI21XL U27789 ( .A0(n5913), .A1(AOPD[47]), .B0(n16002), .Y(n3386) );
  OAI21XL U27790 ( .A0(n5913), .A1(AOPD[46]), .B0(n16006), .Y(n3382) );
  OAI21XL U27791 ( .A0(n16386), .A1(n16154), .B0(n5909), .Y(n16007) );
  OAI21XL U27792 ( .A0(n16390), .A1(n5806), .B0(n5910), .Y(n16010) );
  OAI21XL U27793 ( .A0(n6882), .A1(AOPD[43]), .B0(n16016), .Y(n3370) );
  OAI21XL U27794 ( .A0(n6882), .A1(AOPD[42]), .B0(n16019), .Y(n3366) );
  OAI21XL U27795 ( .A0(n5912), .A1(AOPD[41]), .B0(n16022), .Y(n3362) );
  OAI21XL U27796 ( .A0(n5907), .A1(AOPD[40]), .B0(n16025), .Y(n3358) );
  OAI21XL U27797 ( .A0(n16410), .A1(n5806), .B0(n6880), .Y(n16026) );
  OAI2BB2XL U27798 ( .B0(n5909), .B1(AOPD[39]), .A0N(n16028), .A1N(n16027), 
        .Y(n3350) );
  OAI21XL U27799 ( .A0(n16414), .A1(n16154), .B0(n5917), .Y(n16029) );
  OAI2BB2XL U27800 ( .B0(n5915), .B1(AOPD[38]), .A0N(n16031), .A1N(n16030), 
        .Y(n3346) );
  OAI21XL U27801 ( .A0(n5913), .A1(AOPD[37]), .B0(n16035), .Y(n3342) );
  OAI21XL U27802 ( .A0(n5913), .A1(AOPD[36]), .B0(n16039), .Y(n3338) );
  OAI21XL U27803 ( .A0(n16427), .A1(n16154), .B0(n5800), .Y(n16040) );
  OAI2BB2XL U27804 ( .B0(n5909), .B1(AOPD[35]), .A0N(n16042), .A1N(n16041), 
        .Y(n3334) );
  OAI21XL U27805 ( .A0(n5913), .A1(AOPD[34]), .B0(n16045), .Y(n3330) );
  OAI21XL U27806 ( .A0(n5917), .A1(AOPD[33]), .B0(n16049), .Y(n3326) );
  OAI21XL U27807 ( .A0(n16163), .A1(n16439), .B0(n16052), .Y(n16053) );
  OAI21XL U27808 ( .A0(n6881), .A1(AOPD[32]), .B0(n16053), .Y(n3322) );
  OAI21XL U27809 ( .A0(n6882), .A1(AOPD[31]), .B0(n16057), .Y(n3318) );
  OAI21XL U27810 ( .A0(n5905), .A1(AOPD[30]), .B0(n16060), .Y(n3314) );
  OAI21XL U27811 ( .A0(n6882), .A1(AOPD[29]), .B0(n16064), .Y(n3306) );
  OAI21XL U27812 ( .A0(n5905), .A1(AOPD[28]), .B0(n16067), .Y(n3302) );
  OAI21XL U27813 ( .A0(n16163), .A1(n16459), .B0(n16070), .Y(n16071) );
  OAI21XL U27814 ( .A0(R7_valid), .A1(AOPD[27]), .B0(n16071), .Y(n3298) );
  OAI21XL U27815 ( .A0(n5907), .A1(AOPD[26]), .B0(n16074), .Y(n3294) );
  OAI21XL U27816 ( .A0(n16468), .A1(n16154), .B0(n5913), .Y(n16075) );
  OAI21XL U27817 ( .A0(n5907), .A1(AOPD[24]), .B0(n16080), .Y(n3286) );
  OAI21XL U27818 ( .A0(R7_valid), .A1(AOPD[23]), .B0(n16083), .Y(n3282) );
  OAI21XL U27819 ( .A0(n5905), .A1(AOPD[22]), .B0(n16087), .Y(n3278) );
  OAI21XL U27820 ( .A0(n6884), .A1(AOPD[21]), .B0(n16090), .Y(n3274) );
  OAI21XL U27821 ( .A0(n5906), .A1(AOPD[20]), .B0(n16094), .Y(n3270) );
  OAI21XL U27822 ( .A0(n16494), .A1(n5806), .B0(n5912), .Y(n16095) );
  OAI21XL U27823 ( .A0(n5908), .A1(AOPD[18]), .B0(n16100), .Y(n3258) );
  OAI21XL U27824 ( .A0(n6880), .A1(AOPD[17]), .B0(n16104), .Y(n3254) );
  OAI21XL U27825 ( .A0(n6886), .A1(AOPD[16]), .B0(n16108), .Y(n3250) );
  OAI21XL U27826 ( .A0(n5908), .A1(AOPD[15]), .B0(n16112), .Y(n3246) );
  OAI21XL U27827 ( .A0(n5912), .A1(AOPD[14]), .B0(n16115), .Y(n3242) );
  OAI21XL U27828 ( .A0(n5800), .A1(AOPD[13]), .B0(n16118), .Y(n3238) );
  OAI21XL U27829 ( .A0(n5913), .A1(AOPD[12]), .B0(n16121), .Y(n3234) );
  OAI21XL U27830 ( .A0(n5906), .A1(AOPD[11]), .B0(n16124), .Y(n3230) );
  OAI21XL U27831 ( .A0(n5906), .A1(AOPD[10]), .B0(n16127), .Y(n3226) );
  OAI21XL U27832 ( .A0(n5912), .A1(AOPD[9]), .B0(n16131), .Y(n3426) );
  OAI21XL U27833 ( .A0(n6883), .A1(AOPD[8]), .B0(n16134), .Y(n3422) );
  OAI21XL U27834 ( .A0(n16543), .A1(n16163), .B0(R7_valid), .Y(n16135) );
  OAI21XL U27835 ( .A0(n5913), .A1(AOPD[6]), .B0(n16142), .Y(n3414) );
  OAI21XL U27836 ( .A0(n5906), .A1(AOPD[5]), .B0(n16146), .Y(n3410) );
  OAI21XL U27837 ( .A0(n5907), .A1(AOPD[4]), .B0(n16150), .Y(n3398) );
  OAI21XL U27838 ( .A0(n5906), .A1(AOPD[3]), .B0(n16153), .Y(n3354) );
  OAI21XL U27839 ( .A0(n16562), .A1(n16154), .B0(R7_valid), .Y(n16155) );
  OAI2BB2XL U27840 ( .B0(n5915), .B1(AOPD[2]), .A0N(n16157), .A1N(n16156), .Y(
        n3310) );
  OAI21XL U27841 ( .A0(n16163), .A1(n16567), .B0(n16162), .Y(n16164) );
  OAI21XL U27842 ( .A0(n6883), .A1(AOPD[1]), .B0(n16164), .Y(n3266) );
  OAI21XL U27843 ( .A0(n5907), .A1(AOPD[0]), .B0(n16169), .Y(n3222) );
  OAI21XL U27844 ( .A0(n16361), .A1(n16245), .B0(n5917), .Y(n16170) );
  OAI21XL U27845 ( .A0(n5909), .A1(AOPC[50]), .B0(n16175), .Y(n3401) );
  OAI21XL U27846 ( .A0(n5906), .A1(AOPC[49]), .B0(n16178), .Y(n3393) );
  OAI21XL U27847 ( .A0(n6883), .A1(AOPC[48]), .B0(n16181), .Y(n3389) );
  OAI21XL U27848 ( .A0(n5906), .A1(AOPC[47]), .B0(n16184), .Y(n3385) );
  OAI21XL U27849 ( .A0(n5813), .A1(n16382), .B0(n16187), .Y(n16188) );
  OAI21XL U27850 ( .A0(n5913), .A1(AOPC[46]), .B0(n16188), .Y(n3381) );
  OAI21XL U27851 ( .A0(n5915), .A1(AOPC[45]), .B0(n16192), .Y(n3377) );
  OAI21XL U27852 ( .A0(n5906), .A1(AOPC[44]), .B0(n16195), .Y(n3373) );
  OAI21XL U27853 ( .A0(n5913), .A1(AOPC[43]), .B0(n16199), .Y(n3369) );
  OAI21XL U27854 ( .A0(n5906), .A1(AOPC[42]), .B0(n16202), .Y(n3365) );
  OAI21XL U27855 ( .A0(n5917), .A1(AOPC[41]), .B0(n16206), .Y(n3361) );
  OAI21XL U27856 ( .A0(n6885), .A1(AOPC[40]), .B0(n16209), .Y(n3357) );
  OAI21XL U27857 ( .A0(n5917), .A1(AOPC[39]), .B0(n16212), .Y(n3349) );
  OAI21XL U27858 ( .A0(n5905), .A1(AOPC[38]), .B0(n16216), .Y(n3345) );
  OAI21XL U27859 ( .A0(n16419), .A1(n16245), .B0(R7_valid), .Y(n16217) );
  OAI2BB2XL U27860 ( .B0(n5915), .B1(AOPC[37]), .A0N(n16219), .A1N(n16218), 
        .Y(n3341) );
  OAI21XL U27861 ( .A0(n5908), .A1(AOPC[36]), .B0(n16223), .Y(n3337) );
  OAI21XL U27862 ( .A0(n5912), .A1(AOPC[35]), .B0(n16227), .Y(n3333) );
  OAI21XL U27863 ( .A0(n6884), .A1(AOPC[34]), .B0(n16230), .Y(n3329) );
  OAI21XL U27864 ( .A0(n5917), .A1(AOPC[33]), .B0(n16233), .Y(n3325) );
  OAI21XL U27865 ( .A0(n5813), .A1(n16439), .B0(n16236), .Y(n16237) );
  OAI21XL U27866 ( .A0(n6881), .A1(AOPC[32]), .B0(n16237), .Y(n3321) );
  OAI21XL U27867 ( .A0(n5800), .A1(AOPC[31]), .B0(n16241), .Y(n3317) );
  OAI21XL U27868 ( .A0(n6886), .A1(AOPC[30]), .B0(n16244), .Y(n3313) );
  OAI21XL U27869 ( .A0(n16451), .A1(n16245), .B0(R7_valid), .Y(n16246) );
  OAI2BB2XL U27870 ( .B0(n5915), .B1(AOPC[29]), .A0N(n16248), .A1N(n16247), 
        .Y(n3305) );
  OAI21XL U27871 ( .A0(n5912), .A1(AOPC[28]), .B0(n16252), .Y(n3301) );
  OAI21XL U27872 ( .A0(n6886), .A1(AOPC[27]), .B0(n16256), .Y(n3297) );
  OAI21XL U27873 ( .A0(n5917), .A1(AOPC[26]), .B0(n16260), .Y(n3293) );
  OAI21XL U27874 ( .A0(n6886), .A1(AOPC[25]), .B0(n16264), .Y(n3289) );
  OAI21XL U27875 ( .A0(n6886), .A1(AOPC[24]), .B0(n16267), .Y(n3285) );
  OAI21XL U27876 ( .A0(n5917), .A1(AOPC[23]), .B0(n16270), .Y(n3281) );
  OAI21XL U27877 ( .A0(n5912), .A1(AOPC[22]), .B0(n16273), .Y(n3277) );
  OAI21XL U27878 ( .A0(n5913), .A1(AOPC[21]), .B0(n16276), .Y(n3273) );
  OAI21XL U27879 ( .A0(n5913), .A1(AOPC[20]), .B0(n16281), .Y(n3269) );
  OAI21XL U27880 ( .A0(n5908), .A1(AOPC[19]), .B0(n16284), .Y(n3261) );
  OAI21XL U27881 ( .A0(n6886), .A1(AOPC[18]), .B0(n16288), .Y(n3257) );
  OAI21XL U27882 ( .A0(n5813), .A1(n16504), .B0(n16291), .Y(n16292) );
  OAI21XL U27883 ( .A0(n6886), .A1(AOPC[17]), .B0(n16292), .Y(n3253) );
  OAI21XL U27884 ( .A0(n5917), .A1(AOPC[16]), .B0(n16296), .Y(n3249) );
  OAI21XL U27885 ( .A0(n5917), .A1(AOPC[15]), .B0(n16300), .Y(n3245) );
  OAI21XL U27886 ( .A0(n5912), .A1(AOPC[14]), .B0(n16304), .Y(n3241) );
  OAI21XL U27887 ( .A0(R7_valid), .A1(AOPC[13]), .B0(n16307), .Y(n3237) );
  OAI21XL U27888 ( .A0(n5917), .A1(AOPC[12]), .B0(n16310), .Y(n3233) );
  OAI21XL U27889 ( .A0(n6883), .A1(AOPC[11]), .B0(n16313), .Y(n3229) );
  OAI21XL U27890 ( .A0(n6881), .A1(AOPC[10]), .B0(n16316), .Y(n3225) );
  OAI21XL U27891 ( .A0(n5905), .A1(AOPC[9]), .B0(n16320), .Y(n3425) );
  OAI21XL U27892 ( .A0(n5912), .A1(AOPC[8]), .B0(n16324), .Y(n3421) );
  OAI21XL U27893 ( .A0(n6886), .A1(AOPC[7]), .B0(n16328), .Y(n3417) );
  OAI21XL U27894 ( .A0(n5906), .A1(AOPC[6]), .B0(n16332), .Y(n3413) );
  OAI21XL U27895 ( .A0(n5906), .A1(AOPC[5]), .B0(n16335), .Y(n3409) );
  OAI21XL U27896 ( .A0(n5907), .A1(AOPC[4]), .B0(n16339), .Y(n3397) );
  OAI21XL U27897 ( .A0(n6886), .A1(AOPC[3]), .B0(n16343), .Y(n3353) );
  OAI21XL U27898 ( .A0(n6882), .A1(AOPC[2]), .B0(n16349), .Y(n3309) );
  OAI21XL U27899 ( .A0(n5813), .A1(n16567), .B0(n16352), .Y(n16353) );
  OAI21XL U27900 ( .A0(n5912), .A1(AOPC[1]), .B0(n16353), .Y(n3265) );
  AOI21XL U27901 ( .A0(B0_q[0]), .A1(n15687), .B0(n28985), .Y(n16355) );
  OAI21XL U27902 ( .A0(n5912), .A1(AOPC[0]), .B0(n16358), .Y(n3221) );
  OAI21XL U27903 ( .A0(n6886), .A1(AOPA[51]), .B0(n16362), .Y(n3407) );
  OAI21XL U27904 ( .A0(n5906), .A1(AOPA[50]), .B0(n16366), .Y(n3403) );
  OAI21XL U27905 ( .A0(n6881), .A1(AOPA[49]), .B0(n16370), .Y(n3395) );
  OAI21XL U27906 ( .A0(n5908), .A1(AOPA[48]), .B0(n16374), .Y(n3391) );
  OAI21XL U27907 ( .A0(n6885), .A1(AOPA[47]), .B0(n16379), .Y(n3387) );
  OAI21XL U27908 ( .A0(n5910), .A1(AOPA[46]), .B0(n16383), .Y(n3383) );
  OAI21XL U27909 ( .A0(n5910), .A1(AOPA[45]), .B0(n16387), .Y(n3379) );
  OAI21XL U27910 ( .A0(R7_valid), .A1(AOPA[44]), .B0(n16391), .Y(n3375) );
  OAI21XL U27911 ( .A0(n6882), .A1(AOPA[43]), .B0(n16395), .Y(n3371) );
  OAI21XL U27912 ( .A0(n5907), .A1(AOPA[42]), .B0(n16399), .Y(n3367) );
  OAI21XL U27913 ( .A0(R7_valid), .A1(AOPA[41]), .B0(n16403), .Y(n3363) );
  OAI21XL U27914 ( .A0(n5908), .A1(AOPA[40]), .B0(n16407), .Y(n3359) );
  OAI21XL U27915 ( .A0(n5906), .A1(AOPA[39]), .B0(n16411), .Y(n3351) );
  OAI21XL U27916 ( .A0(n6883), .A1(AOPA[38]), .B0(n16415), .Y(n3347) );
  OAI21XL U27917 ( .A0(n5907), .A1(AOPA[37]), .B0(n16420), .Y(n3343) );
  OAI21XL U27918 ( .A0(R7_valid), .A1(AOPA[36]), .B0(n16424), .Y(n3339) );
  OAI21XL U27919 ( .A0(n6882), .A1(AOPA[35]), .B0(n16428), .Y(n3335) );
  OAI21XL U27920 ( .A0(n5910), .A1(AOPA[34]), .B0(n16432), .Y(n3331) );
  OAI21XL U27921 ( .A0(n5917), .A1(AOPA[33]), .B0(n16436), .Y(n3327) );
  OAI21XL U27922 ( .A0(n5800), .A1(AOPA[32]), .B0(n16440), .Y(n3323) );
  OAI21XL U27923 ( .A0(n6882), .A1(AOPA[31]), .B0(n16444), .Y(n3319) );
  OAI21XL U27924 ( .A0(n6886), .A1(AOPA[30]), .B0(n16448), .Y(n3315) );
  OAI21XL U27925 ( .A0(n6886), .A1(AOPA[29]), .B0(n16452), .Y(n3307) );
  OAI21XL U27926 ( .A0(n5913), .A1(AOPA[28]), .B0(n16456), .Y(n3303) );
  OAI21XL U27927 ( .A0(n6882), .A1(AOPA[27]), .B0(n16460), .Y(n3299) );
  OAI21XL U27928 ( .A0(n6882), .A1(AOPA[26]), .B0(n16465), .Y(n3295) );
  OAI21XL U27929 ( .A0(n5915), .A1(AOPA[25]), .B0(n16469), .Y(n3291) );
  OAI21XL U27930 ( .A0(n6882), .A1(AOPA[24]), .B0(n16474), .Y(n3287) );
  OAI21XL U27931 ( .A0(n5913), .A1(AOPA[23]), .B0(n16478), .Y(n3283) );
  OAI21XL U27932 ( .A0(n5913), .A1(AOPA[22]), .B0(n16482), .Y(n3279) );
  OAI21XL U27933 ( .A0(n5906), .A1(AOPA[21]), .B0(n16486), .Y(n3275) );
  OAI21XL U27934 ( .A0(n6883), .A1(AOPA[20]), .B0(n16491), .Y(n3271) );
  OAI21XL U27935 ( .A0(n5913), .A1(AOPA[19]), .B0(n16495), .Y(n3263) );
  OAI21XL U27936 ( .A0(n5906), .A1(AOPA[18]), .B0(n16500), .Y(n3259) );
  OAI21XL U27937 ( .A0(n5905), .A1(AOPA[17]), .B0(n16505), .Y(n3255) );
  OAI21XL U27938 ( .A0(n6886), .A1(AOPA[16]), .B0(n16509), .Y(n3251) );
  OAI21XL U27939 ( .A0(n5908), .A1(AOPA[15]), .B0(n16512), .Y(n3247) );
  OAI21XL U27940 ( .A0(n6886), .A1(AOPA[14]), .B0(n16516), .Y(n3243) );
  OAI21XL U27941 ( .A0(n6886), .A1(AOPA[13]), .B0(n16520), .Y(n3239) );
  OAI21XL U27942 ( .A0(n5800), .A1(AOPA[12]), .B0(n16524), .Y(n3235) );
  OAI21XL U27943 ( .A0(n5913), .A1(AOPA[11]), .B0(n16528), .Y(n3231) );
  OAI21XL U27944 ( .A0(n6881), .A1(AOPA[10]), .B0(n16532), .Y(n3227) );
  OAI21XL U27945 ( .A0(n5905), .A1(AOPA[9]), .B0(n16536), .Y(n3427) );
  OAI21XL U27946 ( .A0(n5909), .A1(AOPA[8]), .B0(n16540), .Y(n3423) );
  OAI21XL U27947 ( .A0(n6882), .A1(AOPA[7]), .B0(n16544), .Y(n3419) );
  OAI21XL U27948 ( .A0(n5907), .A1(AOPA[6]), .B0(n16547), .Y(n3415) );
  OAI21XL U27949 ( .A0(n5912), .A1(AOPA[5]), .B0(n16551), .Y(n3411) );
  OAI21XL U27950 ( .A0(n5912), .A1(AOPA[4]), .B0(n16555), .Y(n3399) );
  OAI21XL U27951 ( .A0(n6883), .A1(AOPA[3]), .B0(n16558), .Y(n3355) );
  OAI21XL U27952 ( .A0(n6880), .A1(AOPA[2]), .B0(n16563), .Y(n3311) );
  OAI21XL U27953 ( .A0(n5912), .A1(AOPA[1]), .B0(n16568), .Y(n3267) );
  AOI21XL U27954 ( .A0(B3_q[0]), .A1(n7127), .B0(n28985), .Y(n16572) );
  OAI21XL U27955 ( .A0(n5913), .A1(AOPA[0]), .B0(n16574), .Y(n3223) );
  NOR2XL U27956 ( .A(U2_U0_y0[2]), .B(U2_U0_y2[2]), .Y(n16575) );
  NOR2XL U27957 ( .A(U2_U0_y0[3]), .B(U2_U0_y2[3]), .Y(n16581) );
  NOR2XL U27958 ( .A(n16575), .B(n16581), .Y(n16584) );
  NOR2XL U27959 ( .A(U2_U0_y0[1]), .B(U2_U0_y2[1]), .Y(n16578) );
  NAND2XL U27960 ( .A(U2_U0_y0[0]), .B(U2_U0_y2[0]), .Y(n16577) );
  NAND2XL U27961 ( .A(U2_U0_y0[1]), .B(U2_U0_y2[1]), .Y(n16576) );
  OAI21XL U27962 ( .A0(n16578), .A1(n16577), .B0(n16576), .Y(n16583) );
  NAND2XL U27963 ( .A(U2_U0_y0[2]), .B(U2_U0_y2[2]), .Y(n16580) );
  NAND2XL U27964 ( .A(U2_U0_y0[3]), .B(U2_U0_y2[3]), .Y(n16579) );
  OAI21XL U27965 ( .A0(n16581), .A1(n16580), .B0(n16579), .Y(n16582) );
  AOI21XL U27966 ( .A0(n16584), .A1(n16583), .B0(n16582), .Y(n16599) );
  NOR2XL U27967 ( .A(U2_U0_y0[4]), .B(U2_U0_y2[4]), .Y(n16585) );
  NOR2XL U27968 ( .A(U2_U0_y0[5]), .B(U2_U0_y2[5]), .Y(n16590) );
  NOR2XL U27969 ( .A(n16585), .B(n16590), .Y(n16587) );
  NOR2XL U27970 ( .A(U2_U0_y0[6]), .B(U2_U0_y2[6]), .Y(n16586) );
  NAND2XL U27971 ( .A(n16587), .B(n16596), .Y(n16598) );
  NAND2XL U27972 ( .A(U2_U0_y0[4]), .B(U2_U0_y2[4]), .Y(n16589) );
  NAND2XL U27973 ( .A(U2_U0_y0[5]), .B(U2_U0_y2[5]), .Y(n16588) );
  OAI21XL U27974 ( .A0(n16590), .A1(n16589), .B0(n16588), .Y(n16595) );
  NAND2XL U27975 ( .A(U2_U0_y0[6]), .B(U2_U0_y2[6]), .Y(n16592) );
  NAND2XL U27976 ( .A(U2_U0_y0[7]), .B(U2_U0_y2[7]), .Y(n16591) );
  OAI21XL U27977 ( .A0(n16593), .A1(n16592), .B0(n16591), .Y(n16594) );
  OAI21XL U27978 ( .A0(n16599), .A1(n16598), .B0(n16597), .Y(n16623) );
  OR2X2 U27979 ( .A(n16616), .B(n16603), .Y(n16619) );
  NAND2XL U27980 ( .A(U2_U0_y0[8]), .B(U2_U0_y2[8]), .Y(n16606) );
  NAND2XL U27981 ( .A(U2_U0_y0[9]), .B(U2_U0_y2[9]), .Y(n16605) );
  OAI21XL U27982 ( .A0(n16607), .A1(n16606), .B0(n16605), .Y(n16612) );
  NAND2XL U27983 ( .A(U2_U0_y0[10]), .B(U2_U0_y2[10]), .Y(n16609) );
  NAND2XL U27984 ( .A(U2_U0_y0[11]), .B(U2_U0_y2[11]), .Y(n16608) );
  OAI21XL U27985 ( .A0(n16610), .A1(n16609), .B0(n16608), .Y(n16611) );
  NAND2XL U27986 ( .A(U2_U0_y0[12]), .B(U2_U0_y2[12]), .Y(n16615) );
  OAI21XL U27987 ( .A0(n16616), .A1(n16615), .B0(n16614), .Y(n16617) );
  OAI21XL U27988 ( .A0(n16620), .A1(n16619), .B0(n16618), .Y(n16621) );
  INVXL U27989 ( .A(n16940), .Y(n16630) );
  NAND2XL U27990 ( .A(n7537), .B(n16636), .Y(n16941) );
  INVXL U27991 ( .A(n16941), .Y(n16637) );
  INVXL U27992 ( .A(n16641), .Y(n16642) );
  INVXL U27993 ( .A(n16643), .Y(n16645) );
  INVXL U27994 ( .A(n16668), .Y(n16676) );
  AOI21XL U27995 ( .A0(n16676), .A1(n16669), .B0(n6675), .Y(n16672) );
  XOR2X1 U27996 ( .A(n16672), .B(n16671), .Y(n16673) );
  NAND2XL U27997 ( .A(n16674), .B(n16967), .Y(n16973) );
  AOI21XL U27998 ( .A0(n16700), .A1(n16681), .B0(n16680), .Y(n16690) );
  OAI21XL U27999 ( .A0(n16690), .A1(n16683), .B0(n16682), .Y(n16686) );
  NAND2XL U28000 ( .A(n8574), .B(n16684), .Y(n16981) );
  NAND2XL U28001 ( .A(n16688), .B(n16979), .Y(n16984) );
  AOI21XL U28002 ( .A0(n16700), .A1(n16693), .B0(n16692), .Y(n16696) );
  NAND2XL U28003 ( .A(n8580), .B(n16694), .Y(n16989) );
  OAI21XL U28004 ( .A0(n16734), .A1(n16704), .B0(n16703), .Y(n16714) );
  OAI21XL U28005 ( .A0(n16734), .A1(n16717), .B0(n16716), .Y(n16730) );
  INVXL U28006 ( .A(n16718), .Y(n16721) );
  INVXL U28007 ( .A(n6583), .Y(n16749) );
  OAI21XL U28008 ( .A0(n16768), .A1(n16759), .B0(n16758), .Y(n16764) );
  XOR2XL U28009 ( .A(n16774), .B(n16773), .Y(n16775) );
  XOR2XL U28010 ( .A(n16778), .B(n16777), .Y(n16779) );
  CLKINVX3 U28011 ( .A(n17032), .Y(n25267) );
  XNOR2XL U28012 ( .A(n16780), .B(U1_A_i_d0[0]), .Y(n17049) );
  NAND2XL U28013 ( .A(n16783), .B(n16782), .Y(n16784) );
  MXI2X1 U28014 ( .A(U1_pipe7[25]), .B(n16786), .S0(n5812), .Y(n4978) );
  INVXL U28015 ( .A(n16789), .Y(n16791) );
  INVXL U28016 ( .A(n17055), .Y(n16792) );
  INVXL U28017 ( .A(n16794), .Y(n16795) );
  INVX1 U28018 ( .A(n17065), .Y(n16803) );
  AOI21XL U28019 ( .A0(n16821), .A1(n16813), .B0(n16812), .Y(n16816) );
  XOR2X1 U28020 ( .A(n16816), .B(n16815), .Y(n16817) );
  MXI2X1 U28021 ( .A(U1_pipe7[20]), .B(n16817), .S0(n25330), .Y(n4973) );
  AOI21XL U28022 ( .A0(n16832), .A1(n14949), .B0(n16824), .Y(n16828) );
  NAND2XL U28023 ( .A(n16830), .B(n17074), .Y(n17080) );
  OAI21XL U28024 ( .A0(n16845), .A1(n16836), .B0(n16842), .Y(n16840) );
  AOI21XL U28025 ( .A0(n16855), .A1(n14947), .B0(n16847), .Y(n16851) );
  NAND2XL U28026 ( .A(n14947), .B(n16853), .Y(n16854) );
  XNOR2X1 U28027 ( .A(n16855), .B(n16854), .Y(n16856) );
  OAI21XL U28028 ( .A0(n16887), .A1(n16859), .B0(n16858), .Y(n16867) );
  AOI21XL U28029 ( .A0(n16867), .A1(n16860), .B0(n6952), .Y(n16863) );
  INVXL U28030 ( .A(n16875), .Y(n16877) );
  NAND2XL U28031 ( .A(n16885), .B(n17117), .Y(n17128) );
  AOI21XL U28032 ( .A0(n16907), .A1(n16891), .B0(n16890), .Y(n16894) );
  OAI21XL U28033 ( .A0(n16920), .A1(n16911), .B0(n16910), .Y(n16916) );
  XOR2XL U28034 ( .A(n16926), .B(n16925), .Y(n16927) );
  XOR2XL U28035 ( .A(n16930), .B(n16929), .Y(n16931) );
  XNOR2XL U28036 ( .A(n20180), .B(n16932), .Y(n17166) );
  NAND2XL U28037 ( .A(U1_pipe7[0]), .B(U1_pipe6[0]), .Y(n16934) );
  OAI21XL U28038 ( .A0(n16935), .A1(n16934), .B0(n16933), .Y(n17802) );
  OAI21XL U28039 ( .A0(n7535), .A1(n16946), .B0(n16945), .Y(n16948) );
  XNOR2XL U28040 ( .A(n16948), .B(n16947), .Y(n16949) );
  OAI21XL U28041 ( .A0(n7535), .A1(n16951), .B0(n16950), .Y(n16953) );
  XNOR2XL U28042 ( .A(n16953), .B(n16952), .Y(n16954) );
  XOR2X1 U28043 ( .A(n7535), .B(n16955), .Y(n16956) );
  OAI21XL U28044 ( .A0(n16969), .A1(n16968), .B0(n16967), .Y(n16971) );
  XNOR2XL U28045 ( .A(n16971), .B(n16970), .Y(n16972) );
  INVXL U28046 ( .A(n16975), .Y(n16978) );
  INVXL U28047 ( .A(n16976), .Y(n16977) );
  OAI21XL U28048 ( .A0(n16985), .A1(n16980), .B0(n16979), .Y(n16982) );
  XNOR2XL U28049 ( .A(n16982), .B(n16981), .Y(n16983) );
  OAI21XL U28050 ( .A0(n17016), .A1(n16996), .B0(n16995), .Y(n17002) );
  AOI21XL U28051 ( .A0(n17002), .A1(n8553), .B0(n16997), .Y(n16999) );
  OAI21XL U28052 ( .A0(n17016), .A1(n17005), .B0(n17004), .Y(n17013) );
  INVXL U28053 ( .A(n17018), .Y(n17031) );
  AOI21XL U28054 ( .A0(n17031), .A1(n17020), .B0(n17019), .Y(n17022) );
  OAI21XL U28055 ( .A0(n17041), .A1(n17036), .B0(n17035), .Y(n17038) );
  XOR2XL U28056 ( .A(n17044), .B(n17043), .Y(n17045) );
  XNOR2XL U28057 ( .A(n17047), .B(n17046), .Y(n17048) );
  NAND2XL U28058 ( .A(n13987), .B(n17051), .Y(n17052) );
  XNOR2X1 U28059 ( .A(n17053), .B(n17052), .Y(n17054) );
  MXI2X1 U28060 ( .A(U1_pipe5[25]), .B(n17054), .S0(n5804), .Y(n4922) );
  XOR2X1 U28061 ( .A(n17056), .B(n17055), .Y(n17057) );
  OAI21XL U28062 ( .A0(n17069), .A1(n17059), .B0(n17058), .Y(n17061) );
  MXI2X1 U28063 ( .A(U1_pipe5[23]), .B(n17062), .S0(n20025), .Y(n4920) );
  OAI21XL U28064 ( .A0(n17069), .A1(n17064), .B0(n17063), .Y(n17066) );
  XNOR2X1 U28065 ( .A(n17066), .B(n17065), .Y(n17067) );
  MXI2X1 U28066 ( .A(U1_pipe5[22]), .B(n17067), .S0(n24784), .Y(n4919) );
  OAI21XL U28067 ( .A0(n17076), .A1(n17075), .B0(n17074), .Y(n17078) );
  XNOR2X1 U28068 ( .A(n17078), .B(n17077), .Y(n17079) );
  MXI2X1 U28069 ( .A(U1_pipe5[18]), .B(n17079), .S0(n17187), .Y(n4915) );
  OAI21XL U28070 ( .A0(n17095), .A1(n17087), .B0(n17092), .Y(n17090) );
  NAND2XL U28071 ( .A(n6941), .B(n17088), .Y(n17089) );
  NAND2XL U28072 ( .A(n17093), .B(n17092), .Y(n17094) );
  AOI21XL U28073 ( .A0(n5966), .A1(n17104), .B0(n17097), .Y(n17101) );
  NAND2XL U28074 ( .A(n17104), .B(n17103), .Y(n17105) );
  OAI21XL U28075 ( .A0(n17129), .A1(n17109), .B0(n17108), .Y(n17115) );
  OAI21XL U28076 ( .A0(n17129), .A1(n17118), .B0(n17117), .Y(n17126) );
  INVXL U28077 ( .A(n17119), .Y(n17120) );
  AOI21XL U28078 ( .A0(n17149), .A1(n17133), .B0(n17132), .Y(n17136) );
  INVXL U28079 ( .A(n17140), .Y(n17142) );
  OAI21XL U28080 ( .A0(n17158), .A1(n17153), .B0(n17152), .Y(n17155) );
  XOR2XL U28081 ( .A(n17161), .B(n17160), .Y(n17162) );
  XNOR2XL U28082 ( .A(n17164), .B(n17163), .Y(n17165) );
  NAND2XL U28083 ( .A(U1_pipe5[0]), .B(U1_pipe4[0]), .Y(n17168) );
  OAI21XL U28084 ( .A0(n17169), .A1(n17168), .B0(n17167), .Y(n17813) );
  NAND2XL U28085 ( .A(n17178), .B(n17177), .Y(n17458) );
  INVXL U28086 ( .A(n17183), .Y(n17185) );
  XNOR2X1 U28087 ( .A(n17186), .B(n17465), .Y(n17188) );
  MXI2X1 U28088 ( .A(U1_pipe14[23]), .B(n17188), .S0(n17187), .Y(n4774) );
  XNOR2X1 U28089 ( .A(n17192), .B(n17471), .Y(n17193) );
  MXI2X1 U28090 ( .A(U1_pipe14[22]), .B(n17193), .S0(n5809), .Y(n4773) );
  NAND2XL U28091 ( .A(n17195), .B(n17194), .Y(n17475) );
  NAND2XL U28092 ( .A(n17199), .B(n17198), .Y(n17487) );
  OAI21XL U28093 ( .A0(n17203), .A1(n17202), .B0(n17207), .Y(n17205) );
  NAND2XL U28094 ( .A(n7001), .B(n17204), .Y(n17494) );
  XNOR2XL U28095 ( .A(n17205), .B(n17494), .Y(n17206) );
  NAND2XL U28096 ( .A(n17208), .B(n17207), .Y(n17498) );
  INVXL U28097 ( .A(n17211), .Y(n17214) );
  INVXL U28098 ( .A(n17212), .Y(n17213) );
  XNOR2XL U28099 ( .A(n17218), .B(n17508), .Y(n17219) );
  NAND2XL U28100 ( .A(n17229), .B(n17228), .Y(n17522) );
  AOI21XL U28101 ( .A0(n17240), .A1(n9577), .B0(n17235), .Y(n17237) );
  NAND2XL U28102 ( .A(n9577), .B(n17239), .Y(n17535) );
  INVXL U28103 ( .A(n17251), .Y(n17244) );
  NAND2XL U28104 ( .A(n17247), .B(n17246), .Y(n17545) );
  INVXL U28105 ( .A(n17259), .Y(n17275) );
  AOI21XL U28106 ( .A0(n17275), .A1(n17261), .B0(n17260), .Y(n17264) );
  INVXL U28107 ( .A(n17268), .Y(n17270) );
  OAI21XL U28108 ( .A0(n17286), .A1(n17283), .B0(n17284), .Y(n17281) );
  INVXL U28109 ( .A(n17278), .Y(n17280) );
  XOR2XL U28110 ( .A(n17587), .B(n17291), .Y(n17292) );
  XNOR2XL U28111 ( .A(n17591), .B(n17294), .Y(n17295) );
  XNOR2XL U28112 ( .A(n19231), .B(U1_A_i_d0[0]), .Y(n17595) );
  MXI2X1 U28113 ( .A(U1_pipe15[25]), .B(n17298), .S0(n5809), .Y(n4804) );
  INVX1 U28114 ( .A(n17299), .Y(n17301) );
  NAND2X1 U28115 ( .A(n17301), .B(n17300), .Y(n17605) );
  XOR2X1 U28116 ( .A(n17302), .B(n17605), .Y(n17303) );
  MXI2X1 U28117 ( .A(U1_pipe15[24]), .B(n17303), .S0(n25267), .Y(n4803) );
  INVXL U28118 ( .A(n17307), .Y(n17309) );
  MXI2X1 U28119 ( .A(U1_pipe15[23]), .B(n17311), .S0(n25267), .Y(n4802) );
  OAI21XL U28120 ( .A0(n17320), .A1(n17312), .B0(n17317), .Y(n17315) );
  XNOR2X1 U28121 ( .A(n17315), .B(n17617), .Y(n17316) );
  MXI2X1 U28122 ( .A(U1_pipe15[22]), .B(n17316), .S0(n25267), .Y(n4801) );
  NAND2XL U28123 ( .A(n17318), .B(n17317), .Y(n17319) );
  XOR2X1 U28124 ( .A(n17320), .B(n17319), .Y(n17321) );
  INVXL U28125 ( .A(n17324), .Y(n17327) );
  INVXL U28126 ( .A(n17325), .Y(n17326) );
  MXI2X1 U28127 ( .A(U1_pipe15[20]), .B(n17333), .S0(n25267), .Y(n4799) );
  NAND2XL U28128 ( .A(n17335), .B(n17334), .Y(n17336) );
  OAI21XL U28129 ( .A0(n17339), .A1(n17338), .B0(n17344), .Y(n17342) );
  XNOR2X1 U28130 ( .A(n17342), .B(n17634), .Y(n17343) );
  MXI2X1 U28131 ( .A(U1_pipe15[18]), .B(n17343), .S0(n25267), .Y(n4797) );
  NAND2XL U28132 ( .A(n17345), .B(n17344), .Y(n17346) );
  XNOR2X1 U28133 ( .A(n17347), .B(n17346), .Y(n17348) );
  INVXL U28134 ( .A(n17349), .Y(n17352) );
  INVXL U28135 ( .A(n17350), .Y(n17351) );
  OAI21XL U28136 ( .A0(n17360), .A1(n17353), .B0(n17358), .Y(n17356) );
  XNOR2X1 U28137 ( .A(n17356), .B(n17649), .Y(n17357) );
  MXI2X1 U28138 ( .A(U1_pipe15[16]), .B(n17357), .S0(n25267), .Y(n4795) );
  AOI21XL U28139 ( .A0(n17370), .A1(n13554), .B0(n17362), .Y(n17366) );
  NAND2XL U28140 ( .A(n13554), .B(n17368), .Y(n17369) );
  XNOR2X1 U28141 ( .A(n17370), .B(n17369), .Y(n17371) );
  MXI2X1 U28142 ( .A(U1_pipe15[13]), .B(n17371), .S0(n22853), .Y(n4792) );
  OAI21XL U28143 ( .A0(n17401), .A1(n17374), .B0(n17373), .Y(n17383) );
  AOI21XL U28144 ( .A0(n17383), .A1(n13545), .B0(n17375), .Y(n17379) );
  NAND2XL U28145 ( .A(n13545), .B(n17381), .Y(n17382) );
  OAI21XL U28146 ( .A0(n17401), .A1(n17385), .B0(n17399), .Y(n17397) );
  INVXL U28147 ( .A(n17386), .Y(n17395) );
  INVXL U28148 ( .A(n17394), .Y(n17387) );
  NAND2XL U28149 ( .A(n17395), .B(n17394), .Y(n17396) );
  NAND2XL U28150 ( .A(n17400), .B(n17399), .Y(n17695) );
  AOI21XL U28151 ( .A0(n17421), .A1(n17405), .B0(n17404), .Y(n17408) );
  INVXL U28152 ( .A(n17412), .Y(n17414) );
  OAI21XL U28153 ( .A0(n17434), .A1(n17430), .B0(n17431), .Y(n17428) );
  OAI21XL U28154 ( .A0(n17443), .A1(n17436), .B0(n17441), .Y(n17439) );
  XOR2XL U28155 ( .A(n17444), .B(n17443), .Y(n17445) );
  XNOR2XL U28156 ( .A(n17446), .B(n19507), .Y(n17742) );
  INVXL U28157 ( .A(n17458), .Y(n17459) );
  INVXL U28158 ( .A(n17461), .Y(n17464) );
  MXI2X1 U28159 ( .A(U1_pipe10[23]), .B(n17468), .S0(n17641), .Y(n4861) );
  MXI2X1 U28160 ( .A(U1_pipe10[22]), .B(n17474), .S0(n17641), .Y(n4860) );
  AOI21XL U28161 ( .A0(n17489), .A1(n17482), .B0(n17481), .Y(n17485) );
  XOR2X1 U28162 ( .A(n17485), .B(n17484), .Y(n17486) );
  INVXL U28163 ( .A(n17487), .Y(n17488) );
  AOI21XL U28164 ( .A0(n17500), .A1(n17493), .B0(n17492), .Y(n17496) );
  INVXL U28165 ( .A(n17503), .Y(n17504) );
  AOI21XL U28166 ( .A0(n17524), .A1(n17517), .B0(n17516), .Y(n17520) );
  OAI21XL U28167 ( .A0(n17555), .A1(n17528), .B0(n17527), .Y(n17537) );
  OAI21XL U28168 ( .A0(n17555), .A1(n17540), .B0(n17539), .Y(n17551) );
  INVXL U28169 ( .A(n17541), .Y(n17544) );
  INVXL U28170 ( .A(n17542), .Y(n17543) );
  AOI21XL U28171 ( .A0(n17574), .A1(n17559), .B0(n17558), .Y(n17562) );
  OAI21XL U28172 ( .A0(n17585), .A1(n17578), .B0(n17577), .Y(n17581) );
  XOR2XL U28173 ( .A(n17589), .B(n17588), .Y(n17590) );
  XOR2XL U28174 ( .A(n17593), .B(n17592), .Y(n17594) );
  INVXL U28175 ( .A(n17596), .Y(n17598) );
  NAND2XL U28176 ( .A(n17598), .B(n17597), .Y(n17599) );
  XOR2X1 U28177 ( .A(n17600), .B(n17599), .Y(n17601) );
  MXI2X1 U28178 ( .A(U1_pipe11[25]), .B(n17601), .S0(n25330), .Y(n4891) );
  OAI21XL U28179 ( .A0(n17625), .A1(n17604), .B0(n17603), .Y(n17607) );
  XNOR2X1 U28180 ( .A(n17607), .B(n17606), .Y(n17608) );
  MXI2X1 U28181 ( .A(U1_pipe11[24]), .B(n17608), .S0(n5812), .Y(n4890) );
  INVXL U28182 ( .A(n17609), .Y(n17612) );
  OAI21XL U28183 ( .A0(n17625), .A1(n17612), .B0(n17611), .Y(n17615) );
  XNOR2X1 U28184 ( .A(n17615), .B(n17614), .Y(n17616) );
  MXI2X1 U28185 ( .A(U1_pipe11[23]), .B(n17616), .S0(n25330), .Y(n4889) );
  OAI21XL U28186 ( .A0(n17625), .A1(n17621), .B0(n17622), .Y(n17619) );
  XNOR2X1 U28187 ( .A(n17619), .B(n17618), .Y(n17620) );
  MXI2X1 U28188 ( .A(U1_pipe11[22]), .B(n17620), .S0(n25330), .Y(n4888) );
  INVXL U28189 ( .A(n17621), .Y(n17623) );
  XOR2X1 U28190 ( .A(n17625), .B(n17624), .Y(n17626) );
  NAND2XL U28191 ( .A(n17628), .B(n17627), .Y(n17629) );
  MXI2X1 U28192 ( .A(U1_pipe11[19]), .B(n17631), .S0(n20438), .Y(n4885) );
  MXI2X1 U28193 ( .A(U1_pipe11[18]), .B(n17637), .S0(n5812), .Y(n4884) );
  INVXL U28194 ( .A(n17643), .Y(n17646) );
  INVXL U28195 ( .A(n17644), .Y(n17645) );
  OAI21XL U28196 ( .A0(n17655), .A1(n17648), .B0(n17647), .Y(n17651) );
  XNOR2X1 U28197 ( .A(n17651), .B(n17650), .Y(n17652) );
  MXI2X1 U28198 ( .A(U1_pipe11[16]), .B(n17652), .S0(n20438), .Y(n4882) );
  AOI21XL U28199 ( .A0(n17664), .A1(n13034), .B0(n17657), .Y(n17660) );
  NAND2XL U28200 ( .A(n13025), .B(n17658), .Y(n17659) );
  XNOR2X1 U28201 ( .A(n17664), .B(n17663), .Y(n17665) );
  OAI21XL U28202 ( .A0(n17697), .A1(n17668), .B0(n17667), .Y(n17678) );
  AOI21XL U28203 ( .A0(n17678), .A1(n17676), .B0(n17669), .Y(n17673) );
  INVXL U28204 ( .A(n17690), .Y(n17683) );
  INVXL U28205 ( .A(n17684), .Y(n17686) );
  OAI21XL U28206 ( .A0(n17730), .A1(n17726), .B0(n17727), .Y(n17724) );
  INVXL U28207 ( .A(n17720), .Y(n17722) );
  XOR2XL U28208 ( .A(n17736), .B(n17735), .Y(n17737) );
  XOR2XL U28209 ( .A(n17740), .B(n17739), .Y(n17741) );
  NAND2XL U28210 ( .A(U1_pipe11[0]), .B(U1_pipe10[0]), .Y(n17744) );
  OAI21XL U28211 ( .A0(n17745), .A1(n17744), .B0(n17743), .Y(n17831) );
  OAI21XL U28212 ( .A0(n21732), .A1(n17751), .B0(n17750), .Y(n17843) );
  INVXL U28213 ( .A(n23177), .Y(n17790) );
  CMPR22X1 U28214 ( .A(U2_U0_y2[14]), .B(U2_U0_y0[14]), .CO(n23176), .S(n23132) );
  OR2X2 U28215 ( .A(n17753), .B(n17752), .Y(n17788) );
  NOR2XL U28216 ( .A(n17754), .B(U2_A_i_d[1]), .Y(n17837) );
  OAI21XL U28217 ( .A0(n17758), .A1(n17797), .B0(n17799), .Y(n17763) );
  CMPR22X1 U28218 ( .A(U1_pipe7[2]), .B(U1_pipe6[2]), .CO(n17760), .S(n16936)
         );
  OAI21XL U28219 ( .A0(n17765), .A1(n17808), .B0(n17810), .Y(n17770) );
  CMPR22X1 U28220 ( .A(U1_pipe5[2]), .B(U1_pipe4[2]), .CO(n17767), .S(n17170)
         );
  OAI21XL U28221 ( .A0(n17774), .A1(n17773), .B0(n17772), .Y(n17871) );
  CMPR22X1 U28222 ( .A(U1_pipe14[2]), .B(n28744), .CO(n17776), .S(n17447) );
  OAI21XL U28223 ( .A0(n17780), .A1(n17826), .B0(n17828), .Y(n17785) );
  CMPR22X1 U28224 ( .A(U1_pipe11[2]), .B(U1_pipe10[2]), .CO(n17782), .S(n17746) );
  OAI21XL U28225 ( .A0(n17787), .A1(n17837), .B0(n17839), .Y(n17795) );
  CMPR32X1 U28226 ( .A(n17790), .B(n17789), .C(n17788), .CO(n17791), .S(n17754) );
  OAI21XL U28227 ( .A0(n17800), .A1(n17799), .B0(n17798), .Y(n17801) );
  CMPR22X1 U28228 ( .A(U1_pipe7[3]), .B(U1_pipe6[3]), .CO(n17805), .S(n17759)
         );
  OAI21XL U28229 ( .A0(n17811), .A1(n17810), .B0(n17809), .Y(n17812) );
  CMPR22X1 U28230 ( .A(U1_pipe5[3]), .B(U1_pipe4[3]), .CO(n17816), .S(n17766)
         );
  OAI21XL U28231 ( .A0(n17819), .A1(n17866), .B0(n17868), .Y(n17824) );
  CMPR22X1 U28232 ( .A(U1_pipe14[3]), .B(n28743), .CO(n17821), .S(n17775) );
  OAI21XL U28233 ( .A0(n17829), .A1(n17828), .B0(n17827), .Y(n17830) );
  CMPR22X1 U28234 ( .A(U1_pipe11[3]), .B(U1_pipe10[3]), .CO(n17834), .S(n17781) );
  NOR2XL U28235 ( .A(n17840), .B(n17837), .Y(n17842) );
  OAI21XL U28236 ( .A0(n17840), .A1(n17839), .B0(n17838), .Y(n17841) );
  AOI21XL U28237 ( .A0(n17843), .A1(n17842), .B0(n17841), .Y(n18050) );
  INVXL U28238 ( .A(n23276), .Y(n17888) );
  CMPR22X1 U28239 ( .A(U2_U0_y2[16]), .B(U2_U0_y0[16]), .CO(n23275), .S(n23225) );
  CMPR32X1 U28240 ( .A(n17845), .B(n17844), .C(U2_A_i_d[2]), .CO(n17846), .S(
        n17792) );
  NOR2XL U28241 ( .A(n17847), .B(n17846), .Y(n17933) );
  NAND2XL U28242 ( .A(n17847), .B(n17846), .Y(n17935) );
  CMPR22X1 U28243 ( .A(U1_pipe7[4]), .B(U1_pipe6[4]), .CO(n17853), .S(n17804)
         );
  CMPR22X1 U28244 ( .A(U1_pipe5[4]), .B(U1_pipe4[4]), .CO(n17861), .S(n17815)
         );
  NAND2XL U28245 ( .A(n17862), .B(n17906), .Y(n17863) );
  OAI21XL U28246 ( .A0(n17869), .A1(n17868), .B0(n17867), .Y(n17870) );
  CMPR22X1 U28247 ( .A(U1_pipe14[4]), .B(n28887), .CO(n17874), .S(n17820) );
  CMPR22X1 U28248 ( .A(U1_pipe11[4]), .B(U1_pipe10[4]), .CO(n17880), .S(n17833) );
  CMPR22X1 U28249 ( .A(U2_U0_y2[17]), .B(U2_U0_y0[17]), .CO(n23321), .S(n23276) );
  INVXL U28250 ( .A(n23321), .Y(n17938) );
  CMPR32X1 U28251 ( .A(n17888), .B(n17887), .C(U2_A_i_d[3]), .CO(n17889), .S(
        n17847) );
  NAND2XL U28252 ( .A(n17890), .B(n17889), .Y(n17934) );
  OAI21XL U28253 ( .A0(n17898), .A1(n17897), .B0(n17896), .Y(n18030) );
  CMPR22X1 U28254 ( .A(U1_pipe11[5]), .B(U1_pipe10[5]), .CO(n17901), .S(n17879) );
  OAI21XL U28255 ( .A0(n17908), .A1(n17907), .B0(n17906), .Y(n18007) );
  CMPR22X1 U28256 ( .A(U1_pipe5[5]), .B(U1_pipe4[5]), .CO(n17911), .S(n17860)
         );
  CMPR22X1 U28257 ( .A(U1_pipe14[5]), .B(n28886), .CO(n17918), .S(n17873) );
  OAI21XL U28258 ( .A0(n17926), .A1(n17925), .B0(n17924), .Y(n17991) );
  CMPR22X1 U28259 ( .A(U1_pipe7[5]), .B(U1_pipe6[5]), .CO(n17929), .S(n17852)
         );
  NOR2XL U28260 ( .A(n17933), .B(n17936), .Y(n18041) );
  OAI21XL U28261 ( .A0(n17936), .A1(n17935), .B0(n17934), .Y(n18046) );
  INVXL U28262 ( .A(n23366), .Y(n17978) );
  CMPR32X1 U28263 ( .A(n17939), .B(n17938), .C(U2_A_i_d[4]), .CO(n17940), .S(
        n17890) );
  INVXL U28264 ( .A(n18040), .Y(n17942) );
  OAI21XL U28265 ( .A0(n17945), .A1(n17985), .B0(n17988), .Y(n17950) );
  CMPR22X1 U28266 ( .A(U1_pipe7[6]), .B(U1_pipe6[6]), .CO(n17947), .S(n17928)
         );
  OAI21XL U28267 ( .A0(n17952), .A1(n18001), .B0(n18004), .Y(n17957) );
  CMPR22X1 U28268 ( .A(U1_pipe5[6]), .B(U1_pipe4[6]), .CO(n17954), .S(n17910)
         );
  OAI21XL U28269 ( .A0(n17962), .A1(n17961), .B0(n17960), .Y(n18076) );
  CMPR22X1 U28270 ( .A(U1_pipe14[6]), .B(n28742), .CO(n17965), .S(n17917) );
  OAI21XL U28271 ( .A0(n17969), .A1(n18024), .B0(n18027), .Y(n17974) );
  CMPR22X1 U28272 ( .A(U1_pipe11[6]), .B(U1_pipe10[6]), .CO(n17971), .S(n17900) );
  OAI21XL U28273 ( .A0(n17976), .A1(n18040), .B0(n18043), .Y(n17983) );
  INVXL U28274 ( .A(n23428), .Y(n18051) );
  INVXL U28275 ( .A(n18044), .Y(n17981) );
  NAND2XL U28276 ( .A(n17980), .B(n17979), .Y(n18042) );
  OAI21XL U28277 ( .A0(n17989), .A1(n17988), .B0(n17987), .Y(n17990) );
  OAI21XL U28278 ( .A0(n17995), .A1(n17994), .B0(n17993), .Y(n18438) );
  CMPR22X1 U28279 ( .A(U1_pipe7[7]), .B(U1_pipe6[7]), .CO(n17997), .S(n17946)
         );
  OAI21XL U28280 ( .A0(n18005), .A1(n18004), .B0(n18003), .Y(n18006) );
  OAI21XL U28281 ( .A0(n18011), .A1(n18010), .B0(n18009), .Y(n18457) );
  CMPR22X1 U28282 ( .A(U1_pipe5[7]), .B(U1_pipe4[7]), .CO(n18013), .S(n17953)
         );
  OAI21XL U28283 ( .A0(n18017), .A1(n18070), .B0(n18073), .Y(n18022) );
  CMPR22X1 U28284 ( .A(U1_pipe14[7]), .B(n28885), .CO(n18019), .S(n17964) );
  OAI21XL U28285 ( .A0(n18028), .A1(n18027), .B0(n18026), .Y(n18029) );
  OAI21XL U28286 ( .A0(n18034), .A1(n18033), .B0(n18032), .Y(n18476) );
  CMPR22X1 U28287 ( .A(U1_pipe11[7]), .B(U1_pipe10[7]), .CO(n18036), .S(n17970) );
  OAI21XL U28288 ( .A0(n18044), .A1(n18043), .B0(n18042), .Y(n18045) );
  AOI21X1 U28289 ( .A0(n18047), .A1(n18046), .B0(n18045), .Y(n18048) );
  OAI21XL U28290 ( .A0(n18050), .A1(n18049), .B0(n18048), .Y(n18495) );
  INVXL U28291 ( .A(n23482), .Y(n18093) );
  CMPR22X1 U28292 ( .A(U2_U0_y2[20]), .B(U2_U0_y0[20]), .CO(n23481), .S(n23429) );
  CMPR32X1 U28293 ( .A(n18052), .B(n18051), .C(U2_A_i_d[6]), .CO(n18053), .S(
        n17980) );
  INVXL U28294 ( .A(n18136), .Y(n18055) );
  OAI21XL U28295 ( .A0(n18204), .A1(n18126), .B0(n18128), .Y(n18062) );
  CMPR22X1 U28296 ( .A(U1_pipe11[8]), .B(U1_pipe10[8]), .CO(n18059), .S(n18035) );
  OAI21XL U28297 ( .A0(n18217), .A1(n18110), .B0(n18112), .Y(n18068) );
  CMPR22X1 U28298 ( .A(U1_pipe5[8]), .B(U1_pipe4[8]), .CO(n18065), .S(n18012)
         );
  OAI21XL U28299 ( .A0(n18074), .A1(n18073), .B0(n18072), .Y(n18075) );
  OAI21XL U28300 ( .A0(n18080), .A1(n18079), .B0(n18078), .Y(n18514) );
  CMPR22X1 U28301 ( .A(U1_pipe14[8]), .B(n28884), .CO(n18082), .S(n18018) );
  OAI21XL U28302 ( .A0(n18239), .A1(n18100), .B0(n18102), .Y(n18090) );
  CMPR22X1 U28303 ( .A(U1_pipe7[8]), .B(U1_pipe6[8]), .CO(n18087), .S(n17996)
         );
  NAND2XL U28304 ( .A(n18088), .B(n18101), .Y(n18089) );
  OAI21XL U28305 ( .A0(n18252), .A1(n18136), .B0(n18138), .Y(n18098) );
  INVX1 U28306 ( .A(n23524), .Y(n18142) );
  ADDFHX1 U28307 ( .A(n18093), .B(n18092), .CI(U2_A_i_d[7]), .CO(n18094), .S(
        n18054) );
  NOR2X1 U28308 ( .A(n18095), .B(n18094), .Y(n18139) );
  NAND2XL U28309 ( .A(n18095), .B(n18094), .Y(n18137) );
  OAI21XL U28310 ( .A0(n18103), .A1(n18102), .B0(n18101), .Y(n18237) );
  OAI21XL U28311 ( .A0(n18239), .A1(n18105), .B0(n18104), .Y(n18150) );
  CMPR22X1 U28312 ( .A(U1_pipe7[9]), .B(U1_pipe6[9]), .CO(n18107), .S(n18086)
         );
  OAI21XL U28313 ( .A0(n18113), .A1(n18112), .B0(n18111), .Y(n18215) );
  OAI21XL U28314 ( .A0(n18217), .A1(n18115), .B0(n18114), .Y(n18159) );
  CMPR22X1 U28315 ( .A(U1_pipe5[9]), .B(U1_pipe4[9]), .CO(n18117), .S(n18064)
         );
  OAI21XL U28316 ( .A0(n18267), .A1(n18166), .B0(n18168), .Y(n18124) );
  CMPR22X1 U28317 ( .A(U1_pipe14[9]), .B(n28741), .CO(n18121), .S(n18081) );
  OAI21XL U28318 ( .A0(n18129), .A1(n18128), .B0(n18127), .Y(n18202) );
  OAI21XL U28319 ( .A0(n18204), .A1(n18131), .B0(n18130), .Y(n18178) );
  CMPR22X1 U28320 ( .A(U1_pipe11[9]), .B(U1_pipe10[9]), .CO(n18133), .S(n18058) );
  NAND2XL U28321 ( .A(n18177), .B(n18199), .Y(n18134) );
  NOR2XL U28322 ( .A(n18136), .B(n18139), .Y(n18245) );
  INVXL U28323 ( .A(n18245), .Y(n18141) );
  OAI21XL U28324 ( .A0(n18252), .A1(n18141), .B0(n18140), .Y(n18187) );
  CMPR32X1 U28325 ( .A(n18143), .B(n18142), .C(U2_A_i_d[8]), .CO(n18144), .S(
        n18095) );
  NOR2XL U28326 ( .A(n18145), .B(n18144), .Y(n18244) );
  INVXL U28327 ( .A(n18244), .Y(n18186) );
  NAND2XL U28328 ( .A(n18145), .B(n18144), .Y(n18247) );
  NAND2XL U28329 ( .A(n18186), .B(n18247), .Y(n18146) );
  CMPR22X1 U28330 ( .A(U1_pipe7[10]), .B(U1_pipe6[10]), .CO(n18152), .S(n18106) );
  CMPR22X1 U28331 ( .A(U1_pipe5[10]), .B(U1_pipe4[10]), .CO(n18161), .S(n18116) );
  OAI21XL U28332 ( .A0(n18169), .A1(n18168), .B0(n18167), .Y(n18265) );
  OAI21XL U28333 ( .A0(n18267), .A1(n18171), .B0(n18170), .Y(n18224) );
  CMPR22X1 U28334 ( .A(U1_pipe14[10]), .B(n28883), .CO(n18173), .S(n18120) );
  CMPR22X1 U28335 ( .A(U1_pipe11[10]), .B(U1_pipe10[10]), .CO(n18180), .S(
        n18132) );
  CLKINVX3 U28336 ( .A(n28997), .Y(n18351) );
  INVXL U28337 ( .A(n18247), .Y(n18185) );
  AOI21XL U28338 ( .A0(n18187), .A1(n18186), .B0(n18185), .Y(n18194) );
  INVX1 U28339 ( .A(n23633), .Y(n18253) );
  NAND2XL U28340 ( .A(n18191), .B(n18190), .Y(n18246) );
  OAI21XL U28341 ( .A0(n18200), .A1(n18199), .B0(n18198), .Y(n18201) );
  OAI21XL U28342 ( .A0(n18204), .A1(n18464), .B0(n18473), .Y(n18292) );
  CMPR22X1 U28343 ( .A(U1_pipe11[11]), .B(U1_pipe10[11]), .CO(n18206), .S(
        n18179) );
  OAI21XL U28344 ( .A0(n18213), .A1(n18212), .B0(n18211), .Y(n18214) );
  OAI21XL U28345 ( .A0(n18217), .A1(n18445), .B0(n18454), .Y(n18283) );
  CMPR22X1 U28346 ( .A(U1_pipe5[11]), .B(U1_pipe4[11]), .CO(n18219), .S(n18160) );
  CMPR22X1 U28347 ( .A(U1_pipe14[11]), .B(n28882), .CO(n18226), .S(n18172) );
  OAI21XL U28348 ( .A0(n18235), .A1(n18234), .B0(n18233), .Y(n18236) );
  OAI21XL U28349 ( .A0(n18239), .A1(n18426), .B0(n18435), .Y(n18274) );
  CMPR22X1 U28350 ( .A(U1_pipe7[11]), .B(U1_pipe6[11]), .CO(n18241), .S(n18151) );
  NOR2XL U28351 ( .A(n18244), .B(n18248), .Y(n18251) );
  NAND2XL U28352 ( .A(n18245), .B(n18251), .Y(n18483) );
  OAI21XL U28353 ( .A0(n18248), .A1(n18247), .B0(n18246), .Y(n18249) );
  INVX1 U28354 ( .A(n23691), .Y(n18303) );
  NOR2XL U28355 ( .A(n18256), .B(n18255), .Y(n18353) );
  INVXL U28356 ( .A(n18353), .Y(n18300) );
  NAND2XL U28357 ( .A(n18300), .B(n18355), .Y(n18257) );
  OAI21XL U28358 ( .A0(n18263), .A1(n18262), .B0(n18261), .Y(n18264) );
  OAI21XL U28359 ( .A0(n18267), .A1(n18502), .B0(n18511), .Y(n18312) );
  CMPR22X1 U28360 ( .A(U1_pipe14[12]), .B(n28881), .CO(n18269), .S(n18225) );
  CMPR22X1 U28361 ( .A(U1_pipe7[12]), .B(U1_pipe6[12]), .CO(n18276), .S(n18240) );
  CMPR22X1 U28362 ( .A(U1_pipe5[12]), .B(U1_pipe4[12]), .CO(n18285), .S(n18218) );
  CMPR22X1 U28363 ( .A(U1_pipe11[12]), .B(U1_pipe10[12]), .CO(n18294), .S(
        n18205) );
  INVXL U28364 ( .A(n18355), .Y(n18299) );
  AOI21XL U28365 ( .A0(n18301), .A1(n18300), .B0(n18299), .Y(n18308) );
  INVX1 U28366 ( .A(n23743), .Y(n18361) );
  CMPR32X1 U28367 ( .A(n18303), .B(n18302), .C(U2_A_i_d[11]), .CO(n18304), .S(
        n18256) );
  NOR2X1 U28368 ( .A(n18305), .B(n18304), .Y(n18356) );
  INVXL U28369 ( .A(n18356), .Y(n18306) );
  NAND2XL U28370 ( .A(n18305), .B(n18304), .Y(n18354) );
  NAND2XL U28371 ( .A(n18306), .B(n18354), .Y(n18307) );
  CMPR22X1 U28372 ( .A(U1_pipe14[13]), .B(n28880), .CO(n18314), .S(n18268) );
  OAI21XL U28373 ( .A0(n18322), .A1(n18321), .B0(n18320), .Y(n18431) );
  OAI21XL U28374 ( .A0(n18325), .A1(n18324), .B0(n18323), .Y(n18397) );
  CMPR22X1 U28375 ( .A(U1_pipe7[13]), .B(U1_pipe6[13]), .CO(n18327), .S(n18275) );
  OAI21XL U28376 ( .A0(n18333), .A1(n18332), .B0(n18331), .Y(n18450) );
  OAI21XL U28377 ( .A0(n18336), .A1(n18335), .B0(n18334), .Y(n18388) );
  CMPR22X1 U28378 ( .A(U1_pipe5[13]), .B(U1_pipe4[13]), .CO(n18338), .S(n18284) );
  OAI21XL U28379 ( .A0(n18344), .A1(n18343), .B0(n18342), .Y(n18469) );
  OAI21XL U28380 ( .A0(n18347), .A1(n18346), .B0(n18345), .Y(n18379) );
  CMPR22X1 U28381 ( .A(U1_pipe11[13]), .B(U1_pipe10[13]), .CO(n18349), .S(
        n18293) );
  NOR2XL U28382 ( .A(n18353), .B(n18356), .Y(n18482) );
  INVXL U28383 ( .A(n18482), .Y(n18358) );
  INVXL U28384 ( .A(n18488), .Y(n18357) );
  CMPR22X1 U28385 ( .A(U2_U0_y2[26]), .B(U2_U0_y0[26]), .CO(n23795), .S(n23743) );
  CMPR32X1 U28386 ( .A(n18361), .B(n18360), .C(U2_A_i_d[12]), .CO(n18362), .S(
        n18305) );
  INVXL U28387 ( .A(n18481), .Y(n18405) );
  CLKINVX3 U28388 ( .A(n28998), .Y(n18987) );
  OAI21XL U28389 ( .A0(n18369), .A1(n18368), .B0(n18367), .Y(n18507) );
  OAI21XL U28390 ( .A0(n18372), .A1(n18371), .B0(n18370), .Y(n18417) );
  CMPR22X1 U28391 ( .A(U1_pipe14[14]), .B(n28879), .CO(n18374), .S(n18313) );
  CMPR22X1 U28392 ( .A(U1_pipe11[14]), .B(U1_pipe10[14]), .CO(n18381), .S(
        n18348) );
  CMPR22X1 U28393 ( .A(U1_pipe5[14]), .B(U1_pipe4[14]), .CO(n18390), .S(n18337) );
  CMPR22X1 U28394 ( .A(U1_pipe7[14]), .B(U1_pipe6[14]), .CO(n18399), .S(n18326) );
  INVXL U28395 ( .A(n18486), .Y(n18411) );
  NAND2XL U28396 ( .A(n18410), .B(n18409), .Y(n18484) );
  CMPR22X1 U28397 ( .A(U1_pipe14[15]), .B(n28878), .CO(n18419), .S(n18373) );
  OAI21XL U28398 ( .A0(n18429), .A1(n18428), .B0(n18427), .Y(n18430) );
  OAI21XL U28399 ( .A0(n18435), .A1(n18434), .B0(n18433), .Y(n18436) );
  CMPR22X1 U28400 ( .A(U1_pipe7[15]), .B(U1_pipe6[15]), .CO(n18440), .S(n18398) );
  OAI21XL U28401 ( .A0(n18448), .A1(n18447), .B0(n18446), .Y(n18449) );
  OAI21XL U28402 ( .A0(n18454), .A1(n18453), .B0(n18452), .Y(n18455) );
  CMPR22X1 U28403 ( .A(U1_pipe5[15]), .B(U1_pipe4[15]), .CO(n18459), .S(n18389) );
  OAI21XL U28404 ( .A0(n18467), .A1(n18466), .B0(n18465), .Y(n18468) );
  OAI21XL U28405 ( .A0(n18473), .A1(n18472), .B0(n18471), .Y(n18474) );
  CMPR22X1 U28406 ( .A(U1_pipe11[15]), .B(U1_pipe10[15]), .CO(n18478), .S(
        n18380) );
  NAND2XL U28407 ( .A(n18482), .B(n18489), .Y(n18491) );
  NOR2XL U28408 ( .A(n18483), .B(n18491), .Y(n18494) );
  OAI21XL U28409 ( .A0(n18486), .A1(n18485), .B0(n18484), .Y(n18487) );
  AOI21XL U28410 ( .A0(n18489), .A1(n18488), .B0(n18487), .Y(n18490) );
  NAND2XL U28411 ( .A(n18545), .B(n18593), .Y(n18498) );
  XNOR2X1 U28412 ( .A(n18816), .B(n18498), .Y(n18499) );
  MXI2X1 U28413 ( .A(U2_pipe3[15]), .B(n18499), .S0(n18987), .Y(n4229) );
  OAI21XL U28414 ( .A0(n18505), .A1(n18504), .B0(n18503), .Y(n18506) );
  OAI21XL U28415 ( .A0(n18511), .A1(n18510), .B0(n18509), .Y(n18512) );
  NAND2XL U28416 ( .A(n18515), .B(n18554), .Y(n18518) );
  CMPR22X1 U28417 ( .A(U1_pipe7[16]), .B(U1_pipe6[16]), .CO(n18523), .S(n18439) );
  CMPR22X1 U28418 ( .A(U1_pipe5[16]), .B(U1_pipe4[16]), .CO(n18531), .S(n18458) );
  CMPR22X1 U28419 ( .A(U1_pipe11[16]), .B(U1_pipe10[16]), .CO(n18539), .S(
        n18477) );
  INVXL U28420 ( .A(n18593), .Y(n18544) );
  AOI21XL U28421 ( .A0(n18816), .A1(n18545), .B0(n18544), .Y(n18552) );
  INVXL U28422 ( .A(n18594), .Y(n18550) );
  NAND2XL U28423 ( .A(n18550), .B(n18592), .Y(n18551) );
  OAI21XL U28424 ( .A0(n18564), .A1(n18563), .B0(n18562), .Y(n18640) );
  CLKINVX3 U28425 ( .A(n28997), .Y(n18739) );
  OAI21XL U28426 ( .A0(n18574), .A1(n18573), .B0(n18572), .Y(n18628) );
  OAI21XL U28427 ( .A0(n18584), .A1(n18583), .B0(n18582), .Y(n18616) );
  ADDHX2 U28428 ( .A(U2_U0_y2[30]), .B(U2_U0_y0[30]), .CO(n24040), .S(n23982)
         );
  NOR2X1 U28429 ( .A(n18598), .B(n18597), .Y(n18700) );
  NAND2X1 U28430 ( .A(n18598), .B(n18597), .Y(n18703) );
  XOR2X1 U28431 ( .A(n18649), .B(n18600), .Y(n18601) );
  CMPR22X1 U28432 ( .A(U1_pipe14[18]), .B(n28875), .CO(n18608), .S(n18556) );
  CMPR22X1 U28433 ( .A(U1_pipe7[18]), .B(U1_pipe6[18]), .CO(n18620), .S(n18586) );
  CMPR22X1 U28434 ( .A(U1_pipe5[18]), .B(U1_pipe4[18]), .CO(n18632), .S(n18576) );
  CMPR22X1 U28435 ( .A(U1_pipe11[18]), .B(U1_pipe10[18]), .CO(n18644), .S(
        n18566) );
  CLKINVX2 U28436 ( .A(n24097), .Y(n18710) );
  NOR2X2 U28437 ( .A(n18653), .B(n18652), .Y(n18704) );
  NAND2XL U28438 ( .A(n18653), .B(n18652), .Y(n18702) );
  OAI21XL U28439 ( .A0(n18659), .A1(n18658), .B0(n18657), .Y(n18719) );
  OAI21XL U28440 ( .A0(n18670), .A1(n18669), .B0(n18668), .Y(n18731) );
  OAI21XL U28441 ( .A0(n18681), .A1(n18680), .B0(n18679), .Y(n18744) );
  OAI21XL U28442 ( .A0(n18692), .A1(n18691), .B0(n18690), .Y(n18756) );
  NAND2XL U28443 ( .A(n18701), .B(n18707), .Y(n18807) );
  INVXL U28444 ( .A(n18815), .Y(n18708) );
  NOR2X1 U28445 ( .A(n18713), .B(n18712), .Y(n18765) );
  XOR2X1 U28446 ( .A(n18766), .B(n18714), .Y(n18715) );
  OAI21XL U28447 ( .A0(n18722), .A1(n18721), .B0(n18720), .Y(n18776) );
  OAI21XL U28448 ( .A0(n18734), .A1(n18733), .B0(n18732), .Y(n18800) );
  OAI21XL U28449 ( .A0(n18747), .A1(n18746), .B0(n18745), .Y(n18792) );
  CLKINVX3 U28450 ( .A(n28997), .Y(n18893) );
  OAI21XL U28451 ( .A0(n18759), .A1(n18758), .B0(n18757), .Y(n18784) );
  CLKINVX2 U28452 ( .A(n24206), .Y(n18817) );
  NAND2XL U28453 ( .A(n18770), .B(n18769), .Y(n18809) );
  XNOR2X1 U28454 ( .A(n18772), .B(n18771), .Y(n18773) );
  MXI2X1 U28455 ( .A(U2_pipe3[20]), .B(n18773), .S0(n18987), .Y(n4239) );
  CMPR22X1 U28456 ( .A(U1_pipe14[21]), .B(n28872), .CO(n18778), .S(n18724) );
  CMPR22X1 U28457 ( .A(U1_pipe7[21]), .B(U1_pipe6[21]), .CO(n18786), .S(n18761) );
  CMPR22X1 U28458 ( .A(U1_pipe5[21]), .B(U1_pipe4[21]), .CO(n18794), .S(n18749) );
  CMPR22X1 U28459 ( .A(U1_pipe11[21]), .B(U1_pipe10[21]), .CO(n18802), .S(
        n18736) );
  NAND2X1 U28460 ( .A(n18806), .B(n18812), .Y(n18814) );
  INVXL U28461 ( .A(n18808), .Y(n18811) );
  INVXL U28462 ( .A(n18809), .Y(n18810) );
  AOI21XL U28463 ( .A0(n18816), .A1(n18856), .B0(n18859), .Y(n18822) );
  CMPR22X1 U28464 ( .A(U2_U0_y2[34]), .B(U2_U0_y0[34]), .CO(n24248), .S(n24207) );
  INVX1 U28465 ( .A(n24248), .Y(n18863) );
  NAND2XL U28466 ( .A(n18820), .B(n18819), .Y(n18857) );
  OAI21XL U28467 ( .A0(n18826), .A1(n18825), .B0(n18824), .Y(n18872) );
  OAI21XL U28468 ( .A0(n18834), .A1(n18833), .B0(n18832), .Y(n18880) );
  OAI21XL U28469 ( .A0(n18842), .A1(n18841), .B0(n18840), .Y(n18888) );
  OAI21XL U28470 ( .A0(n18850), .A1(n18849), .B0(n18848), .Y(n18897) );
  INVXL U28471 ( .A(n18857), .Y(n18858) );
  OAI21X1 U28472 ( .A0(n18862), .A1(n18861), .B0(n18860), .Y(n18905) );
  INVXL U28473 ( .A(n24290), .Y(n18907) );
  CMPR22X1 U28474 ( .A(U1_pipe14[23]), .B(n28953), .CO(n18874), .S(n18828) );
  CMPR22X1 U28475 ( .A(U1_pipe11[23]), .B(U1_pipe10[23]), .CO(n18882), .S(
        n18836) );
  CMPR22X1 U28476 ( .A(U1_pipe5[23]), .B(U1_pipe4[23]), .CO(n18890), .S(n18844) );
  CMPR22X1 U28477 ( .A(U1_pipe7[23]), .B(U1_pipe6[23]), .CO(n18899), .S(n18852) );
  OAI21XL U28478 ( .A0(n18913), .A1(n18912), .B0(n18911), .Y(n18949) );
  OAI21XL U28479 ( .A0(n18921), .A1(n18920), .B0(n18919), .Y(n18957) );
  OAI21XL U28480 ( .A0(n18929), .A1(n18928), .B0(n18927), .Y(n18965) );
  OAI21XL U28481 ( .A0(n18937), .A1(n18936), .B0(n18935), .Y(n18973) );
  CMPR22X1 U28482 ( .A(U2_U0_y2[37]), .B(U2_U0_y0[37]), .CO(n24372), .S(n24332) );
  CMPR32X1 U28483 ( .A(n18944), .B(n18943), .C(U2_A_i_d[23]), .CO(n18979), .S(
        n18909) );
  CMPR22X1 U28484 ( .A(U1_pipe14[25]), .B(n28951), .CO(n18951), .S(n18915) );
  CMPR22X1 U28485 ( .A(U1_pipe11[25]), .B(U1_pipe10[25]), .CO(n18959), .S(
        n18923) );
  CMPR22X1 U28486 ( .A(U1_pipe5[25]), .B(U1_pipe4[25]), .CO(n18967), .S(n18931) );
  CMPR22X1 U28487 ( .A(U1_pipe7[25]), .B(U1_pipe6[25]), .CO(n18975), .S(n18939) );
  CMPR22X1 U28488 ( .A(U2_U0_y2[38]), .B(U2_U0_y0[38]), .CO(n18981), .S(n24373) );
  XOR3X2 U28489 ( .A(n5784), .B(n18982), .C(U2_A_i_d[25]), .Y(n24375) );
  CMPR32X1 U28490 ( .A(n18984), .B(n18983), .C(U2_A_i_d[24]), .CO(n18985), .S(
        n18980) );
  CMPR22X1 U28491 ( .A(U1_pipe14[26]), .B(n29006), .CO(n18992), .S(n18950) );
  OAI21XL U28492 ( .A0(n18990), .A1(n18989), .B0(n18988), .Y(n18991) );
  CMPR32X1 U28493 ( .A(n18993), .B(n18992), .C(n18991), .S(n18994) );
  CMPR22X1 U28494 ( .A(U1_pipe7[26]), .B(U1_pipe6[26]), .CO(n18999), .S(n18974) );
  OAI21XL U28495 ( .A0(n18997), .A1(n18996), .B0(n18995), .Y(n18998) );
  CMPR32X1 U28496 ( .A(n19000), .B(n18999), .C(n18998), .S(n19001) );
  CMPR22X1 U28497 ( .A(U1_pipe5[26]), .B(U1_pipe4[26]), .CO(n19006), .S(n18966) );
  OAI21XL U28498 ( .A0(n19004), .A1(n19003), .B0(n19002), .Y(n19005) );
  CMPR32X1 U28499 ( .A(n19007), .B(n19006), .C(n19005), .S(n19008) );
  CMPR22X1 U28500 ( .A(U1_pipe11[26]), .B(U1_pipe10[26]), .CO(n19013), .S(
        n18958) );
  OAI21XL U28501 ( .A0(n19011), .A1(n19010), .B0(n19009), .Y(n19012) );
  CMPR32X1 U28502 ( .A(n19014), .B(n19013), .C(n19012), .S(n19015) );
  NOR2XL U28503 ( .A(U2_U0_y0[2]), .B(U2_U0_y1[2]), .Y(n19016) );
  NOR2XL U28504 ( .A(U2_U0_y0[3]), .B(U2_U0_y1[3]), .Y(n19022) );
  NOR2XL U28505 ( .A(n19016), .B(n19022), .Y(n19025) );
  NOR2XL U28506 ( .A(U2_U0_y0[1]), .B(U2_U0_y1[1]), .Y(n19019) );
  NAND2XL U28507 ( .A(U2_U0_y0[0]), .B(U2_U0_y1[0]), .Y(n19018) );
  NAND2XL U28508 ( .A(U2_U0_y0[1]), .B(U2_U0_y1[1]), .Y(n19017) );
  OAI21XL U28509 ( .A0(n19019), .A1(n19018), .B0(n19017), .Y(n19024) );
  NAND2XL U28510 ( .A(U2_U0_y0[2]), .B(U2_U0_y1[2]), .Y(n19021) );
  NAND2XL U28511 ( .A(U2_U0_y0[3]), .B(U2_U0_y1[3]), .Y(n19020) );
  OAI21XL U28512 ( .A0(n19022), .A1(n19021), .B0(n19020), .Y(n19023) );
  AOI21XL U28513 ( .A0(n19025), .A1(n19024), .B0(n19023), .Y(n19040) );
  NOR2XL U28514 ( .A(U2_U0_y0[4]), .B(U2_U0_y1[4]), .Y(n19026) );
  NOR2XL U28515 ( .A(U2_U0_y0[5]), .B(U2_U0_y1[5]), .Y(n19031) );
  NOR2XL U28516 ( .A(n19026), .B(n19031), .Y(n19028) );
  NOR2XL U28517 ( .A(U2_U0_y0[6]), .B(U2_U0_y1[6]), .Y(n19027) );
  NAND2XL U28518 ( .A(n19028), .B(n19037), .Y(n19039) );
  NAND2XL U28519 ( .A(U2_U0_y0[4]), .B(U2_U0_y1[4]), .Y(n19030) );
  NAND2XL U28520 ( .A(U2_U0_y0[5]), .B(U2_U0_y1[5]), .Y(n19029) );
  OAI21XL U28521 ( .A0(n19031), .A1(n19030), .B0(n19029), .Y(n19036) );
  NAND2XL U28522 ( .A(U2_U0_y0[6]), .B(U2_U0_y1[6]), .Y(n19033) );
  NAND2XL U28523 ( .A(U2_U0_y0[7]), .B(U2_U0_y1[7]), .Y(n19032) );
  OAI21XL U28524 ( .A0(n19034), .A1(n19033), .B0(n19032), .Y(n19035) );
  OAI21XL U28525 ( .A0(n19040), .A1(n19039), .B0(n19038), .Y(n19064) );
  OR2X2 U28526 ( .A(n19057), .B(n19044), .Y(n19060) );
  NAND2XL U28527 ( .A(U2_U0_y0[8]), .B(U2_U0_y1[8]), .Y(n19047) );
  NAND2XL U28528 ( .A(U2_U0_y0[9]), .B(U2_U0_y1[9]), .Y(n19046) );
  OAI21XL U28529 ( .A0(n19048), .A1(n19047), .B0(n19046), .Y(n19053) );
  NAND2XL U28530 ( .A(U2_U0_y0[10]), .B(U2_U0_y1[10]), .Y(n19050) );
  NAND2XL U28531 ( .A(U2_U0_y0[11]), .B(U2_U0_y1[11]), .Y(n19049) );
  OAI21XL U28532 ( .A0(n19051), .A1(n19050), .B0(n19049), .Y(n19052) );
  NAND2XL U28533 ( .A(U2_U0_y0[12]), .B(U2_U0_y1[12]), .Y(n19056) );
  OAI21XL U28534 ( .A0(n19057), .A1(n19056), .B0(n19055), .Y(n19058) );
  OAI21XL U28535 ( .A0(n19061), .A1(n19060), .B0(n19059), .Y(n19062) );
  CLKINVX3 U28536 ( .A(n28998), .Y(n21023) );
  INVXL U28537 ( .A(n19069), .Y(n19070) );
  OAI21XL U28538 ( .A0(n19100), .A1(n19074), .B0(n19073), .Y(n19079) );
  INVXL U28539 ( .A(n19075), .Y(n19077) );
  INVXL U28540 ( .A(n19390), .Y(n19078) );
  INVXL U28541 ( .A(n19081), .Y(n19084) );
  INVXL U28542 ( .A(n19082), .Y(n19083) );
  OAI21XL U28543 ( .A0(n19100), .A1(n19084), .B0(n19083), .Y(n19089) );
  INVXL U28544 ( .A(n19085), .Y(n19087) );
  NAND2XL U28545 ( .A(n19087), .B(n19086), .Y(n19395) );
  INVXL U28546 ( .A(n19395), .Y(n19088) );
  XNOR2X1 U28547 ( .A(n19089), .B(n19088), .Y(n19090) );
  MXI2X1 U28548 ( .A(U1_pipe2[23]), .B(n19090), .S0(n5812), .Y(n5035) );
  OAI21XL U28549 ( .A0(n19100), .A1(n19092), .B0(n19091), .Y(n19096) );
  NAND2XL U28550 ( .A(n19098), .B(n19398), .Y(n19403) );
  INVXL U28551 ( .A(n19403), .Y(n19099) );
  AOI21XL U28552 ( .A0(n19114), .A1(n19107), .B0(n19106), .Y(n19110) );
  INVXL U28553 ( .A(n19419), .Y(n19113) );
  INVXL U28554 ( .A(n19116), .Y(n19125) );
  AOI21XL U28555 ( .A0(n19125), .A1(n9689), .B0(n19117), .Y(n19121) );
  INVXL U28556 ( .A(n19127), .Y(n19130) );
  INVXL U28557 ( .A(n19128), .Y(n19129) );
  OAI21XL U28558 ( .A0(n19140), .A1(n19132), .B0(n19131), .Y(n19136) );
  AOI21XL U28559 ( .A0(n19150), .A1(n19143), .B0(n19142), .Y(n19146) );
  NAND2XL U28560 ( .A(n7024), .B(n19144), .Y(n19445) );
  NAND2XL U28561 ( .A(n19444), .B(n19148), .Y(n19448) );
  OAI21XL U28562 ( .A0(n19184), .A1(n19167), .B0(n19166), .Y(n19180) );
  INVXL U28563 ( .A(n19168), .Y(n19171) );
  INVXL U28564 ( .A(n19169), .Y(n19170) );
  INVXL U28565 ( .A(n19172), .Y(n19174) );
  NAND2XL U28566 ( .A(n19174), .B(n19173), .Y(n19465) );
  AOI21XL U28567 ( .A0(n19205), .A1(n19188), .B0(n19187), .Y(n19191) );
  INVXL U28568 ( .A(n19197), .Y(n19199) );
  OAI21XL U28569 ( .A0(n19219), .A1(n19209), .B0(n19208), .Y(n19214) );
  INVXL U28570 ( .A(n19210), .Y(n19212) );
  XOR2XL U28571 ( .A(n19225), .B(n19224), .Y(n19226) );
  XOR2XL U28572 ( .A(n19229), .B(n19228), .Y(n19230) );
  XNOR2XL U28573 ( .A(n19231), .B(U1_A_r_d0[0]), .Y(n19504) );
  MXI2X1 U28574 ( .A(U1_pipe3[27]), .B(n19232), .S0(n19215), .Y(n5067) );
  OR2X2 U28575 ( .A(n20029), .B(n19233), .Y(n19566) );
  MXI2X1 U28576 ( .A(U1_pipe3[24]), .B(n19238), .S0(n19215), .Y(n5064) );
  INVXL U28577 ( .A(n19239), .Y(n19242) );
  NAND2XL U28578 ( .A(n20041), .B(n19243), .Y(n19561) );
  XNOR2X1 U28579 ( .A(n19246), .B(n19245), .Y(n19247) );
  MXI2X1 U28580 ( .A(U1_pipe3[23]), .B(n19247), .S0(n19215), .Y(n5063) );
  NAND2XL U28581 ( .A(n20048), .B(n19248), .Y(n19558) );
  MXI2X1 U28582 ( .A(U1_pipe3[22]), .B(n19250), .S0(n19215), .Y(n5062) );
  NAND2XL U28583 ( .A(n7790), .B(n19252), .Y(n19253) );
  XOR2X1 U28584 ( .A(n19254), .B(n19253), .Y(n19255) );
  MXI2X1 U28585 ( .A(U1_pipe3[21]), .B(n19255), .S0(n19215), .Y(n5061) );
  NAND2XL U28586 ( .A(n19259), .B(n20015), .Y(n19554) );
  AOI21XL U28587 ( .A0(n19274), .A1(n19268), .B0(n8003), .Y(n19270) );
  INVXL U28588 ( .A(n19610), .Y(n19538) );
  INVXL U28589 ( .A(n19277), .Y(n19278) );
  OAI21XL U28590 ( .A0(n19289), .A1(n19280), .B0(n19286), .Y(n19284) );
  NAND2XL U28591 ( .A(n20007), .B(n19282), .Y(n19545) );
  NAND2XL U28592 ( .A(n19287), .B(n19286), .Y(n19288) );
  AOI21XL U28593 ( .A0(n19299), .A1(n14824), .B0(n19291), .Y(n19295) );
  NAND2XL U28594 ( .A(n19984), .B(n19311), .Y(n19531) );
  NAND2XL U28595 ( .A(n19310), .B(n19531), .Y(n19647) );
  OAI21XL U28596 ( .A0(n19332), .A1(n19316), .B0(n19315), .Y(n19328) );
  INVXL U28597 ( .A(n19317), .Y(n19320) );
  INVXL U28598 ( .A(n19527), .Y(n19322) );
  NAND2XL U28599 ( .A(n19979), .B(n19321), .Y(n19526) );
  NOR2XL U28600 ( .A(n19978), .B(n19326), .Y(n19524) );
  NAND2XL U28601 ( .A(n19978), .B(n19326), .Y(n19652) );
  NOR2XL U28602 ( .A(n19330), .B(n19976), .Y(n19651) );
  INVXL U28603 ( .A(n19651), .Y(n19525) );
  NAND2XL U28604 ( .A(n19330), .B(n19976), .Y(n19650) );
  NAND2XL U28605 ( .A(n19525), .B(n19650), .Y(n19661) );
  AOI21XL U28606 ( .A0(n19353), .A1(n19336), .B0(n19335), .Y(n19340) );
  OAI21XL U28607 ( .A0(n19366), .A1(n19357), .B0(n19356), .Y(n19361) );
  NOR2XL U28608 ( .A(n19358), .B(n19962), .Y(n19515) );
  INVXL U28609 ( .A(n19515), .Y(n19359) );
  NAND2XL U28610 ( .A(n19358), .B(n19962), .Y(n19514) );
  NOR2XL U28611 ( .A(n19363), .B(n19960), .Y(n19686) );
  NAND2XL U28612 ( .A(n19363), .B(n19960), .Y(n19685) );
  NOR2XL U28613 ( .A(n19369), .B(n19956), .Y(n19368) );
  INVXL U28614 ( .A(n19368), .Y(n19511) );
  NAND2XL U28615 ( .A(n19369), .B(n19956), .Y(n19508) );
  XOR2XL U28616 ( .A(n19371), .B(n19370), .Y(n19372) );
  NOR2XL U28617 ( .A(n19373), .B(n19954), .Y(n19694) );
  INVXL U28618 ( .A(n19694), .Y(n19506) );
  NAND2XL U28619 ( .A(n19373), .B(n19954), .Y(n19693) );
  XOR2XL U28620 ( .A(n19375), .B(n19374), .Y(n19376) );
  XNOR2XL U28621 ( .A(n19377), .B(n19507), .Y(n19701) );
  OAI21XL U28622 ( .A0(n19404), .A1(n19394), .B0(n19393), .Y(n19396) );
  OAI21XL U28623 ( .A0(n19404), .A1(n19399), .B0(n19398), .Y(n19401) );
  INVXL U28624 ( .A(n19410), .Y(n19413) );
  INVXL U28625 ( .A(n19411), .Y(n19412) );
  OAI21X1 U28626 ( .A0(n19420), .A1(n19415), .B0(n19414), .Y(n19417) );
  OAI21XL U28627 ( .A0(n19424), .A1(n19423), .B0(n19422), .Y(n19426) );
  XNOR2XL U28628 ( .A(n19426), .B(n19425), .Y(n19427) );
  INVXL U28629 ( .A(n19431), .Y(n19434) );
  INVXL U28630 ( .A(n19432), .Y(n19433) );
  OAI21XL U28631 ( .A0(n19441), .A1(n19436), .B0(n19435), .Y(n19438) );
  XNOR2XL U28632 ( .A(n19438), .B(n19437), .Y(n19439) );
  AOI21XL U28633 ( .A0(n19458), .A1(n13680), .B0(n19453), .Y(n19455) );
  OAI21XL U28634 ( .A0(n19472), .A1(n19461), .B0(n19460), .Y(n19469) );
  INVXL U28635 ( .A(n19462), .Y(n19463) );
  INVXL U28636 ( .A(n19474), .Y(n19487) );
  AOI21XL U28637 ( .A0(n19487), .A1(n19476), .B0(n19475), .Y(n19478) );
  OAI21XL U28638 ( .A0(n19496), .A1(n19491), .B0(n19490), .Y(n19493) );
  XOR2XL U28639 ( .A(n19499), .B(n19498), .Y(n19500) );
  XNOR2XL U28640 ( .A(n19502), .B(n19501), .Y(n19503) );
  NOR2XL U28641 ( .A(n19673), .B(n19671), .Y(n19666) );
  NAND2XL U28642 ( .A(n19666), .B(n19505), .Y(n19523) );
  NAND2XL U28643 ( .A(n19511), .B(n19506), .Y(n19513) );
  INVXL U28644 ( .A(n19693), .Y(n19510) );
  INVXL U28645 ( .A(n19508), .Y(n19509) );
  AOI21XL U28646 ( .A0(n19511), .A1(n19510), .B0(n19509), .Y(n19512) );
  OAI21XL U28647 ( .A0(n19513), .A1(n19698), .B0(n19512), .Y(n19684) );
  NOR2XL U28648 ( .A(n19515), .B(n19686), .Y(n19517) );
  OAI21XL U28649 ( .A0(n19515), .A1(n19685), .B0(n19514), .Y(n19516) );
  NAND2XL U28650 ( .A(n19518), .B(n19965), .Y(n19679) );
  NAND2XL U28651 ( .A(n19519), .B(n19967), .Y(n19674) );
  OAI21XL U28652 ( .A0(n19673), .A1(n19679), .B0(n19674), .Y(n19665) );
  NAND2XL U28653 ( .A(n19520), .B(n19969), .Y(n19667) );
  INVXL U28654 ( .A(n19667), .Y(n19521) );
  AOI21XL U28655 ( .A0(n19665), .A1(n19505), .B0(n19521), .Y(n19522) );
  NOR2XL U28656 ( .A(n19527), .B(n19524), .Y(n19530) );
  NAND2XL U28657 ( .A(n19530), .B(n19525), .Y(n19641) );
  NAND2X1 U28658 ( .A(n5788), .B(n19310), .Y(n19535) );
  NOR2X1 U28659 ( .A(n19641), .B(n19535), .Y(n19537) );
  INVXL U28660 ( .A(n19650), .Y(n19529) );
  OAI21XL U28661 ( .A0(n19527), .A1(n19652), .B0(n19526), .Y(n19528) );
  AOI21XL U28662 ( .A0(n19530), .A1(n19529), .B0(n19528), .Y(n19640) );
  NAND2XL U28663 ( .A(n19986), .B(n19532), .Y(n19643) );
  INVXL U28664 ( .A(n19643), .Y(n19533) );
  OAI21X1 U28665 ( .A0(n19640), .A1(n19535), .B0(n19534), .Y(n19536) );
  NOR2XL U28666 ( .A(n20003), .B(n19542), .Y(n19539) );
  NAND2XL U28667 ( .A(n20001), .B(n19541), .Y(n19635) );
  INVXL U28668 ( .A(n19635), .Y(n19629) );
  NAND2XL U28669 ( .A(n20003), .B(n19542), .Y(n19630) );
  INVXL U28670 ( .A(n19630), .Y(n19543) );
  NAND2XL U28671 ( .A(n20005), .B(n19544), .Y(n19624) );
  INVXL U28672 ( .A(n19624), .Y(n19547) );
  INVXL U28673 ( .A(n19545), .Y(n19546) );
  INVXL U28674 ( .A(n19550), .Y(n19551) );
  INVXL U28675 ( .A(n19554), .Y(n19555) );
  NOR2XL U28676 ( .A(n19557), .B(n20051), .Y(n19584) );
  INVXL U28677 ( .A(n19584), .Y(n19589) );
  INVXL U28678 ( .A(n19558), .Y(n19559) );
  MXI2X1 U28679 ( .A(U1_pipe1[27]), .B(n19570), .S0(n19405), .Y(n5011) );
  INVXL U28680 ( .A(n19571), .Y(n19573) );
  MXI2X1 U28681 ( .A(U1_pipe1[25]), .B(n19576), .S0(n19405), .Y(n5009) );
  MXI2X1 U28682 ( .A(U1_pipe1[24]), .B(n19577), .S0(n19405), .Y(n5008) );
  OAI21XL U28683 ( .A0(n19591), .A1(n19580), .B0(n19579), .Y(n19582) );
  XNOR2X1 U28684 ( .A(n19582), .B(n19581), .Y(n19583) );
  MXI2X1 U28685 ( .A(U1_pipe1[23]), .B(n19583), .S0(n25330), .Y(n5154) );
  OAI21XL U28686 ( .A0(n19591), .A1(n19584), .B0(n19588), .Y(n19586) );
  XNOR2X1 U28687 ( .A(n19586), .B(n19585), .Y(n19587) );
  MXI2X1 U28688 ( .A(U1_pipe1[22]), .B(n19587), .S0(n25330), .Y(n5153) );
  NAND2XL U28689 ( .A(n19589), .B(n19588), .Y(n19590) );
  MXI2X1 U28690 ( .A(U1_pipe1[21]), .B(n19592), .S0(n25330), .Y(n5152) );
  CLKINVX3 U28691 ( .A(n19593), .Y(n19637) );
  INVXL U28692 ( .A(n19596), .Y(n19599) );
  XNOR2X1 U28693 ( .A(n19602), .B(n19601), .Y(n19603) );
  MXI2X1 U28694 ( .A(U1_pipe1[20]), .B(n19603), .S0(n25330), .Y(n5151) );
  NAND2XL U28695 ( .A(n19605), .B(n19604), .Y(n19606) );
  XOR2X1 U28696 ( .A(n19607), .B(n19606), .Y(n19608) );
  OAI21XL U28697 ( .A0(n6232), .A1(n19610), .B0(n19609), .Y(n19612) );
  XNOR2X1 U28698 ( .A(n19612), .B(n19611), .Y(n19613) );
  MXI2X1 U28699 ( .A(U1_pipe1[18]), .B(n19613), .S0(n19405), .Y(n5149) );
  INVXL U28700 ( .A(n19616), .Y(n19619) );
  INVXL U28701 ( .A(n19617), .Y(n19618) );
  OAI21XL U28702 ( .A0(n19627), .A1(n19620), .B0(n19624), .Y(n19622) );
  XNOR2XL U28703 ( .A(n19622), .B(n19621), .Y(n19623) );
  MXI2X1 U28704 ( .A(U1_pipe1[16]), .B(n19623), .S0(n20025), .Y(n5147) );
  NAND2XL U28705 ( .A(n19625), .B(n19624), .Y(n19626) );
  XOR2X1 U28706 ( .A(n19627), .B(n19626), .Y(n19628) );
  NAND2XL U28707 ( .A(n19631), .B(n19630), .Y(n19632) );
  NAND2XL U28708 ( .A(n19540), .B(n19635), .Y(n19636) );
  XNOR2X1 U28709 ( .A(n19637), .B(n19636), .Y(n19638) );
  OAI21XL U28710 ( .A0(n19662), .A1(n19651), .B0(n19650), .Y(n19659) );
  AOI21XL U28711 ( .A0(n19682), .A1(n19666), .B0(n19665), .Y(n19669) );
  INVXL U28712 ( .A(n19673), .Y(n19675) );
  INVXL U28713 ( .A(n19684), .Y(n19691) );
  OAI21XL U28714 ( .A0(n19691), .A1(n19686), .B0(n19685), .Y(n19688) );
  OAI21XL U28715 ( .A0(n19698), .A1(n19694), .B0(n19693), .Y(n19696) );
  XOR2XL U28716 ( .A(n19699), .B(n19698), .Y(n19700) );
  NAND2XL U28717 ( .A(U1_pipe1[0]), .B(U1_pipe0[0]), .Y(n19703) );
  OAI21XL U28718 ( .A0(n19704), .A1(n19703), .B0(n19702), .Y(n20527) );
  NOR2XL U28719 ( .A(n19724), .B(U1_A_r_d0[6]), .Y(n19726) );
  NOR2XL U28720 ( .A(n19723), .B(U1_A_r_d0[5]), .Y(n19913) );
  NOR2XL U28721 ( .A(n19726), .B(n19913), .Y(n19908) );
  OR2X2 U28722 ( .A(n19727), .B(U1_A_r_d0[7]), .Y(n19729) );
  NAND2XL U28723 ( .A(n19908), .B(n19729), .Y(n19731) );
  NOR2XL U28724 ( .A(n19718), .B(U1_A_r_d0[4]), .Y(n19720) );
  NOR2XL U28725 ( .A(n19720), .B(n19929), .Y(n19722) );
  AOI21XL U28726 ( .A0(n19713), .A1(n19710), .B0(n19712), .Y(n19943) );
  OAI21XL U28727 ( .A0(n19943), .A1(n19716), .B0(n19715), .Y(n19927) );
  NAND2XL U28728 ( .A(n19718), .B(U1_A_r_d0[4]), .Y(n19719) );
  OAI21XL U28729 ( .A0(n19720), .A1(n19928), .B0(n19719), .Y(n19721) );
  AOI21XL U28730 ( .A0(n19722), .A1(n19927), .B0(n19721), .Y(n19906) );
  NAND2XL U28731 ( .A(n19723), .B(U1_A_r_d0[5]), .Y(n19914) );
  NAND2XL U28732 ( .A(n19724), .B(U1_A_r_d0[6]), .Y(n19725) );
  OAI21XL U28733 ( .A0(n19726), .A1(n19914), .B0(n19725), .Y(n19907) );
  AOI21XL U28734 ( .A0(n19907), .A1(n19729), .B0(n19728), .Y(n19730) );
  OAI21XL U28735 ( .A0(n19731), .A1(n19906), .B0(n19730), .Y(n19872) );
  NOR2XL U28736 ( .A(n8657), .B(U1_A_r_d0[9]), .Y(n19888) );
  NOR2XL U28737 ( .A(n19740), .B(n19888), .Y(n19743) );
  NOR2XL U28738 ( .A(n19737), .B(U1_A_r_d0[8]), .Y(n19887) );
  INVXL U28739 ( .A(n19887), .Y(n19733) );
  NAND2XL U28740 ( .A(n19743), .B(n19733), .Y(n19874) );
  OR2X2 U28741 ( .A(n19744), .B(U1_A_r_d0[11]), .Y(n19876) );
  NAND2XL U28742 ( .A(n19735), .B(n19876), .Y(n19748) );
  NOR2XL U28743 ( .A(n19874), .B(n19748), .Y(n19750) );
  INVXL U28744 ( .A(n19886), .Y(n19742) );
  NAND2XL U28745 ( .A(n8657), .B(U1_A_r_d0[9]), .Y(n19889) );
  NAND2XL U28746 ( .A(n19738), .B(U1_A_r_d0[10]), .Y(n19739) );
  OAI21XL U28747 ( .A0(n19740), .A1(n19889), .B0(n19739), .Y(n19741) );
  AOI21XL U28748 ( .A0(n19735), .A1(n19875), .B0(n19746), .Y(n19747) );
  NOR2XL U28749 ( .A(n19761), .B(U1_A_r_d0[16]), .Y(n19752) );
  NOR2XL U28750 ( .A(n19760), .B(U1_A_r_d0[15]), .Y(n19852) );
  INVXL U28751 ( .A(n19852), .Y(n19753) );
  OR2X2 U28752 ( .A(n19757), .B(U1_A_r_d0[13]), .Y(n19863) );
  NAND2XL U28753 ( .A(n19755), .B(n19863), .Y(n19847) );
  OR2X2 U28754 ( .A(n19767), .B(U1_A_r_d0[19]), .Y(n19827) );
  OR2X2 U28755 ( .A(n19765), .B(U1_A_r_d0[17]), .Y(n19837) );
  NAND2X1 U28756 ( .A(n19766), .B(n19837), .Y(n19825) );
  AND2X2 U28757 ( .A(n19757), .B(U1_A_r_d0[13]), .Y(n19862) );
  NAND2XL U28758 ( .A(n19760), .B(U1_A_r_d0[15]), .Y(n19851) );
  AND2X2 U28759 ( .A(n19765), .B(U1_A_r_d0[17]), .Y(n19836) );
  AND2X2 U28760 ( .A(n19767), .B(U1_A_r_d0[19]), .Y(n19826) );
  NOR2XL U28761 ( .A(n19776), .B(U1_A_r_d0[21]), .Y(n19812) );
  NOR2XL U28762 ( .A(n19782), .B(U1_A_r_d0[24]), .Y(n19784) );
  NAND2XL U28763 ( .A(n19776), .B(U1_A_r_d0[21]), .Y(n19811) );
  NAND2XL U28764 ( .A(n19777), .B(U1_A_r_d0[22]), .Y(n19778) );
  NAND2XL U28765 ( .A(n19782), .B(U1_A_r_d0[24]), .Y(n19783) );
  NOR2XL U28766 ( .A(n19786), .B(U1_A_r_d0[25]), .Y(n19788) );
  NAND2XL U28767 ( .A(n19786), .B(U1_A_r_d0[25]), .Y(n19787) );
  MXI2X1 U28768 ( .A(U1_pipe12[27]), .B(n19789), .S0(n25330), .Y(n4722) );
  INVXL U28769 ( .A(n20189), .Y(n19792) );
  XOR2X1 U28770 ( .A(n19793), .B(n19792), .Y(n19794) );
  OAI21XL U28771 ( .A0(n19820), .A1(n19796), .B0(n19795), .Y(n19800) );
  NAND2XL U28772 ( .A(n19797), .B(n19798), .Y(n20192) );
  INVXL U28773 ( .A(n20192), .Y(n19799) );
  INVXL U28774 ( .A(n19803), .Y(n19804) );
  INVXL U28775 ( .A(n19805), .Y(n19807) );
  XNOR2X1 U28776 ( .A(n19809), .B(n19808), .Y(n19810) );
  OAI21XL U28777 ( .A0(n19820), .A1(n19812), .B0(n19811), .Y(n19816) );
  XNOR2X1 U28778 ( .A(n19816), .B(n19815), .Y(n19817) );
  XOR2X1 U28779 ( .A(n19831), .B(n19830), .Y(n19832) );
  NAND2XL U28780 ( .A(n19833), .B(n20215), .Y(n20220) );
  INVXL U28781 ( .A(n19835), .Y(n19845) );
  AOI21XL U28782 ( .A0(n19845), .A1(n19837), .B0(n19836), .Y(n19841) );
  INVXL U28783 ( .A(n19848), .Y(n19849) );
  OAI21XL U28784 ( .A0(n19860), .A1(n19852), .B0(n19851), .Y(n19856) );
  AOI21XL U28785 ( .A0(n19870), .A1(n19863), .B0(n19862), .Y(n19866) );
  OAI21XL U28786 ( .A0(n19904), .A1(n19874), .B0(n19873), .Y(n19884) );
  AOI21XL U28787 ( .A0(n19884), .A1(n19876), .B0(n19875), .Y(n19880) );
  OAI21XL U28788 ( .A0(n19904), .A1(n19887), .B0(n19886), .Y(n19900) );
  AOI21XL U28789 ( .A0(n19925), .A1(n19908), .B0(n19907), .Y(n19911) );
  OAI21XL U28790 ( .A0(n19938), .A1(n19929), .B0(n19928), .Y(n19934) );
  XOR2XL U28791 ( .A(n19944), .B(n19943), .Y(n19945) );
  XOR2XL U28792 ( .A(n19948), .B(n19947), .Y(n19949) );
  XNOR2XL U28793 ( .A(n16780), .B(U1_A_r_d0[0]), .Y(n20307) );
  NOR2XL U28794 ( .A(n20145), .B(n20143), .Y(n20138) );
  NAND2XL U28795 ( .A(n20138), .B(n19950), .Y(n19973) );
  NOR2XL U28796 ( .A(n5883), .B(n19962), .Y(n20159) );
  NOR2XL U28797 ( .A(n19961), .B(n19960), .Y(n20158) );
  NOR2XL U28798 ( .A(n20159), .B(n20158), .Y(n19964) );
  NOR2XL U28799 ( .A(n20180), .B(n20179), .Y(n20176) );
  AOI21XL U28800 ( .A0(n19955), .A1(n19953), .B0(n8010), .Y(n20172) );
  NOR2XL U28801 ( .A(n19957), .B(n19956), .Y(n19959) );
  NAND2XL U28802 ( .A(n19957), .B(n19956), .Y(n19958) );
  OAI21XL U28803 ( .A0(n20172), .A1(n19959), .B0(n19958), .Y(n20156) );
  NAND2XL U28804 ( .A(n19961), .B(n19960), .Y(n20157) );
  NAND2XL U28805 ( .A(n5883), .B(n19962), .Y(n20160) );
  OAI21XL U28806 ( .A0(n20159), .A1(n20157), .B0(n20160), .Y(n19963) );
  AOI21XL U28807 ( .A0(n19964), .A1(n20156), .B0(n19963), .Y(n20136) );
  NAND2XL U28808 ( .A(n19968), .B(n19967), .Y(n20146) );
  OAI21XL U28809 ( .A0(n20145), .A1(n20151), .B0(n20146), .Y(n20137) );
  AOI21XL U28810 ( .A0(n20137), .A1(n19950), .B0(n19971), .Y(n19972) );
  OAI21XL U28811 ( .A0(n19973), .A1(n20136), .B0(n19972), .Y(n20103) );
  NOR2XL U28812 ( .A(n14934), .B(n19978), .Y(n20119) );
  NOR2XL U28813 ( .A(n19977), .B(n19976), .Y(n20118) );
  INVXL U28814 ( .A(n20118), .Y(n19975) );
  NAND2XL U28815 ( .A(n19983), .B(n19975), .Y(n20105) );
  NOR2XL U28816 ( .A(n20105), .B(n19990), .Y(n19992) );
  NAND2XL U28817 ( .A(n14934), .B(n19978), .Y(n20127) );
  NAND2XL U28818 ( .A(n19980), .B(n19979), .Y(n20122) );
  OAI21XL U28819 ( .A0(n20121), .A1(n20127), .B0(n20122), .Y(n19981) );
  AOI21XL U28820 ( .A0(n19983), .A1(n19982), .B0(n19981), .Y(n20104) );
  NAND2XL U28821 ( .A(n19985), .B(n19984), .Y(n20112) );
  INVXL U28822 ( .A(n20112), .Y(n20106) );
  NAND2XL U28823 ( .A(n19987), .B(n19986), .Y(n20107) );
  INVXL U28824 ( .A(n20107), .Y(n19988) );
  OAI21XL U28825 ( .A0(n20104), .A1(n19990), .B0(n19989), .Y(n19991) );
  NOR2XL U28826 ( .A(n20006), .B(n20005), .Y(n20083) );
  NAND2XL U28827 ( .A(n6938), .B(n19995), .Y(n20079) );
  NOR2XL U28828 ( .A(n20014), .B(n20013), .Y(n19997) );
  INVXL U28829 ( .A(n19997), .Y(n20059) );
  INVXL U28830 ( .A(n20000), .Y(n20070) );
  NAND2XL U28831 ( .A(n20002), .B(n20001), .Y(n20099) );
  INVXL U28832 ( .A(n20099), .Y(n20094) );
  NAND2XL U28833 ( .A(n7434), .B(n20003), .Y(n20095) );
  NAND2XL U28834 ( .A(n20006), .B(n20005), .Y(n20089) );
  INVXL U28835 ( .A(n20089), .Y(n20009) );
  NAND2XL U28836 ( .A(n5859), .B(n20007), .Y(n20084) );
  INVXL U28837 ( .A(n20084), .Y(n20008) );
  NAND2XL U28838 ( .A(n5817), .B(n20015), .Y(n20060) );
  NAND2XL U28839 ( .A(n20016), .B(n20051), .Y(n20045) );
  NAND2XL U28840 ( .A(n5850), .B(n20048), .Y(n20017) );
  NAND2XL U28841 ( .A(n20020), .B(n20033), .Y(n20021) );
  MXI2X1 U28842 ( .A(U1_pipe13[26]), .B(n20027), .S0(n20025), .Y(n4749) );
  OAI21XL U28843 ( .A0(n20053), .A1(n20031), .B0(n20030), .Y(n20035) );
  XNOR2X1 U28844 ( .A(n20035), .B(n20034), .Y(n20036) );
  MXI2X1 U28845 ( .A(U1_pipe13[24]), .B(n20036), .S0(n20025), .Y(n4747) );
  INVXL U28846 ( .A(n20038), .Y(n20039) );
  MXI2X1 U28847 ( .A(U1_pipe13[23]), .B(n20044), .S0(n20025), .Y(n4746) );
  NAND2XL U28848 ( .A(n20048), .B(n20047), .Y(n20322) );
  XOR2X1 U28849 ( .A(n20053), .B(n20052), .Y(n20054) );
  AOI21X1 U28850 ( .A0(n20101), .A1(n20056), .B0(n20055), .Y(n20069) );
  XOR2X1 U28851 ( .A(n20063), .B(n20062), .Y(n20064) );
  MXI2X1 U28852 ( .A(U1_pipe13[20]), .B(n20064), .S0(n20025), .Y(n4743) );
  XNOR2X1 U28853 ( .A(n20067), .B(n20066), .Y(n20068) );
  AOI21XL U28854 ( .A0(n20077), .A1(n20070), .B0(n6901), .Y(n20074) );
  XOR2X1 U28855 ( .A(n20074), .B(n20073), .Y(n20075) );
  NAND2XL U28856 ( .A(n20356), .B(n20355), .Y(n20360) );
  INVXL U28857 ( .A(n20080), .Y(n20081) );
  OAI21XL U28858 ( .A0(n20092), .A1(n20083), .B0(n20089), .Y(n20087) );
  AOI21XL U28859 ( .A0(n20101), .A1(n19995), .B0(n20094), .Y(n20097) );
  NAND2XL U28860 ( .A(n6938), .B(n20095), .Y(n20096) );
  NAND2XL U28861 ( .A(n19995), .B(n20099), .Y(n20100) );
  OAI21XL U28862 ( .A0(n20134), .A1(n20105), .B0(n20104), .Y(n20115) );
  AOI21XL U28863 ( .A0(n20115), .A1(n20113), .B0(n20106), .Y(n20110) );
  NAND2XL U28864 ( .A(n20113), .B(n20112), .Y(n20114) );
  OAI21XL U28865 ( .A0(n20134), .A1(n20118), .B0(n20117), .Y(n20130) );
  INVXL U28866 ( .A(n20119), .Y(n20128) );
  INVXL U28867 ( .A(n20127), .Y(n20120) );
  NAND2XL U28868 ( .A(n20128), .B(n20127), .Y(n20129) );
  NAND2XL U28869 ( .A(n20132), .B(n20401), .Y(n20416) );
  INVXL U28870 ( .A(n20136), .Y(n20154) );
  AOI21XL U28871 ( .A0(n20154), .A1(n20138), .B0(n20137), .Y(n20141) );
  OAI21XL U28872 ( .A0(n20167), .A1(n20158), .B0(n20157), .Y(n20163) );
  INVXL U28873 ( .A(n20159), .Y(n20161) );
  NAND2XL U28874 ( .A(n20165), .B(n20441), .Y(n20449) );
  INVXL U28875 ( .A(n20169), .Y(n20171) );
  XOR2XL U28876 ( .A(n20173), .B(n20172), .Y(n20174) );
  XOR2XL U28877 ( .A(n20177), .B(n20176), .Y(n20178) );
  XNOR2XL U28878 ( .A(n20180), .B(n20179), .Y(n20458) );
  OR2XL U28879 ( .A(U1_pipe13[1]), .B(U1_pipe12[1]), .Y(n20185) );
  OR2XL U28880 ( .A(n28910), .B(U1_pipe12[0]), .Y(n20184) );
  MXI2X1 U28881 ( .A(U1_pipe8[26]), .B(n20188), .S0(n20240), .Y(n4808) );
  XNOR2X1 U28882 ( .A(n20190), .B(n20189), .Y(n20191) );
  OAI21XL U28883 ( .A0(n20206), .A1(n20196), .B0(n20195), .Y(n20198) );
  XNOR2XL U28884 ( .A(n20198), .B(n20197), .Y(n20199) );
  OAI21XL U28885 ( .A0(n20206), .A1(n20201), .B0(n20200), .Y(n20203) );
  XNOR2XL U28886 ( .A(n20203), .B(n20202), .Y(n20204) );
  INVX1 U28887 ( .A(n20208), .Y(n20251) );
  AOI21X1 U28888 ( .A0(n20251), .A1(n20210), .B0(n20209), .Y(n20225) );
  OAI21XL U28889 ( .A0(n20221), .A1(n20216), .B0(n20215), .Y(n20218) );
  XNOR2X1 U28890 ( .A(n20218), .B(n20217), .Y(n20219) );
  OAI21XL U28891 ( .A0(n20225), .A1(n20224), .B0(n20223), .Y(n20227) );
  XNOR2XL U28892 ( .A(n20227), .B(n20226), .Y(n20228) );
  INVXL U28893 ( .A(n20233), .Y(n20234) );
  AOI21XL U28894 ( .A0(n20251), .A1(n20235), .B0(n20234), .Y(n20243) );
  OAI21XL U28895 ( .A0(n20243), .A1(n20237), .B0(n20236), .Y(n20239) );
  XNOR2XL U28896 ( .A(n20239), .B(n20238), .Y(n20241) );
  OAI21XL U28897 ( .A0(n20275), .A1(n20255), .B0(n20254), .Y(n20261) );
  AOI21XL U28898 ( .A0(n20261), .A1(n12300), .B0(n20256), .Y(n20258) );
  OAI21XL U28899 ( .A0(n20275), .A1(n20264), .B0(n20263), .Y(n20272) );
  OAI21XL U28900 ( .A0(n20299), .A1(n20294), .B0(n20293), .Y(n20296) );
  XOR2XL U28901 ( .A(n20302), .B(n20301), .Y(n20303) );
  XNOR2XL U28902 ( .A(n20305), .B(n20304), .Y(n20306) );
  INVXL U28903 ( .A(n20311), .Y(n20314) );
  INVXL U28904 ( .A(n20312), .Y(n20313) );
  INVXL U28905 ( .A(n20344), .Y(n20325) );
  INVXL U28906 ( .A(n20322), .Y(n20323) );
  MXI2X1 U28907 ( .A(U1_pipe9[27]), .B(n20334), .S0(n20240), .Y(n4837) );
  MXI2X1 U28908 ( .A(U1_pipe9[24]), .B(n20340), .S0(n20240), .Y(n4834) );
  MXI2X1 U28909 ( .A(U1_pipe9[23]), .B(n20343), .S0(n20240), .Y(n4833) );
  XNOR2X1 U28910 ( .A(n20347), .B(n20346), .Y(n20348) );
  MXI2X1 U28911 ( .A(U1_pipe9[22]), .B(n20348), .S0(n20240), .Y(n4832) );
  XOR2X1 U28912 ( .A(n20350), .B(n20349), .Y(n20351) );
  XNOR2XL U28913 ( .A(n20358), .B(n20357), .Y(n20359) );
  INVXL U28914 ( .A(n20363), .Y(n20366) );
  INVXL U28915 ( .A(n20364), .Y(n20365) );
  OAI21XL U28916 ( .A0(n20375), .A1(n20367), .B0(n20372), .Y(n20370) );
  NAND2XL U28917 ( .A(n7005), .B(n20368), .Y(n20369) );
  NAND2XL U28918 ( .A(n20373), .B(n20372), .Y(n20374) );
  OAI21XL U28919 ( .A0(n20417), .A1(n20390), .B0(n20389), .Y(n20399) );
  AOI21XL U28920 ( .A0(n20399), .A1(n14874), .B0(n20391), .Y(n20395) );
  NAND2XL U28921 ( .A(n14874), .B(n20397), .Y(n20398) );
  OAI21XL U28922 ( .A0(n20417), .A1(n20402), .B0(n20401), .Y(n20414) );
  INVXL U28923 ( .A(n20403), .Y(n20412) );
  INVXL U28924 ( .A(n20411), .Y(n20404) );
  NAND2XL U28925 ( .A(n20412), .B(n20411), .Y(n20413) );
  AOI21XL U28926 ( .A0(n20437), .A1(n20421), .B0(n20420), .Y(n20424) );
  INVXL U28927 ( .A(n20428), .Y(n20430) );
  INVXL U28928 ( .A(n20440), .Y(n20450) );
  OAI21XL U28929 ( .A0(n20450), .A1(n20442), .B0(n20441), .Y(n20447) );
  INVXL U28930 ( .A(n20443), .Y(n20445) );
  XOR2XL U28931 ( .A(n20453), .B(n20452), .Y(n20454) );
  XNOR2XL U28932 ( .A(n20456), .B(n20455), .Y(n20457) );
  OAI21XL U28933 ( .A0(n24411), .A1(n20467), .B0(n20466), .Y(n20553) );
  INVXL U28934 ( .A(n25848), .Y(n20508) );
  CMPR22X1 U28935 ( .A(U2_U0_y1[14]), .B(U2_U0_y0[14]), .CO(n25847), .S(n25800) );
  OR2X2 U28936 ( .A(n20469), .B(n20468), .Y(n20506) );
  NOR2XL U28937 ( .A(n20470), .B(U2_A_r_d[1]), .Y(n20547) );
  OAI21XL U28938 ( .A0(n20476), .A1(n20475), .B0(n20474), .Y(n20595) );
  CMPR22X1 U28939 ( .A(U1_pipe2[2]), .B(n28736), .CO(n20478), .S(n19378) );
  OAI21XL U28940 ( .A0(n20482), .A1(n20522), .B0(n20524), .Y(n20487) );
  CMPR22X1 U28941 ( .A(U1_pipe1[2]), .B(U1_pipe0[2]), .CO(n20484), .S(n19705)
         );
  OAI21XL U28942 ( .A0(n20491), .A1(n20490), .B0(n20489), .Y(n20584) );
  CMPR22X1 U28943 ( .A(U1_pipe12[2]), .B(n28740), .CO(n20493), .S(n20181) );
  OAI21XL U28944 ( .A0(n20499), .A1(n20498), .B0(n20497), .Y(n20565) );
  CMPR22X1 U28945 ( .A(U1_pipe8[2]), .B(n28732), .CO(n20501), .S(n20459) );
  OAI21XL U28946 ( .A0(n20505), .A1(n20547), .B0(n20549), .Y(n20513) );
  INVXL U28947 ( .A(n25887), .Y(n20554) );
  CMPR32X1 U28948 ( .A(n20508), .B(n20507), .C(n20506), .CO(n20509), .S(n20470) );
  OAI21XL U28949 ( .A0(n20515), .A1(n20590), .B0(n20592), .Y(n20520) );
  CMPR22X1 U28950 ( .A(U1_pipe2[3]), .B(n28735), .CO(n20517), .S(n20477) );
  OAI21XL U28951 ( .A0(n20525), .A1(n20524), .B0(n20523), .Y(n20526) );
  CMPR22X1 U28952 ( .A(U1_pipe1[3]), .B(U1_pipe0[3]), .CO(n20530), .S(n20483)
         );
  OAI21XL U28953 ( .A0(n20533), .A1(n20579), .B0(n20581), .Y(n20538) );
  CMPR22X1 U28954 ( .A(U1_pipe12[3]), .B(n28739), .CO(n20535), .S(n20492) );
  OAI21XL U28955 ( .A0(n20540), .A1(n20560), .B0(n20562), .Y(n20545) );
  CMPR22X1 U28956 ( .A(U1_pipe8[3]), .B(n28731), .CO(n20542), .S(n20500) );
  NOR2XL U28957 ( .A(n20550), .B(n20547), .Y(n20552) );
  OAI21XL U28958 ( .A0(n20550), .A1(n20549), .B0(n20548), .Y(n20551) );
  AOI21XL U28959 ( .A0(n20553), .A1(n20552), .B0(n20551), .Y(n20750) );
  INVXL U28960 ( .A(n25944), .Y(n20604) );
  INVXL U28961 ( .A(n25943), .Y(n20603) );
  CMPR32X1 U28962 ( .A(n20555), .B(n20554), .C(U2_A_r_d[2]), .CO(n20556), .S(
        n20510) );
  NAND2XL U28963 ( .A(n20557), .B(n20556), .Y(n20647) );
  OAI21XL U28964 ( .A0(n20563), .A1(n20562), .B0(n20561), .Y(n20564) );
  CMPR22X1 U28965 ( .A(U1_pipe8[4]), .B(n28839), .CO(n20568), .S(n20541) );
  CMPR22X1 U28966 ( .A(U1_pipe1[4]), .B(U1_pipe0[4]), .CO(n20574), .S(n20529)
         );
  OAI21XL U28967 ( .A0(n20582), .A1(n20581), .B0(n20580), .Y(n20583) );
  CMPR22X1 U28968 ( .A(U1_pipe12[4]), .B(n28871), .CO(n20587), .S(n20534) );
  OAI21XL U28969 ( .A0(n20593), .A1(n20592), .B0(n20591), .Y(n20594) );
  CMPR22X1 U28970 ( .A(U1_pipe2[4]), .B(n28855), .CO(n20598), .S(n20516) );
  INVXL U28971 ( .A(n25986), .Y(n20651) );
  INVXL U28972 ( .A(n25985), .Y(n20650) );
  CMPR32X1 U28973 ( .A(n20604), .B(n20603), .C(U2_A_r_d[3]), .CO(n20605), .S(
        n20557) );
  INVXL U28974 ( .A(n20648), .Y(n20607) );
  NAND2XL U28975 ( .A(n20606), .B(n20605), .Y(n20646) );
  CMPR22X1 U28976 ( .A(U1_pipe2[5]), .B(n28854), .CO(n20614), .S(n20597) );
  OAI21XL U28977 ( .A0(n20622), .A1(n20621), .B0(n20620), .Y(n20716) );
  CMPR22X1 U28978 ( .A(U1_pipe1[5]), .B(U1_pipe0[5]), .CO(n20625), .S(n20573)
         );
  CMPR22X1 U28979 ( .A(U1_pipe12[5]), .B(n28870), .CO(n20632), .S(n20586) );
  CMPR22X1 U28980 ( .A(U1_pipe8[5]), .B(n28838), .CO(n20640), .S(n20567) );
  NOR2XL U28981 ( .A(n20645), .B(n20648), .Y(n20741) );
  OAI21XL U28982 ( .A0(n20648), .A1(n20647), .B0(n20646), .Y(n20746) );
  AOI21XL U28983 ( .A0(n20649), .A1(n20741), .B0(n20746), .Y(n20694) );
  INVXL U28984 ( .A(n26036), .Y(n20696) );
  INVXL U28985 ( .A(n26035), .Y(n20695) );
  CMPR32X1 U28986 ( .A(n20651), .B(n20650), .C(U2_A_r_d[4]), .CO(n20652), .S(
        n20606) );
  INVXL U28987 ( .A(n20740), .Y(n20654) );
  NAND2XL U28988 ( .A(n20653), .B(n20652), .Y(n20743) );
  OAI21XL U28989 ( .A0(n20660), .A1(n20659), .B0(n20658), .Y(n20802) );
  CMPR22X1 U28990 ( .A(U1_pipe2[6]), .B(n28734), .CO(n20663), .S(n20613) );
  OAI21XL U28991 ( .A0(n20667), .A1(n20710), .B0(n20713), .Y(n20672) );
  CMPR22X1 U28992 ( .A(U1_pipe1[6]), .B(U1_pipe0[6]), .CO(n20669), .S(n20624)
         );
  OAI21XL U28993 ( .A0(n20677), .A1(n20676), .B0(n20675), .Y(n20786) );
  CMPR22X1 U28994 ( .A(U1_pipe12[6]), .B(n28738), .CO(n20680), .S(n20631) );
  OAI21XL U28995 ( .A0(n20687), .A1(n20686), .B0(n20685), .Y(n20764) );
  CMPR22X1 U28996 ( .A(U1_pipe8[6]), .B(n28730), .CO(n20690), .S(n20639) );
  OAI21XL U28997 ( .A0(n20694), .A1(n20740), .B0(n20743), .Y(n20701) );
  INVXL U28998 ( .A(n26081), .Y(n20752) );
  INVXL U28999 ( .A(n26080), .Y(n20751) );
  CMPR32X1 U29000 ( .A(n20696), .B(n20695), .C(U2_A_r_d[5]), .CO(n20697), .S(
        n20653) );
  INVXL U29001 ( .A(n20744), .Y(n20699) );
  NAND2XL U29002 ( .A(n20698), .B(n20697), .Y(n20742) );
  OAI21XL U29003 ( .A0(n20703), .A1(n20758), .B0(n20761), .Y(n20708) );
  CMPR22X1 U29004 ( .A(U1_pipe8[7]), .B(n28837), .CO(n20705), .S(n20689) );
  OAI21XL U29005 ( .A0(n20714), .A1(n20713), .B0(n20712), .Y(n20715) );
  OAI21XL U29006 ( .A0(n20720), .A1(n20719), .B0(n20718), .Y(n21161) );
  CMPR22X1 U29007 ( .A(U1_pipe1[7]), .B(U1_pipe0[7]), .CO(n20722), .S(n20668)
         );
  OAI21XL U29008 ( .A0(n20726), .A1(n20780), .B0(n20783), .Y(n20731) );
  CMPR22X1 U29009 ( .A(U1_pipe12[7]), .B(n28869), .CO(n20728), .S(n20679) );
  OAI21XL U29010 ( .A0(n20733), .A1(n20796), .B0(n20799), .Y(n20738) );
  CMPR22X1 U29011 ( .A(U1_pipe2[7]), .B(n28853), .CO(n20735), .S(n20662) );
  NOR2XL U29012 ( .A(n20740), .B(n20744), .Y(n20747) );
  NAND2XL U29013 ( .A(n20741), .B(n20747), .Y(n20749) );
  OAI21XL U29014 ( .A0(n20744), .A1(n20743), .B0(n20742), .Y(n20745) );
  AOI21XL U29015 ( .A0(n20747), .A1(n20746), .B0(n20745), .Y(n20748) );
  OAI21XL U29016 ( .A0(n20750), .A1(n20749), .B0(n20748), .Y(n21189) );
  INVXL U29017 ( .A(n26154), .Y(n20813) );
  INVXL U29018 ( .A(n26153), .Y(n20812) );
  CMPR32X1 U29019 ( .A(n20752), .B(n20751), .C(U2_A_r_d[6]), .CO(n20753), .S(
        n20698) );
  NAND2XL U29020 ( .A(n20755), .B(n20850), .Y(n20756) );
  OAI21XL U29021 ( .A0(n20762), .A1(n20761), .B0(n20760), .Y(n20763) );
  OAI21XL U29022 ( .A0(n20768), .A1(n20767), .B0(n20766), .Y(n21258) );
  CMPR22X1 U29023 ( .A(U1_pipe8[8]), .B(n28836), .CO(n20770), .S(n20704) );
  NAND2XL U29024 ( .A(n20771), .B(n20891), .Y(n20772) );
  OAI21XL U29025 ( .A0(n20927), .A1(n20826), .B0(n20828), .Y(n20778) );
  CMPR22X1 U29026 ( .A(U1_pipe1[8]), .B(U1_pipe0[8]), .CO(n20775), .S(n20721)
         );
  OAI21XL U29027 ( .A0(n20784), .A1(n20783), .B0(n20782), .Y(n20785) );
  OAI21XL U29028 ( .A0(n20790), .A1(n20789), .B0(n20788), .Y(n21210) );
  CMPR22X1 U29029 ( .A(U1_pipe12[8]), .B(n28868), .CO(n20792), .S(n20727) );
  OAI21XL U29030 ( .A0(n20800), .A1(n20799), .B0(n20798), .Y(n20801) );
  OAI21XL U29031 ( .A0(n20806), .A1(n20805), .B0(n20804), .Y(n21230) );
  CMPR22X1 U29032 ( .A(U1_pipe2[8]), .B(n28852), .CO(n20808), .S(n20734) );
  OAI21XL U29033 ( .A0(n20958), .A1(n20848), .B0(n20850), .Y(n20818) );
  CMPR32X1 U29034 ( .A(n20813), .B(n20812), .C(U2_A_r_d[7]), .CO(n20814), .S(
        n20754) );
  INVXL U29035 ( .A(n20851), .Y(n20816) );
  OAI21XL U29036 ( .A0(n21008), .A1(n20860), .B0(n20862), .Y(n20824) );
  CMPR22X1 U29037 ( .A(U1_pipe2[9]), .B(n28733), .CO(n20821), .S(n20807) );
  NAND2XL U29038 ( .A(n20822), .B(n20861), .Y(n20823) );
  OAI21XL U29039 ( .A0(n20829), .A1(n20828), .B0(n20827), .Y(n20925) );
  OAI21XL U29040 ( .A0(n20927), .A1(n20831), .B0(n20830), .Y(n20872) );
  CMPR22X1 U29041 ( .A(U1_pipe1[9]), .B(U1_pipe0[9]), .CO(n20833), .S(n20774)
         );
  OAI21XL U29042 ( .A0(n20973), .A1(n20879), .B0(n20881), .Y(n20840) );
  CMPR22X1 U29043 ( .A(U1_pipe12[9]), .B(n28737), .CO(n20837), .S(n20791) );
  OAI21XL U29044 ( .A0(n20986), .A1(n20889), .B0(n20891), .Y(n20846) );
  CMPR22X1 U29045 ( .A(U1_pipe8[9]), .B(n28729), .CO(n20843), .S(n20769) );
  NOR2XL U29046 ( .A(n20848), .B(n20851), .Y(n20951) );
  OAI21XL U29047 ( .A0(n20851), .A1(n20850), .B0(n20849), .Y(n20956) );
  INVXL U29048 ( .A(n20956), .Y(n20852) );
  CMPR32X1 U29049 ( .A(n20855), .B(n20854), .C(U2_A_r_d[8]), .CO(n20856), .S(
        n20815) );
  NOR2XL U29050 ( .A(n20857), .B(n20856), .Y(n20950) );
  NAND2XL U29051 ( .A(n20857), .B(n20856), .Y(n20953) );
  NAND2XL U29052 ( .A(n20900), .B(n20953), .Y(n20858) );
  OAI21XL U29053 ( .A0(n20863), .A1(n20862), .B0(n20861), .Y(n21006) );
  OAI21XL U29054 ( .A0(n21008), .A1(n20865), .B0(n20864), .Y(n20912) );
  CMPR22X1 U29055 ( .A(U1_pipe2[10]), .B(n28851), .CO(n20867), .S(n20820) );
  CMPR22X1 U29056 ( .A(U1_pipe1[10]), .B(U1_pipe0[10]), .CO(n20874), .S(n20832) );
  OAI21XL U29057 ( .A0(n20882), .A1(n20881), .B0(n20880), .Y(n20971) );
  OAI21XL U29058 ( .A0(n20973), .A1(n20884), .B0(n20883), .Y(n20934) );
  CMPR22X1 U29059 ( .A(U1_pipe12[10]), .B(n28867), .CO(n20886), .S(n20836) );
  OAI21XL U29060 ( .A0(n20892), .A1(n20891), .B0(n20890), .Y(n20984) );
  OAI21XL U29061 ( .A0(n20986), .A1(n20894), .B0(n20893), .Y(n20943) );
  CMPR22X1 U29062 ( .A(U1_pipe8[10]), .B(n28835), .CO(n20896), .S(n20842) );
  INVX1 U29063 ( .A(n26291), .Y(n20960) );
  NAND2XL U29064 ( .A(n20905), .B(n20904), .Y(n20952) );
  CMPR22X1 U29065 ( .A(U1_pipe2[11]), .B(n28850), .CO(n20914), .S(n20866) );
  OAI21XL U29066 ( .A0(n20923), .A1(n20922), .B0(n20921), .Y(n20924) );
  OAI21XL U29067 ( .A0(n20927), .A1(n21149), .B0(n21158), .Y(n20993) );
  CMPR22X1 U29068 ( .A(U1_pipe1[11]), .B(U1_pipe0[11]), .CO(n20929), .S(n20873) );
  NAND2XL U29069 ( .A(n20992), .B(n21045), .Y(n20930) );
  CMPR22X1 U29070 ( .A(U1_pipe12[11]), .B(n28866), .CO(n20936), .S(n20885) );
  CMPR22X1 U29071 ( .A(U1_pipe8[11]), .B(n28834), .CO(n20945), .S(n20895) );
  NOR2XL U29072 ( .A(n20950), .B(n20954), .Y(n20957) );
  NAND2XL U29073 ( .A(n20951), .B(n20957), .Y(n21177) );
  OAI21XL U29074 ( .A0(n20954), .A1(n20953), .B0(n20952), .Y(n20955) );
  OAI21XL U29075 ( .A0(n20958), .A1(n21177), .B0(n21186), .Y(n21015) );
  INVXL U29076 ( .A(n21015), .Y(n21069) );
  NAND2XL U29077 ( .A(n21014), .B(n21065), .Y(n20963) );
  OAI21XL U29078 ( .A0(n20969), .A1(n20968), .B0(n20967), .Y(n20970) );
  OAI21XL U29079 ( .A0(n20973), .A1(n21198), .B0(n21207), .Y(n21027) );
  CMPR22X1 U29080 ( .A(U1_pipe12[12]), .B(n28865), .CO(n20975), .S(n20935) );
  OAI21XL U29081 ( .A0(n20982), .A1(n20981), .B0(n20980), .Y(n20983) );
  OAI21XL U29082 ( .A0(n20986), .A1(n21246), .B0(n21255), .Y(n21036) );
  CMPR22X1 U29083 ( .A(U1_pipe8[12]), .B(n28833), .CO(n20988), .S(n20944) );
  CMPR22X1 U29084 ( .A(U1_pipe1[12]), .B(U1_pipe0[12]), .CO(n20995), .S(n20928) );
  OAI21XL U29085 ( .A0(n21004), .A1(n21003), .B0(n21002), .Y(n21005) );
  OAI21XL U29086 ( .A0(n21008), .A1(n21218), .B0(n21227), .Y(n21056) );
  CMPR22X1 U29087 ( .A(U1_pipe2[12]), .B(n28849), .CO(n21010), .S(n20913) );
  INVXL U29088 ( .A(n21065), .Y(n21013) );
  CMPR22X1 U29089 ( .A(U1_pipe12[13]), .B(n28864), .CO(n21029), .S(n20974) );
  CMPR22X1 U29090 ( .A(U1_pipe8[13]), .B(n28832), .CO(n21038), .S(n20987) );
  OAI21XL U29091 ( .A0(n21046), .A1(n21045), .B0(n21044), .Y(n21154) );
  OAI21XL U29092 ( .A0(n21049), .A1(n21048), .B0(n21047), .Y(n21100) );
  CMPR22X1 U29093 ( .A(U1_pipe1[13]), .B(U1_pipe0[13]), .CO(n21051), .S(n20994) );
  CMPR22X1 U29094 ( .A(U1_pipe2[13]), .B(n28848), .CO(n21058), .S(n21009) );
  OAI21XL U29095 ( .A0(n21066), .A1(n21065), .B0(n21064), .Y(n21182) );
  OAI21XL U29096 ( .A0(n21069), .A1(n21068), .B0(n21067), .Y(n21120) );
  ADDHX2 U29097 ( .A(U2_U0_y1[26]), .B(U2_U0_y0[26]), .CO(n26460), .S(n26404)
         );
  CLKINVX3 U29098 ( .A(n26460), .Y(n21121) );
  OAI21XL U29099 ( .A0(n21079), .A1(n21078), .B0(n21077), .Y(n21203) );
  OAI21XL U29100 ( .A0(n21082), .A1(n21081), .B0(n21080), .Y(n21131) );
  CMPR22X1 U29101 ( .A(U1_pipe12[14]), .B(n28863), .CO(n21084), .S(n21028) );
  OAI21XL U29102 ( .A0(n21090), .A1(n21089), .B0(n21088), .Y(n21251) );
  OAI21XL U29103 ( .A0(n21093), .A1(n21092), .B0(n21091), .Y(n21140) );
  CMPR22X1 U29104 ( .A(U1_pipe8[14]), .B(n28831), .CO(n21095), .S(n21037) );
  CMPR22X1 U29105 ( .A(U1_pipe1[14]), .B(U1_pipe0[14]), .CO(n21102), .S(n21050) );
  OAI21XL U29106 ( .A0(n21110), .A1(n21109), .B0(n21108), .Y(n21223) );
  OAI21XL U29107 ( .A0(n21113), .A1(n21112), .B0(n21111), .Y(n21168) );
  CMPR22X1 U29108 ( .A(U1_pipe2[14]), .B(n28847), .CO(n21115), .S(n21057) );
  AOI21XL U29109 ( .A0(n21120), .A1(n21119), .B0(n21118), .Y(n21127) );
  INVXL U29110 ( .A(n21180), .Y(n21125) );
  NAND2XL U29111 ( .A(n21124), .B(n21123), .Y(n21178) );
  XOR2X1 U29112 ( .A(n21127), .B(n21126), .Y(n21128) );
  CMPR22X1 U29113 ( .A(U1_pipe12[15]), .B(n28862), .CO(n21133), .S(n21083) );
  CMPR22X1 U29114 ( .A(U1_pipe8[15]), .B(n28830), .CO(n21142), .S(n21094) );
  OAI21XL U29115 ( .A0(n21152), .A1(n21151), .B0(n21150), .Y(n21153) );
  OAI21XL U29116 ( .A0(n21158), .A1(n21157), .B0(n21156), .Y(n21159) );
  CMPR22X1 U29117 ( .A(U1_pipe1[15]), .B(U1_pipe0[15]), .CO(n21163), .S(n21101) );
  CMPR22X1 U29118 ( .A(U1_pipe2[15]), .B(n28846), .CO(n21170), .S(n21114) );
  NAND2XL U29119 ( .A(n21176), .B(n21183), .Y(n21185) );
  NOR2XL U29120 ( .A(n21177), .B(n21185), .Y(n21188) );
  OAI21XL U29121 ( .A0(n21180), .A1(n21179), .B0(n21178), .Y(n21181) );
  AOI21XL U29122 ( .A0(n21183), .A1(n21182), .B0(n21181), .Y(n21184) );
  OAI21XL U29123 ( .A0(n21186), .A1(n21185), .B0(n21184), .Y(n21187) );
  INVX1 U29124 ( .A(n26607), .Y(n21266) );
  NOR2XL U29125 ( .A(n21193), .B(n21192), .Y(n21304) );
  NAND2XL U29126 ( .A(n21265), .B(n21306), .Y(n21194) );
  OAI21XL U29127 ( .A0(n21201), .A1(n21200), .B0(n21199), .Y(n21202) );
  OAI21XL U29128 ( .A0(n21207), .A1(n21206), .B0(n21205), .Y(n21208) );
  OAI21XL U29129 ( .A0(n21221), .A1(n21220), .B0(n21219), .Y(n21222) );
  OAI21XL U29130 ( .A0(n21227), .A1(n21226), .B0(n21225), .Y(n21228) );
  CMPR22X1 U29131 ( .A(U1_pipe1[16]), .B(U1_pipe0[16]), .CO(n21239), .S(n21162) );
  OAI21XL U29132 ( .A0(n21249), .A1(n21248), .B0(n21247), .Y(n21250) );
  OAI21XL U29133 ( .A0(n21255), .A1(n21254), .B0(n21253), .Y(n21256) );
  INVXL U29134 ( .A(n21306), .Y(n21264) );
  AOI21XL U29135 ( .A0(n21528), .A1(n21265), .B0(n21264), .Y(n21271) );
  INVX1 U29136 ( .A(n26645), .Y(n21308) );
  CMPR32X1 U29137 ( .A(n21266), .B(n7560), .C(U2_A_r_d[15]), .CO(n21267), .S(
        n21193) );
  NAND2XL U29138 ( .A(n21269), .B(n21305), .Y(n21270) );
  OAI21XL U29139 ( .A0(n21290), .A1(n21289), .B0(n21288), .Y(n21340) );
  NOR2XL U29140 ( .A(n21304), .B(n21307), .Y(n21414) );
  OAI21X1 U29141 ( .A0(n21307), .A1(n21306), .B0(n21305), .Y(n21419) );
  AOI21XL U29142 ( .A0(n21528), .A1(n21414), .B0(n21419), .Y(n21360) );
  INVX1 U29143 ( .A(n26703), .Y(n21362) );
  CLKINVX2 U29144 ( .A(n26702), .Y(n21361) );
  NOR2X1 U29145 ( .A(n21311), .B(n21310), .Y(n21413) );
  CMPR22X1 U29146 ( .A(U1_pipe12[18]), .B(n28859), .CO(n21321), .S(n21275) );
  CMPR22X1 U29147 ( .A(U1_pipe2[18]), .B(n28843), .CO(n21332), .S(n21299) );
  CMPR22X1 U29148 ( .A(U1_pipe1[18]), .B(U1_pipe0[18]), .CO(n21344), .S(n21292) );
  CMPR22X1 U29149 ( .A(U1_pipe8[18]), .B(n28827), .CO(n21355), .S(n21282) );
  OAI21XL U29150 ( .A0(n21360), .A1(n21413), .B0(n21416), .Y(n21367) );
  INVX1 U29151 ( .A(n26760), .Y(n21424) );
  NOR2X2 U29152 ( .A(n21364), .B(n21363), .Y(n21417) );
  NAND2X1 U29153 ( .A(n21364), .B(n21363), .Y(n21415) );
  OAI21XL U29154 ( .A0(n21372), .A1(n21371), .B0(n21370), .Y(n21432) );
  OAI21XL U29155 ( .A0(n21383), .A1(n21382), .B0(n21381), .Y(n21444) );
  OAI21XL U29156 ( .A0(n21394), .A1(n21393), .B0(n21392), .Y(n21456) );
  OAI21XL U29157 ( .A0(n21405), .A1(n21404), .B0(n21403), .Y(n21468) );
  NAND2X1 U29158 ( .A(n21414), .B(n21420), .Y(n21519) );
  INVXL U29159 ( .A(n21519), .Y(n21422) );
  OAI21XL U29160 ( .A0(n21417), .A1(n21416), .B0(n21415), .Y(n21418) );
  AOI21X1 U29161 ( .A0(n21420), .A1(n21419), .B0(n21418), .Y(n21527) );
  AOI21XL U29162 ( .A0(n21528), .A1(n21422), .B0(n21421), .Y(n21478) );
  NOR2X1 U29163 ( .A(n21426), .B(n21425), .Y(n21477) );
  INVXL U29164 ( .A(n21477), .Y(n21518) );
  OAI21XL U29165 ( .A0(n21435), .A1(n21434), .B0(n21433), .Y(n21488) );
  OAI21XL U29166 ( .A0(n21447), .A1(n21446), .B0(n21445), .Y(n21512) );
  OAI21XL U29167 ( .A0(n21459), .A1(n21458), .B0(n21457), .Y(n21504) );
  OAI21XL U29168 ( .A0(n21471), .A1(n21470), .B0(n21469), .Y(n21496) );
  OAI21XL U29169 ( .A0(n21478), .A1(n21477), .B0(n21520), .Y(n21484) );
  NAND2XL U29170 ( .A(n21482), .B(n21481), .Y(n21521) );
  CMPR22X1 U29171 ( .A(U1_pipe12[21]), .B(n28856), .CO(n21490), .S(n21437) );
  CMPR22X1 U29172 ( .A(U1_pipe8[21]), .B(n28824), .CO(n21498), .S(n21473) );
  CMPR22X1 U29173 ( .A(U1_pipe1[21]), .B(U1_pipe0[21]), .CO(n21506), .S(n21461) );
  CMPR22X1 U29174 ( .A(U1_pipe2[21]), .B(n28840), .CO(n21514), .S(n21449) );
  NOR2X1 U29175 ( .A(n21519), .B(n21526), .Y(n21568) );
  INVXL U29176 ( .A(n21520), .Y(n21523) );
  INVXL U29177 ( .A(n21521), .Y(n21522) );
  AOI21X1 U29178 ( .A0(n21524), .A1(n21523), .B0(n21522), .Y(n21525) );
  OAI21X1 U29179 ( .A0(n21527), .A1(n21526), .B0(n21525), .Y(n21571) );
  AOI21XL U29180 ( .A0(n21528), .A1(n21568), .B0(n21571), .Y(n21534) );
  NAND2XL U29181 ( .A(n21532), .B(n21531), .Y(n21569) );
  OAI21XL U29182 ( .A0(n21538), .A1(n21537), .B0(n21536), .Y(n21582) );
  OAI21XL U29183 ( .A0(n21546), .A1(n21545), .B0(n21544), .Y(n21590) );
  OAI21XL U29184 ( .A0(n21554), .A1(n21553), .B0(n21552), .Y(n21598) );
  OAI21XL U29185 ( .A0(n21562), .A1(n21561), .B0(n21560), .Y(n21606) );
  INVXL U29186 ( .A(n21569), .Y(n21570) );
  INVXL U29187 ( .A(n26949), .Y(n21616) );
  CMPR22X1 U29188 ( .A(U1_pipe12[23]), .B(n28949), .CO(n21584), .S(n21540) );
  CMPR22X1 U29189 ( .A(U1_pipe8[23]), .B(n28941), .CO(n21592), .S(n21548) );
  CMPR22X1 U29190 ( .A(U1_pipe1[23]), .B(U1_pipe0[23]), .CO(n21600), .S(n21556) );
  CMPR22X1 U29191 ( .A(U1_pipe2[23]), .B(n28945), .CO(n21608), .S(n21564) );
  NOR2X1 U29192 ( .A(n21618), .B(n21617), .Y(n21657) );
  OAI21XL U29193 ( .A0(n21624), .A1(n21623), .B0(n21622), .Y(n21662) );
  OAI21XL U29194 ( .A0(n21632), .A1(n21631), .B0(n21630), .Y(n21670) );
  OAI21XL U29195 ( .A0(n21640), .A1(n21639), .B0(n21638), .Y(n21678) );
  OAI21XL U29196 ( .A0(n21648), .A1(n21647), .B0(n21646), .Y(n21686) );
  CMPR22X1 U29197 ( .A(U2_U0_y1[37]), .B(U2_U0_y0[37]), .CO(n27032), .S(n26991) );
  CMPR32X1 U29198 ( .A(n21655), .B(n21654), .C(U2_A_r_d[23]), .CO(n21692), .S(
        n21618) );
  CMPR22X1 U29199 ( .A(U1_pipe12[25]), .B(n28947), .CO(n21664), .S(n21626) );
  CMPR22X1 U29200 ( .A(U1_pipe2[25]), .B(n28943), .CO(n21672), .S(n21634) );
  CMPR22X1 U29201 ( .A(U1_pipe1[25]), .B(U1_pipe0[25]), .CO(n21680), .S(n21642) );
  CMPR22X1 U29202 ( .A(U1_pipe8[25]), .B(n28939), .CO(n21688), .S(n21650) );
  CMPR22X1 U29203 ( .A(U2_U0_y1[38]), .B(U2_U0_y0[38]), .CO(n21694), .S(n27033) );
  XOR3X2 U29204 ( .A(n5785), .B(n21695), .C(U2_A_r_d[25]), .Y(n27035) );
  CMPR32X1 U29205 ( .A(n21697), .B(n21696), .C(U2_A_r_d[24]), .CO(n21698), .S(
        n21693) );
  MXI2X1 U29206 ( .A(U2_pipe2[25]), .B(n21701), .S0(n21700), .Y(n4197) );
  CMPR22X1 U29207 ( .A(U1_pipe12[26]), .B(n29005), .CO(n21706), .S(n21663) );
  OAI21XL U29208 ( .A0(n21704), .A1(n21703), .B0(n21702), .Y(n21705) );
  CMPR32X1 U29209 ( .A(n21707), .B(n21706), .C(n21705), .S(n21708) );
  CMPR22X1 U29210 ( .A(U1_pipe2[26]), .B(n29004), .CO(n21713), .S(n21671) );
  OAI21XL U29211 ( .A0(n21711), .A1(n21710), .B0(n21709), .Y(n21712) );
  CMPR32X1 U29212 ( .A(n21714), .B(n21713), .C(n21712), .S(n21715) );
  CMPR22X1 U29213 ( .A(U1_pipe1[26]), .B(U1_pipe0[26]), .CO(n21720), .S(n21679) );
  OAI21XL U29214 ( .A0(n21718), .A1(n21717), .B0(n21716), .Y(n21719) );
  CMPR32X1 U29215 ( .A(n21721), .B(n21720), .C(n21719), .S(n21722) );
  CMPR22X1 U29216 ( .A(U1_pipe8[26]), .B(n29003), .CO(n21727), .S(n21687) );
  OAI21XL U29217 ( .A0(n21725), .A1(n21724), .B0(n21723), .Y(n21726) );
  CMPR32X1 U29218 ( .A(n21728), .B(n21727), .C(n21726), .S(n21729) );
  CLKINVX3 U29219 ( .A(n28998), .Y(n23695) );
  NOR2XL U29220 ( .A(n21748), .B(U2_A_i_d[6]), .Y(n21750) );
  NOR2XL U29221 ( .A(n21747), .B(U2_A_i_d[5]), .Y(n21916) );
  OR2X2 U29222 ( .A(n21751), .B(U2_A_i_d[7]), .Y(n21753) );
  NAND2XL U29223 ( .A(n21912), .B(n21753), .Y(n21755) );
  NOR2XL U29224 ( .A(n14338), .B(U2_A_i_d[4]), .Y(n21744) );
  NOR2XL U29225 ( .A(n21742), .B(U2_A_i_d[3]), .Y(n21929) );
  NOR2XL U29226 ( .A(n21744), .B(n21929), .Y(n21746) );
  NOR2XL U29227 ( .A(n25285), .B(U2_A_i_d[0]), .Y(n21943) );
  INVXL U29228 ( .A(n21943), .Y(n21738) );
  NOR2XL U29229 ( .A(n21735), .B(U2_A_i_d[1]), .Y(n21734) );
  INVXL U29230 ( .A(n21734), .Y(n21737) );
  AOI21XL U29231 ( .A0(n21738), .A1(n21737), .B0(n21736), .Y(n21939) );
  NOR2XL U29232 ( .A(n21739), .B(U2_A_i_d[2]), .Y(n21741) );
  OAI21XL U29233 ( .A0(n21939), .A1(n21741), .B0(n21740), .Y(n21927) );
  NAND2XL U29234 ( .A(n21742), .B(U2_A_i_d[3]), .Y(n21928) );
  NAND2XL U29235 ( .A(n14338), .B(U2_A_i_d[4]), .Y(n21743) );
  OAI21XL U29236 ( .A0(n21744), .A1(n21928), .B0(n21743), .Y(n21745) );
  AOI21XL U29237 ( .A0(n21746), .A1(n21927), .B0(n21745), .Y(n21910) );
  NAND2XL U29238 ( .A(n21747), .B(U2_A_i_d[5]), .Y(n21917) );
  NAND2XL U29239 ( .A(n21748), .B(U2_A_i_d[6]), .Y(n21749) );
  OAI21XL U29240 ( .A0(n21750), .A1(n21917), .B0(n21749), .Y(n21911) );
  NOR2XL U29241 ( .A(n5871), .B(U2_A_i_d[10]), .Y(n21760) );
  NOR2XL U29242 ( .A(n14380), .B(U2_A_i_d[9]), .Y(n21896) );
  NOR2XL U29243 ( .A(n21758), .B(U2_A_i_d[8]), .Y(n21895) );
  INVXL U29244 ( .A(n21895), .Y(n21756) );
  NAND2XL U29245 ( .A(n21763), .B(n21756), .Y(n21883) );
  NOR2XL U29246 ( .A(n21764), .B(U2_A_i_d[12]), .Y(n21757) );
  INVXL U29247 ( .A(n21757), .Y(n21766) );
  OR2XL U29248 ( .A(n14386), .B(U2_A_i_d[11]), .Y(n21885) );
  NAND2XL U29249 ( .A(n21766), .B(n21885), .Y(n21768) );
  NOR2XL U29250 ( .A(n21883), .B(n21768), .Y(n21770) );
  NAND2XL U29251 ( .A(n21758), .B(U2_A_i_d[8]), .Y(n21894) );
  INVXL U29252 ( .A(n21894), .Y(n21762) );
  NAND2XL U29253 ( .A(n14380), .B(U2_A_i_d[9]), .Y(n21897) );
  NAND2XL U29254 ( .A(n5871), .B(U2_A_i_d[10]), .Y(n21759) );
  OAI21XL U29255 ( .A0(n21760), .A1(n21897), .B0(n21759), .Y(n21761) );
  AOI21XL U29256 ( .A0(n21763), .A1(n21762), .B0(n21761), .Y(n21882) );
  AOI21XL U29257 ( .A0(n21766), .A1(n21884), .B0(n21765), .Y(n21767) );
  OAI21XL U29258 ( .A0(n21882), .A1(n21768), .B0(n21767), .Y(n21769) );
  NOR2XL U29259 ( .A(n14445), .B(U2_A_i_d[16]), .Y(n21771) );
  INVXL U29260 ( .A(n21771), .Y(n21778) );
  NOR2XL U29261 ( .A(n14444), .B(U2_A_i_d[15]), .Y(n21865) );
  INVXL U29262 ( .A(n21865), .Y(n21772) );
  NAND2XL U29263 ( .A(n21778), .B(n21772), .Y(n21780) );
  INVXL U29264 ( .A(n25203), .Y(n21773) );
  OR2X2 U29265 ( .A(n21773), .B(U2_A_i_d[13]), .Y(n21874) );
  NAND2XL U29266 ( .A(n8058), .B(n21874), .Y(n21860) );
  NOR2XL U29267 ( .A(n21780), .B(n21860), .Y(n21841) );
  OR2X2 U29268 ( .A(n21784), .B(U2_A_i_d[20]), .Y(n21786) );
  OR2X2 U29269 ( .A(n14453), .B(U2_A_i_d[19]), .Y(n21845) );
  NAND2X1 U29270 ( .A(n21786), .B(n21845), .Y(n21788) );
  OR2X2 U29271 ( .A(n5863), .B(U2_A_i_d[17]), .Y(n21853) );
  NAND2X1 U29272 ( .A(n21783), .B(n21853), .Y(n21843) );
  NOR2XL U29273 ( .A(n21788), .B(n21843), .Y(n21790) );
  NAND2XL U29274 ( .A(n21841), .B(n21790), .Y(n21792) );
  AND2X2 U29275 ( .A(n21773), .B(U2_A_i_d[13]), .Y(n21873) );
  AOI21XL U29276 ( .A0(n8058), .A1(n21873), .B0(n21775), .Y(n21861) );
  NAND2XL U29277 ( .A(n14444), .B(U2_A_i_d[15]), .Y(n21864) );
  INVXL U29278 ( .A(n21864), .Y(n21777) );
  AOI21XL U29279 ( .A0(n21778), .A1(n21777), .B0(n21776), .Y(n21779) );
  OAI21XL U29280 ( .A0(n21780), .A1(n21861), .B0(n21779), .Y(n21840) );
  AND2X2 U29281 ( .A(n21781), .B(U2_A_i_d[18]), .Y(n21782) );
  AOI21X1 U29282 ( .A0(n21783), .A1(n21852), .B0(n21782), .Y(n21842) );
  AND2X2 U29283 ( .A(n14453), .B(U2_A_i_d[19]), .Y(n21844) );
  AOI21XL U29284 ( .A0(n21786), .A1(n21844), .B0(n21785), .Y(n21787) );
  OAI21XL U29285 ( .A0(n21788), .A1(n21842), .B0(n21787), .Y(n21789) );
  AOI21X1 U29286 ( .A0(n21840), .A1(n21790), .B0(n21789), .Y(n21791) );
  OAI21X1 U29287 ( .A0(n21839), .A1(n21792), .B0(n21791), .Y(n21815) );
  NOR2XL U29288 ( .A(n21794), .B(U2_A_i_d[21]), .Y(n21831) );
  INVXL U29289 ( .A(n25147), .Y(n21795) );
  NOR2XL U29290 ( .A(n21795), .B(U2_A_i_d[22]), .Y(n21797) );
  NOR2XL U29291 ( .A(n21831), .B(n21797), .Y(n21822) );
  NOR2XL U29292 ( .A(n14484), .B(U2_A_i_d[23]), .Y(n21793) );
  INVXL U29293 ( .A(n21793), .Y(n21799) );
  NAND2XL U29294 ( .A(n21822), .B(n21799), .Y(n21817) );
  NOR2XL U29295 ( .A(n21800), .B(U2_A_i_d[24]), .Y(n21802) );
  NOR2XL U29296 ( .A(n21817), .B(n21802), .Y(n21804) );
  NAND2XL U29297 ( .A(n21794), .B(U2_A_i_d[21]), .Y(n21830) );
  NAND2XL U29298 ( .A(n21795), .B(U2_A_i_d[22]), .Y(n21796) );
  NAND2XL U29299 ( .A(n21800), .B(U2_A_i_d[24]), .Y(n21801) );
  OAI21XL U29300 ( .A0(n21816), .A1(n21802), .B0(n21801), .Y(n21803) );
  AOI21X1 U29301 ( .A0(n21815), .A1(n21804), .B0(n21803), .Y(n21813) );
  NOR2XL U29302 ( .A(n21805), .B(U2_A_i_d[25]), .Y(n21807) );
  NAND2XL U29303 ( .A(n21805), .B(U2_A_i_d[25]), .Y(n21806) );
  INVX1 U29304 ( .A(n21808), .Y(n21809) );
  MXI2X1 U29305 ( .A(U0_pipe6[27]), .B(n21809), .S0(n20438), .Y(n4463) );
  OR2X2 U29306 ( .A(n25125), .B(U2_A_i_d[25]), .Y(n22177) );
  NAND2X1 U29307 ( .A(n25125), .B(U2_A_i_d[25]), .Y(n22176) );
  NAND2X1 U29308 ( .A(n22177), .B(n22176), .Y(n22181) );
  XOR2X1 U29309 ( .A(n21813), .B(n21812), .Y(n21814) );
  OAI21XL U29310 ( .A0(n21837), .A1(n21817), .B0(n21816), .Y(n21820) );
  XNOR2X1 U29311 ( .A(n21820), .B(n21819), .Y(n21821) );
  INVXL U29312 ( .A(n21823), .Y(n21824) );
  OAI21XL U29313 ( .A0(n21837), .A1(n21825), .B0(n21824), .Y(n21828) );
  NOR2XL U29314 ( .A(n25140), .B(U2_A_i_d[23]), .Y(n22171) );
  INVXL U29315 ( .A(n22171), .Y(n21826) );
  XNOR2X1 U29316 ( .A(n21828), .B(n21827), .Y(n21829) );
  OAI21XL U29317 ( .A0(n21837), .A1(n21831), .B0(n21830), .Y(n21834) );
  NOR2XL U29318 ( .A(n25147), .B(U2_A_i_d[22]), .Y(n21832) );
  NAND2XL U29319 ( .A(n25147), .B(U2_A_i_d[22]), .Y(n22166) );
  XNOR2X1 U29320 ( .A(n21834), .B(n21833), .Y(n21835) );
  NOR2XL U29321 ( .A(n25151), .B(U2_A_i_d[21]), .Y(n22192) );
  INVXL U29322 ( .A(n22192), .Y(n22165) );
  NAND2XL U29323 ( .A(n25151), .B(U2_A_i_d[21]), .Y(n22191) );
  OAI21X1 U29324 ( .A0(n21851), .A1(n21843), .B0(n21842), .Y(n21849) );
  NAND2XL U29325 ( .A(n25162), .B(U2_A_i_d[20]), .Y(n22156) );
  XOR2X1 U29326 ( .A(n21846), .B(n22206), .Y(n21847) );
  INVXL U29327 ( .A(n22205), .Y(n22141) );
  NAND2XL U29328 ( .A(n25166), .B(U2_A_i_d[19]), .Y(n22204) );
  NAND2XL U29329 ( .A(n22141), .B(n22204), .Y(n22207) );
  AOI21XL U29330 ( .A0(n21858), .A1(n21853), .B0(n21852), .Y(n21855) );
  OR2X2 U29331 ( .A(n25174), .B(U2_A_i_d[18]), .Y(n22155) );
  NAND2XL U29332 ( .A(n25174), .B(U2_A_i_d[18]), .Y(n22152) );
  NOR2XL U29333 ( .A(n25178), .B(U2_A_i_d[17]), .Y(n22211) );
  INVXL U29334 ( .A(n22211), .Y(n22142) );
  NAND2XL U29335 ( .A(n25178), .B(U2_A_i_d[17]), .Y(n22210) );
  NAND2XL U29336 ( .A(n22142), .B(n22210), .Y(n22216) );
  OAI21XL U29337 ( .A0(n21871), .A1(n21865), .B0(n21864), .Y(n21868) );
  NOR2XL U29338 ( .A(n25189), .B(U2_A_i_d[16]), .Y(n21866) );
  INVXL U29339 ( .A(n21866), .Y(n22149) );
  NAND2XL U29340 ( .A(n25189), .B(U2_A_i_d[16]), .Y(n22146) );
  NOR2XL U29341 ( .A(n25193), .B(U2_A_i_d[15]), .Y(n22223) );
  INVXL U29342 ( .A(n22223), .Y(n22140) );
  NAND2XL U29343 ( .A(n25193), .B(U2_A_i_d[15]), .Y(n22222) );
  AOI21XL U29344 ( .A0(n21879), .A1(n21874), .B0(n21873), .Y(n21876) );
  NAND2XL U29345 ( .A(n25199), .B(U2_A_i_d[14]), .Y(n22144) );
  OR2X1 U29346 ( .A(n25203), .B(U2_A_i_d[13]), .Y(n22231) );
  NAND2XL U29347 ( .A(n25203), .B(U2_A_i_d[13]), .Y(n22143) );
  OAI21XL U29348 ( .A0(n21908), .A1(n21883), .B0(n21882), .Y(n21892) );
  NAND2XL U29349 ( .A(n25212), .B(U2_A_i_d[12]), .Y(n22114) );
  NOR2XL U29350 ( .A(n25216), .B(U2_A_i_d[11]), .Y(n21890) );
  INVXL U29351 ( .A(n21890), .Y(n22242) );
  NAND2XL U29352 ( .A(n25216), .B(U2_A_i_d[11]), .Y(n22113) );
  OAI21XL U29353 ( .A0(n21908), .A1(n21895), .B0(n21894), .Y(n21905) );
  INVXL U29354 ( .A(n21896), .Y(n21899) );
  INVXL U29355 ( .A(n22110), .Y(n21900) );
  NAND2XL U29356 ( .A(n25226), .B(U2_A_i_d[10]), .Y(n22109) );
  NOR2XL U29357 ( .A(n25231), .B(U2_A_i_d[9]), .Y(n22108) );
  NAND2XL U29358 ( .A(n25231), .B(U2_A_i_d[9]), .Y(n22252) );
  NOR2XL U29359 ( .A(n25235), .B(U2_A_i_d[8]), .Y(n22251) );
  INVXL U29360 ( .A(n22251), .Y(n22118) );
  NAND2XL U29361 ( .A(n25235), .B(U2_A_i_d[8]), .Y(n22250) );
  AOI21XL U29362 ( .A0(n21925), .A1(n21912), .B0(n21911), .Y(n21914) );
  OR2X2 U29363 ( .A(n25243), .B(U2_A_i_d[7]), .Y(n22134) );
  NAND2XL U29364 ( .A(n25243), .B(U2_A_i_d[7]), .Y(n22132) );
  NOR2XL U29365 ( .A(n25251), .B(U2_A_i_d[6]), .Y(n22131) );
  INVXL U29366 ( .A(n22131), .Y(n21920) );
  NAND2XL U29367 ( .A(n25251), .B(U2_A_i_d[6]), .Y(n22130) );
  NOR2XL U29368 ( .A(n25256), .B(U2_A_i_d[5]), .Y(n22121) );
  NAND2XL U29369 ( .A(n25256), .B(U2_A_i_d[5]), .Y(n22270) );
  OAI21XL U29370 ( .A0(n21936), .A1(n21929), .B0(n21928), .Y(n21932) );
  NOR2XL U29371 ( .A(n25263), .B(U2_A_i_d[4]), .Y(n22127) );
  NAND2XL U29372 ( .A(n25263), .B(U2_A_i_d[4]), .Y(n22126) );
  NOR2XL U29373 ( .A(n25269), .B(U2_A_i_d[3]), .Y(n22281) );
  NAND2XL U29374 ( .A(n25269), .B(U2_A_i_d[3]), .Y(n22280) );
  NOR2XL U29375 ( .A(n25275), .B(U2_A_i_d[2]), .Y(n22125) );
  NAND2XL U29376 ( .A(n25275), .B(U2_A_i_d[2]), .Y(n22124) );
  XOR2XL U29377 ( .A(n21940), .B(n21939), .Y(n21941) );
  NAND2XL U29378 ( .A(n25281), .B(U2_A_i_d[1]), .Y(n22122) );
  XOR2XL U29379 ( .A(n21944), .B(n21943), .Y(n21945) );
  XNOR2XL U29380 ( .A(n25285), .B(U2_A_i_d[0]), .Y(n22294) );
  MXI2X1 U29381 ( .A(U0_pipe7[26]), .B(n21947), .S0(n22248), .Y(n4436) );
  XOR2X1 U29382 ( .A(n21950), .B(n22298), .Y(n21951) );
  INVXL U29383 ( .A(n21958), .Y(n21959) );
  OAI21XL U29384 ( .A0(n21976), .A1(n21960), .B0(n21959), .Y(n21965) );
  INVXL U29385 ( .A(n21961), .Y(n21963) );
  XNOR2X1 U29386 ( .A(n21965), .B(n21964), .Y(n21966) );
  OAI21XL U29387 ( .A0(n21976), .A1(n21968), .B0(n21967), .Y(n21971) );
  XNOR2X1 U29388 ( .A(n21971), .B(n21970), .Y(n21973) );
  XOR2X1 U29389 ( .A(n21985), .B(n22324), .Y(n21986) );
  AOI21XL U29390 ( .A0(n21998), .A1(n14552), .B0(n14561), .Y(n21994) );
  INVXL U29391 ( .A(n22000), .Y(n22003) );
  INVXL U29392 ( .A(n22001), .Y(n22002) );
  OAI21XL U29393 ( .A0(n22012), .A1(n22004), .B0(n22009), .Y(n22007) );
  NAND2XL U29394 ( .A(n22010), .B(n22009), .Y(n22011) );
  AOI21XL U29395 ( .A0(n22022), .A1(n14549), .B0(n22014), .Y(n22018) );
  NAND2XL U29396 ( .A(n14549), .B(n22020), .Y(n22021) );
  INVXL U29397 ( .A(n22024), .Y(n22056) );
  OAI21XL U29398 ( .A0(n22056), .A1(n22026), .B0(n22025), .Y(n22036) );
  OAI21XL U29399 ( .A0(n22056), .A1(n22039), .B0(n22038), .Y(n22052) );
  INVXL U29400 ( .A(n22041), .Y(n22042) );
  NAND2XL U29401 ( .A(n22046), .B(n22045), .Y(n22377) );
  NAND2XL U29402 ( .A(n22376), .B(n22374), .Y(n22380) );
  INVXL U29403 ( .A(n22058), .Y(n22076) );
  AOI21XL U29404 ( .A0(n22076), .A1(n22060), .B0(n22059), .Y(n22063) );
  INVXL U29405 ( .A(n22067), .Y(n22069) );
  NAND2XL U29406 ( .A(n22074), .B(n22073), .Y(n22075) );
  OAI21XL U29407 ( .A0(n22089), .A1(n22080), .B0(n22079), .Y(n22085) );
  INVXL U29408 ( .A(n22081), .Y(n22083) );
  INVXL U29409 ( .A(n22408), .Y(n22087) );
  XOR2XL U29410 ( .A(n22095), .B(n22094), .Y(n22096) );
  XOR2XL U29411 ( .A(n22099), .B(n22098), .Y(n22100) );
  XNOR2XL U29412 ( .A(n25449), .B(n22727), .Y(n22424) );
  NAND2XL U29413 ( .A(U0_pipe7[0]), .B(U0_pipe6[0]), .Y(n22102) );
  OAI21XL U29414 ( .A0(n22103), .A1(n22102), .B0(n22101), .Y(n23217) );
  INVXL U29415 ( .A(n22250), .Y(n22112) );
  OAI21XL U29416 ( .A0(n22110), .A1(n22252), .B0(n22109), .Y(n22111) );
  AOI21XL U29417 ( .A0(n22119), .A1(n22112), .B0(n22111), .Y(n22239) );
  INVXL U29418 ( .A(n22113), .Y(n22241) );
  INVXL U29419 ( .A(n22114), .Y(n22115) );
  AOI21XL U29420 ( .A0(n22116), .A1(n22241), .B0(n22115), .Y(n22117) );
  OAI21XL U29421 ( .A0(n22239), .A1(n22120), .B0(n22117), .Y(n22139) );
  NAND2XL U29422 ( .A(n22119), .B(n22118), .Y(n22240) );
  NOR2XL U29423 ( .A(n22240), .B(n22120), .Y(n22137) );
  NOR2XL U29424 ( .A(n22131), .B(n22121), .Y(n22266) );
  NAND2XL U29425 ( .A(n22266), .B(n22134), .Y(n22136) );
  NOR2XL U29426 ( .A(n22127), .B(n22281), .Y(n22129) );
  INVXL U29427 ( .A(n22122), .Y(n22123) );
  AOI21XL U29428 ( .A0(n22291), .A1(n21942), .B0(n22123), .Y(n22288) );
  OAI21XL U29429 ( .A0(n22288), .A1(n22125), .B0(n22124), .Y(n22279) );
  OAI21XL U29430 ( .A0(n22127), .A1(n22280), .B0(n22126), .Y(n22128) );
  AOI21XL U29431 ( .A0(n22129), .A1(n22279), .B0(n22128), .Y(n22264) );
  OAI21XL U29432 ( .A0(n22131), .A1(n22270), .B0(n22130), .Y(n22265) );
  INVXL U29433 ( .A(n22132), .Y(n22133) );
  AOI21X1 U29434 ( .A0(n22265), .A1(n22134), .B0(n22133), .Y(n22135) );
  OAI21XL U29435 ( .A0(n22136), .A1(n22264), .B0(n22135), .Y(n22238) );
  AND2X2 U29436 ( .A(n22137), .B(n22238), .Y(n22138) );
  NAND2XL U29437 ( .A(n22149), .B(n22140), .Y(n22151) );
  NAND2XL U29438 ( .A(n8057), .B(n22231), .Y(n22218) );
  NOR2XL U29439 ( .A(n22151), .B(n22218), .Y(n22200) );
  NAND2X1 U29440 ( .A(n6951), .B(n22141), .Y(n22160) );
  NAND2X1 U29441 ( .A(n22155), .B(n22142), .Y(n22201) );
  NOR2X1 U29442 ( .A(n22160), .B(n22201), .Y(n22162) );
  INVXL U29443 ( .A(n22143), .Y(n22230) );
  INVXL U29444 ( .A(n22144), .Y(n22145) );
  AOI21X1 U29445 ( .A0(n8057), .A1(n22230), .B0(n22145), .Y(n22219) );
  INVXL U29446 ( .A(n22222), .Y(n22148) );
  INVXL U29447 ( .A(n22146), .Y(n22147) );
  AOI21XL U29448 ( .A0(n22149), .A1(n22148), .B0(n22147), .Y(n22150) );
  OAI21XL U29449 ( .A0(n22151), .A1(n22219), .B0(n22150), .Y(n22199) );
  INVXL U29450 ( .A(n22210), .Y(n22154) );
  INVXL U29451 ( .A(n22152), .Y(n22153) );
  AOI21X1 U29452 ( .A0(n22155), .A1(n22154), .B0(n22153), .Y(n22202) );
  INVXL U29453 ( .A(n22204), .Y(n22158) );
  INVXL U29454 ( .A(n22156), .Y(n22157) );
  AOI21X1 U29455 ( .A0(n6951), .A1(n22158), .B0(n22157), .Y(n22159) );
  AOI21X1 U29456 ( .A0(n22199), .A1(n22162), .B0(n22161), .Y(n22163) );
  NAND2XL U29457 ( .A(n22165), .B(n22168), .Y(n22187) );
  INVXL U29458 ( .A(n22191), .Y(n22169) );
  INVXL U29459 ( .A(n22166), .Y(n22167) );
  AOI21X1 U29460 ( .A0(n22169), .A1(n22168), .B0(n22167), .Y(n22186) );
  MXI2X1 U29461 ( .A(U0_pipe4[27]), .B(n22178), .S0(n21972), .Y(n4320) );
  MXI2X1 U29462 ( .A(U0_pipe4[26]), .B(n22179), .S0(n21972), .Y(n4321) );
  MXI2X1 U29463 ( .A(U0_pipe4[25]), .B(n22182), .S0(n21972), .Y(n4322) );
  OAI21XL U29464 ( .A0(n22197), .A1(n22187), .B0(n22186), .Y(n22189) );
  XNOR2XL U29465 ( .A(n22189), .B(n22188), .Y(n22190) );
  OAI21XL U29466 ( .A0(n22197), .A1(n22192), .B0(n22191), .Y(n22194) );
  XNOR2XL U29467 ( .A(n22194), .B(n22193), .Y(n22195) );
  INVXL U29468 ( .A(n22202), .Y(n22203) );
  OAI21XL U29469 ( .A0(n22212), .A1(n22211), .B0(n22210), .Y(n22214) );
  XNOR2XL U29470 ( .A(n22214), .B(n22213), .Y(n22215) );
  CLKINVX3 U29471 ( .A(n5837), .Y(n22543) );
  MXI2X1 U29472 ( .A(U0_pipe4[17]), .B(n22217), .S0(n22543), .Y(n4330) );
  OAI21XL U29473 ( .A0(n22228), .A1(n22223), .B0(n22222), .Y(n22225) );
  XNOR2XL U29474 ( .A(n22225), .B(n22224), .Y(n22226) );
  OAI21XL U29475 ( .A0(n22262), .A1(n22240), .B0(n22239), .Y(n22247) );
  AOI21XL U29476 ( .A0(n22247), .A1(n22242), .B0(n22241), .Y(n22244) );
  OAI21XL U29477 ( .A0(n22262), .A1(n22251), .B0(n22250), .Y(n22259) );
  AOI21XL U29478 ( .A0(n22277), .A1(n22266), .B0(n22265), .Y(n22268) );
  OAI21XL U29479 ( .A0(n22286), .A1(n22281), .B0(n22280), .Y(n22283) );
  XOR2XL U29480 ( .A(n22289), .B(n22288), .Y(n22290) );
  XNOR2XL U29481 ( .A(n22292), .B(n22291), .Y(n22293) );
  MXI2X1 U29482 ( .A(U0_pipe5[27]), .B(n22297), .S0(n22248), .Y(n4491) );
  OAI21XL U29483 ( .A0(n22315), .A1(n22305), .B0(n22304), .Y(n22307) );
  XNOR2XL U29484 ( .A(n22307), .B(n22306), .Y(n22308) );
  OAI21XL U29485 ( .A0(n22315), .A1(n22310), .B0(n22309), .Y(n22312) );
  MXI2X1 U29486 ( .A(U0_pipe5[20]), .B(n22325), .S0(n22248), .Y(n4498) );
  OAI21XL U29487 ( .A0(n22331), .A1(n22330), .B0(n22329), .Y(n22333) );
  XNOR2XL U29488 ( .A(n22333), .B(n22332), .Y(n22334) );
  INVXL U29489 ( .A(n22337), .Y(n22340) );
  AOI21XL U29490 ( .A0(n22359), .A1(n22340), .B0(n22339), .Y(n22349) );
  OAI21XL U29491 ( .A0(n22349), .A1(n22341), .B0(n22346), .Y(n22344) );
  NAND2XL U29492 ( .A(n6988), .B(n22342), .Y(n22343) );
  NAND2XL U29493 ( .A(n22347), .B(n22346), .Y(n22348) );
  AOI21XL U29494 ( .A0(n22359), .A1(n13122), .B0(n22351), .Y(n22355) );
  NAND2XL U29495 ( .A(n13122), .B(n22357), .Y(n22358) );
  INVXL U29496 ( .A(n22361), .Y(n22384) );
  OAI21XL U29497 ( .A0(n22384), .A1(n22363), .B0(n22362), .Y(n22370) );
  OAI21XL U29498 ( .A0(n22384), .A1(n22373), .B0(n22372), .Y(n22381) );
  INVXL U29499 ( .A(n22374), .Y(n22375) );
  AOI21XL U29500 ( .A0(n22381), .A1(n22376), .B0(n22375), .Y(n22378) );
  INVXL U29501 ( .A(n22386), .Y(n22404) );
  AOI21XL U29502 ( .A0(n22404), .A1(n22388), .B0(n22387), .Y(n22391) );
  INVXL U29503 ( .A(n22395), .Y(n22397) );
  OAI21XL U29504 ( .A0(n22416), .A1(n22408), .B0(n22407), .Y(n22413) );
  INVXL U29505 ( .A(n22409), .Y(n22411) );
  XOR2XL U29506 ( .A(n22419), .B(n22418), .Y(n22420) );
  XNOR2XL U29507 ( .A(n22422), .B(n22421), .Y(n22423) );
  NAND2XL U29508 ( .A(U0_pipe5[0]), .B(U0_pipe4[0]), .Y(n22426) );
  OAI21XL U29509 ( .A0(n22427), .A1(n22426), .B0(n22425), .Y(n23199) );
  INVXL U29510 ( .A(n22432), .Y(n22489) );
  NAND2X1 U29511 ( .A(n5796), .B(n22489), .Y(n22440) );
  INVXL U29512 ( .A(n22488), .Y(n22437) );
  INVXL U29513 ( .A(n22435), .Y(n22436) );
  AOI21X1 U29514 ( .A0(n5796), .A1(n22437), .B0(n22436), .Y(n22438) );
  AOI21X1 U29515 ( .A0(n22443), .A1(n22442), .B0(n22441), .Y(n22444) );
  NOR2XL U29516 ( .A(n22448), .B(U2_A_i_d[21]), .Y(n22480) );
  INVXL U29517 ( .A(n22480), .Y(n22485) );
  NAND2XL U29518 ( .A(n22485), .B(n22447), .Y(n22475) );
  NOR2XL U29519 ( .A(n22452), .B(U2_A_i_d[23]), .Y(n22476) );
  NAND2X1 U29520 ( .A(n22448), .B(U2_A_i_d[21]), .Y(n22484) );
  INVXL U29521 ( .A(n22484), .Y(n22451) );
  NAND2XL U29522 ( .A(n22449), .B(U2_A_i_d[22]), .Y(n22481) );
  INVXL U29523 ( .A(n22481), .Y(n22450) );
  AOI21XL U29524 ( .A0(n22451), .A1(n22447), .B0(n22450), .Y(n22474) );
  NOR2X1 U29525 ( .A(n22453), .B(U2_A_i_d[24]), .Y(n22468) );
  OR2X2 U29526 ( .A(n22454), .B(U2_A_i_d[25]), .Y(n22464) );
  OAI21XL U29527 ( .A0(n22461), .A1(n22459), .B0(n22460), .Y(n22457) );
  MXI2X1 U29528 ( .A(U0_pipe14[27]), .B(n22458), .S0(n5805), .Y(n4637) );
  MXI2X1 U29529 ( .A(U0_pipe14[26]), .B(n22462), .S0(n5805), .Y(n4638) );
  XNOR2X1 U29530 ( .A(n22466), .B(n22465), .Y(n22467) );
  MXI2X1 U29531 ( .A(U0_pipe14[25]), .B(n22467), .S0(n5805), .Y(n4639) );
  XOR2X1 U29532 ( .A(n22471), .B(n22747), .Y(n22472) );
  INVXL U29533 ( .A(n22473), .Y(n22486) );
  OAI21XL U29534 ( .A0(n22486), .A1(n22475), .B0(n22474), .Y(n22478) );
  XNOR2X1 U29535 ( .A(n22478), .B(n22755), .Y(n22479) );
  MXI2X1 U29536 ( .A(U0_pipe14[23]), .B(n22479), .S0(n5805), .Y(n4641) );
  OAI21XL U29537 ( .A0(n22486), .A1(n22480), .B0(n22484), .Y(n22482) );
  XNOR2X1 U29538 ( .A(n22482), .B(n22761), .Y(n22483) );
  MXI2X1 U29539 ( .A(U0_pipe14[22]), .B(n22483), .S0(n5805), .Y(n4642) );
  NAND2XL U29540 ( .A(n22485), .B(n22484), .Y(n22765) );
  XOR2X1 U29541 ( .A(n22486), .B(n22765), .Y(n22487) );
  CLKINVX3 U29542 ( .A(n5837), .Y(n25318) );
  NAND2XL U29543 ( .A(n22489), .B(n22488), .Y(n22769) );
  XNOR2XL U29544 ( .A(n22495), .B(n22775), .Y(n22496) );
  NAND2XL U29545 ( .A(n5818), .B(n22497), .Y(n22779) );
  OAI21XL U29546 ( .A0(n22511), .A1(n22504), .B0(n22509), .Y(n22507) );
  XNOR2XL U29547 ( .A(n22507), .B(n22789), .Y(n22508) );
  NAND2XL U29548 ( .A(n22510), .B(n22509), .Y(n22793) );
  OAI21XL U29549 ( .A0(n22547), .A1(n22523), .B0(n22522), .Y(n22530) );
  AOI21XL U29550 ( .A0(n22530), .A1(n14029), .B0(n22524), .Y(n22527) );
  OAI21XL U29551 ( .A0(n22547), .A1(n22532), .B0(n22545), .Y(n22542) );
  INVXL U29552 ( .A(n22533), .Y(n22541) );
  AOI21XL U29553 ( .A0(n22542), .A1(n22541), .B0(n22534), .Y(n22538) );
  AOI21XL U29554 ( .A0(n22567), .A1(n22551), .B0(n22550), .Y(n22554) );
  OAI21XL U29555 ( .A0(n22580), .A1(n22576), .B0(n22577), .Y(n22574) );
  XOR2XL U29556 ( .A(n22586), .B(n22585), .Y(n22587) );
  XNOR2XL U29557 ( .A(n22879), .B(n22589), .Y(n22590) );
  XNOR2XL U29558 ( .A(n24581), .B(U2_A_i_d[0]), .Y(n22883) );
  MXI2X1 U29559 ( .A(U0_pipe15[27]), .B(n5795), .S0(n22620), .Y(n4609) );
  OAI21XL U29560 ( .A0(n22614), .A1(n22601), .B0(n22600), .Y(n22606) );
  OAI21XL U29561 ( .A0(n22614), .A1(n22608), .B0(n22612), .Y(n22610) );
  NAND2XL U29562 ( .A(n22617), .B(n22616), .Y(n22618) );
  OAI21XL U29563 ( .A0(n22623), .A1(n22622), .B0(n22628), .Y(n22626) );
  NAND2XL U29564 ( .A(n6904), .B(n22624), .Y(n22625) );
  NAND2XL U29565 ( .A(n22629), .B(n22628), .Y(n22630) );
  INVXL U29566 ( .A(n22632), .Y(n22635) );
  INVXL U29567 ( .A(n22633), .Y(n22634) );
  OAI21XL U29568 ( .A0(n22645), .A1(n22636), .B0(n22642), .Y(n22640) );
  NAND2XL U29569 ( .A(n22638), .B(n22637), .Y(n22639) );
  NAND2XL U29570 ( .A(n22643), .B(n22642), .Y(n22644) );
  NAND2XL U29571 ( .A(n22649), .B(n22648), .Y(n22650) );
  NAND2XL U29572 ( .A(n12612), .B(n22653), .Y(n22654) );
  OAI21XL U29573 ( .A0(n22685), .A1(n22659), .B0(n22658), .Y(n22667) );
  AOI21XL U29574 ( .A0(n22667), .A1(n12572), .B0(n22660), .Y(n22663) );
  NAND2XL U29575 ( .A(n6997), .B(n22661), .Y(n22662) );
  NAND2XL U29576 ( .A(n12572), .B(n22665), .Y(n22666) );
  OAI21XL U29577 ( .A0(n22685), .A1(n22669), .B0(n22683), .Y(n22681) );
  INVXL U29578 ( .A(n22670), .Y(n22679) );
  INVXL U29579 ( .A(n22678), .Y(n22671) );
  INVXL U29580 ( .A(n22672), .Y(n22674) );
  NAND2XL U29581 ( .A(n22674), .B(n22673), .Y(n22675) );
  NAND2XL U29582 ( .A(n22679), .B(n22678), .Y(n22680) );
  NAND2XL U29583 ( .A(n22684), .B(n22683), .Y(n23079) );
  AOI21XL U29584 ( .A0(n22705), .A1(n22689), .B0(n22688), .Y(n22692) );
  INVXL U29585 ( .A(n22696), .Y(n22698) );
  OAI21XL U29586 ( .A0(n22716), .A1(n22713), .B0(n22714), .Y(n22711) );
  OAI21XL U29587 ( .A0(n22725), .A1(n22718), .B0(n22723), .Y(n22721) );
  XOR2XL U29588 ( .A(n23119), .B(n22725), .Y(n22726) );
  XNOR2XL U29589 ( .A(n22891), .B(n24851), .Y(n23123) );
  CMPR32X1 U29590 ( .A(n24414), .B(n29009), .C(n22735), .CO(n22736), .S(n14159) );
  MXI2X1 U29591 ( .A(U0_pipe10[27]), .B(n22737), .S0(n5812), .Y(n4550) );
  XOR2X1 U29592 ( .A(n22742), .B(n22741), .Y(n22743) );
  OAI21XL U29593 ( .A0(n22767), .A1(n22746), .B0(n22745), .Y(n22749) );
  MXI2X1 U29594 ( .A(U0_pipe10[24]), .B(n22750), .S0(n5812), .Y(n4553) );
  INVXL U29595 ( .A(n22752), .Y(n22753) );
  OAI21XL U29596 ( .A0(n22767), .A1(n22754), .B0(n22753), .Y(n22757) );
  MXI2X1 U29597 ( .A(U0_pipe10[23]), .B(n22758), .S0(n5812), .Y(n4554) );
  OAI21XL U29598 ( .A0(n22767), .A1(n22760), .B0(n22759), .Y(n22763) );
  MXI2X1 U29599 ( .A(U0_pipe10[22]), .B(n22764), .S0(n5812), .Y(n4555) );
  XOR2X1 U29600 ( .A(n22767), .B(n22766), .Y(n22768) );
  AOI21XL U29601 ( .A0(n22781), .A1(n14098), .B0(n22774), .Y(n22777) );
  INVXL U29602 ( .A(n22784), .Y(n22785) );
  AOI21XL U29603 ( .A0(n22805), .A1(n22786), .B0(n22785), .Y(n22795) );
  OAI21XL U29604 ( .A0(n22795), .A1(n22788), .B0(n22787), .Y(n22791) );
  AOI21XL U29605 ( .A0(n22805), .A1(n22798), .B0(n22797), .Y(n22801) );
  AOI21XL U29606 ( .A0(n22818), .A1(n22811), .B0(n22810), .Y(n22814) );
  OAI21XL U29607 ( .A0(n22836), .A1(n22821), .B0(n22820), .Y(n22832) );
  INVXL U29608 ( .A(n22822), .Y(n22825) );
  INVXL U29609 ( .A(n22823), .Y(n22824) );
  AOI21XL U29610 ( .A0(n22858), .A1(n22840), .B0(n22839), .Y(n22844) );
  INVXL U29611 ( .A(n22848), .Y(n22850) );
  OAI21XL U29612 ( .A0(n22871), .A1(n22867), .B0(n22868), .Y(n22865) );
  XOR2XL U29613 ( .A(n22877), .B(n22876), .Y(n22878) );
  XOR2XL U29614 ( .A(n22881), .B(n22880), .Y(n22882) );
  INVXL U29615 ( .A(n22885), .Y(n22908) );
  INVXL U29616 ( .A(n22886), .Y(n22907) );
  NOR2XL U29617 ( .A(n22907), .B(n24606), .Y(n23091) );
  NOR2XL U29618 ( .A(n23093), .B(n23091), .Y(n23085) );
  INVXL U29619 ( .A(n22887), .Y(n22909) );
  NOR2XL U29620 ( .A(n22909), .B(n24610), .Y(n22888) );
  NAND2XL U29621 ( .A(n23085), .B(n23087), .Y(n22912) );
  INVXL U29622 ( .A(n22889), .Y(n22902) );
  NOR2XL U29623 ( .A(n22902), .B(n24602), .Y(n22904) );
  INVXL U29624 ( .A(n22890), .Y(n22901) );
  NOR2XL U29625 ( .A(n22901), .B(n24600), .Y(n23106) );
  NOR2XL U29626 ( .A(n22904), .B(n23106), .Y(n22906) );
  NOR2XL U29627 ( .A(n22891), .B(n24851), .Y(n23120) );
  INVXL U29628 ( .A(n23120), .Y(n22896) );
  INVXL U29629 ( .A(n22892), .Y(n22894) );
  NOR2XL U29630 ( .A(n22894), .B(n24590), .Y(n22893) );
  INVXL U29631 ( .A(n22893), .Y(n22895) );
  AOI21XL U29632 ( .A0(n22896), .A1(n22895), .B0(n8002), .Y(n23116) );
  INVXL U29633 ( .A(n22897), .Y(n22898) );
  NOR2XL U29634 ( .A(n22898), .B(n24596), .Y(n22900) );
  NAND2XL U29635 ( .A(n22898), .B(n24596), .Y(n22899) );
  OAI21XL U29636 ( .A0(n23116), .A1(n22900), .B0(n22899), .Y(n23104) );
  NAND2XL U29637 ( .A(n22901), .B(n24600), .Y(n23105) );
  NAND2XL U29638 ( .A(n22902), .B(n24602), .Y(n22903) );
  OAI21XL U29639 ( .A0(n22904), .A1(n23105), .B0(n22903), .Y(n22905) );
  AOI21XL U29640 ( .A0(n22906), .A1(n23104), .B0(n22905), .Y(n23083) );
  NAND2XL U29641 ( .A(n22907), .B(n24606), .Y(n23099) );
  NAND2XL U29642 ( .A(n22908), .B(n24608), .Y(n23094) );
  OAI21XL U29643 ( .A0(n23093), .A1(n23099), .B0(n23094), .Y(n23084) );
  NAND2XL U29644 ( .A(n22909), .B(n24610), .Y(n23086) );
  INVXL U29645 ( .A(n23086), .Y(n22910) );
  INVXL U29646 ( .A(n22914), .Y(n22921) );
  NOR2XL U29647 ( .A(n22921), .B(n24623), .Y(n23066) );
  INVXL U29648 ( .A(n22915), .Y(n22920) );
  INVXL U29649 ( .A(n23065), .Y(n22916) );
  NAND2X1 U29650 ( .A(n23056), .B(n22919), .Y(n22929) );
  NAND2XL U29651 ( .A(n22920), .B(n24621), .Y(n23064) );
  INVXL U29652 ( .A(n23064), .Y(n22924) );
  NAND2XL U29653 ( .A(n22921), .B(n24623), .Y(n23074) );
  NAND2XL U29654 ( .A(n22925), .B(n24631), .Y(n23060) );
  INVXL U29655 ( .A(n23060), .Y(n23054) );
  NAND2XL U29656 ( .A(n22926), .B(n24633), .Y(n23055) );
  INVXL U29657 ( .A(n23055), .Y(n22927) );
  INVX1 U29658 ( .A(n22933), .Y(n22947) );
  OR2X2 U29659 ( .A(n24661), .B(n22947), .Y(n23022) );
  OR2X2 U29660 ( .A(n22942), .B(n24654), .Y(n23032) );
  INVXL U29661 ( .A(n22934), .Y(n22941) );
  NOR2XL U29662 ( .A(n22941), .B(n24652), .Y(n23030) );
  INVXL U29663 ( .A(n23030), .Y(n23037) );
  INVXL U29664 ( .A(n22936), .Y(n22938) );
  NOR2X1 U29665 ( .A(n22946), .B(n23026), .Y(n23001) );
  NAND2X1 U29666 ( .A(n22954), .B(n23001), .Y(n22956) );
  NAND2XL U29667 ( .A(n22938), .B(n24649), .Y(n23047) );
  INVXL U29668 ( .A(n23047), .Y(n23041) );
  INVXL U29669 ( .A(n23042), .Y(n22940) );
  NAND2XL U29670 ( .A(n22941), .B(n24652), .Y(n23036) );
  INVXL U29671 ( .A(n23036), .Y(n22944) );
  NAND2XL U29672 ( .A(n22942), .B(n24654), .Y(n23031) );
  INVXL U29673 ( .A(n23031), .Y(n22943) );
  NAND2X1 U29674 ( .A(n24661), .B(n22947), .Y(n23021) );
  INVXL U29675 ( .A(n23021), .Y(n23015) );
  INVXL U29676 ( .A(n23016), .Y(n22948) );
  NAND2XL U29677 ( .A(n24666), .B(n22949), .Y(n23005) );
  INVXL U29678 ( .A(n23005), .Y(n22950) );
  INVXL U29679 ( .A(n22957), .Y(n22961) );
  NOR2XL U29680 ( .A(n24679), .B(n22961), .Y(n22990) );
  INVXL U29681 ( .A(n22958), .Y(n22962) );
  NAND2XL U29682 ( .A(n24679), .B(n22961), .Y(n22989) );
  NAND2XL U29683 ( .A(n22962), .B(n24680), .Y(n22963) );
  INVXL U29684 ( .A(n22985), .Y(n22964) );
  AOI21X2 U29685 ( .A0(n22984), .A1(n22986), .B0(n22964), .Y(n22977) );
  NAND2XL U29686 ( .A(n22965), .B(n24687), .Y(n22966) );
  MXI2X1 U29687 ( .A(U0_pipe11[26]), .B(n22973), .S0(n24784), .Y(n4523) );
  XOR2X1 U29688 ( .A(n22975), .B(n22974), .Y(n22976) );
  MXI2X1 U29689 ( .A(U0_pipe11[25]), .B(n22976), .S0(n6888), .Y(n4524) );
  OAI21XL U29690 ( .A0(n22997), .A1(n22978), .B0(n22977), .Y(n22981) );
  XNOR2X1 U29691 ( .A(n22981), .B(n22980), .Y(n22982) );
  MXI2X1 U29692 ( .A(U0_pipe11[24]), .B(n22982), .S0(n6888), .Y(n4525) );
  OAI21XL U29693 ( .A0(n22997), .A1(n22990), .B0(n22989), .Y(n22993) );
  XNOR2X1 U29694 ( .A(n22993), .B(n22992), .Y(n22994) );
  MXI2X1 U29695 ( .A(U0_pipe11[20]), .B(n23008), .S0(n22620), .Y(n4529) );
  INVXL U29696 ( .A(n23014), .Y(n23024) );
  AOI21XL U29697 ( .A0(n23024), .A1(n23022), .B0(n23015), .Y(n23019) );
  XOR2X1 U29698 ( .A(n23019), .B(n23018), .Y(n23020) );
  MXI2X1 U29699 ( .A(U0_pipe11[18]), .B(n23020), .S0(n22620), .Y(n4531) );
  INVXL U29700 ( .A(n23027), .Y(n23028) );
  OAI21XL U29701 ( .A0(n23039), .A1(n23030), .B0(n23036), .Y(n23034) );
  NAND2XL U29702 ( .A(n23037), .B(n23036), .Y(n23038) );
  AOI21XL U29703 ( .A0(n23049), .A1(n22937), .B0(n23041), .Y(n23045) );
  NAND2XL U29704 ( .A(n23043), .B(n23042), .Y(n23044) );
  NAND2XL U29705 ( .A(n22937), .B(n23047), .Y(n23048) );
  OAI21XL U29706 ( .A0(n23081), .A1(n23053), .B0(n23052), .Y(n23062) );
  AOI21XL U29707 ( .A0(n23062), .A1(n22919), .B0(n23054), .Y(n23058) );
  INVXL U29708 ( .A(n23066), .Y(n23075) );
  INVXL U29709 ( .A(n23068), .Y(n23070) );
  NAND2XL U29710 ( .A(n23075), .B(n23074), .Y(n23076) );
  INVXL U29711 ( .A(n23083), .Y(n23102) );
  AOI21XL U29712 ( .A0(n23102), .A1(n23085), .B0(n23084), .Y(n23089) );
  INVXL U29713 ( .A(n23093), .Y(n23095) );
  OAI21XL U29714 ( .A0(n23113), .A1(n23106), .B0(n23105), .Y(n23109) );
  XOR2XL U29715 ( .A(n23117), .B(n23116), .Y(n23118) );
  XOR2XL U29716 ( .A(n23121), .B(n23120), .Y(n23122) );
  NAND2XL U29717 ( .A(U0_pipe11[0]), .B(U0_pipe10[0]), .Y(n23125) );
  OAI21XL U29718 ( .A0(n23126), .A1(n23125), .B0(n23124), .Y(n23188) );
  OAI21XL U29719 ( .A0(n23174), .A1(n23131), .B0(n23167), .Y(n23135) );
  OR2X2 U29720 ( .A(n23133), .B(U2_A_i_d[1]), .Y(n23171) );
  NAND2XL U29721 ( .A(n23133), .B(U2_A_i_d[1]), .Y(n23168) );
  OAI21XL U29722 ( .A0(n23137), .A1(n23183), .B0(n23185), .Y(n23142) );
  CMPR22X1 U29723 ( .A(U0_pipe11[2]), .B(U0_pipe10[2]), .CO(n23139), .S(n23127) );
  OAI21XL U29724 ( .A0(n23144), .A1(n23194), .B0(n23196), .Y(n23149) );
  CMPR22X1 U29725 ( .A(U0_pipe5[2]), .B(U0_pipe4[2]), .CO(n23146), .S(n22428)
         );
  OAI21XL U29726 ( .A0(n23153), .A1(n23152), .B0(n23151), .Y(n23254) );
  CMPR22X1 U29727 ( .A(U0_pipe14[2]), .B(n28728), .CO(n23155), .S(n22728) );
  OAI21XL U29728 ( .A0(n23159), .A1(n23212), .B0(n23214), .Y(n23164) );
  CMPR22X1 U29729 ( .A(U0_pipe7[2]), .B(U0_pipe6[2]), .CO(n23161), .S(n22104)
         );
  NAND2XL U29730 ( .A(n23171), .B(n23166), .Y(n23173) );
  INVXL U29731 ( .A(n23168), .Y(n23169) );
  AOI21XL U29732 ( .A0(n23171), .A1(n23170), .B0(n23169), .Y(n23172) );
  OAI21XL U29733 ( .A0(n23174), .A1(n23173), .B0(n23172), .Y(n23274) );
  INVXL U29734 ( .A(n23274), .Y(n23223) );
  CMPR32X1 U29735 ( .A(n23177), .B(n23176), .C(n23175), .CO(n23178), .S(n23133) );
  OAI21XL U29736 ( .A0(n23186), .A1(n23185), .B0(n23184), .Y(n23187) );
  CMPR22X1 U29737 ( .A(U0_pipe11[3]), .B(U0_pipe10[3]), .CO(n23191), .S(n23138) );
  OAI21XL U29738 ( .A0(n23197), .A1(n23196), .B0(n23195), .Y(n23198) );
  CMPR22X1 U29739 ( .A(U0_pipe5[3]), .B(U0_pipe4[3]), .CO(n23202), .S(n23145)
         );
  OAI21XL U29740 ( .A0(n23205), .A1(n23249), .B0(n23251), .Y(n23210) );
  CMPR22X1 U29741 ( .A(U0_pipe14[3]), .B(n28727), .CO(n23207), .S(n23154) );
  OAI21XL U29742 ( .A0(n23215), .A1(n23214), .B0(n23213), .Y(n23216) );
  CMPR22X1 U29743 ( .A(U0_pipe7[3]), .B(U0_pipe6[3]), .CO(n23220), .S(n23160)
         );
  OAI21XL U29744 ( .A0(n23223), .A1(n23268), .B0(n23270), .Y(n23230) );
  CMPR32X1 U29745 ( .A(n23225), .B(n23224), .C(U2_A_i_d[2]), .CO(n23226), .S(
        n23179) );
  NAND2XL U29746 ( .A(n23227), .B(n23226), .Y(n23269) );
  CMPR22X1 U29747 ( .A(U0_pipe11[4]), .B(U0_pipe10[4]), .CO(n23235), .S(n23190) );
  CMPR22X1 U29748 ( .A(U0_pipe5[4]), .B(U0_pipe4[4]), .CO(n23244), .S(n23201)
         );
  NAND2XL U29749 ( .A(n23245), .B(n23292), .Y(n23246) );
  OAI21XL U29750 ( .A0(n23252), .A1(n23251), .B0(n23250), .Y(n23253) );
  CMPR22X1 U29751 ( .A(U0_pipe14[4]), .B(n28823), .CO(n23257), .S(n23206) );
  CMPR22X1 U29752 ( .A(U0_pipe7[4]), .B(U0_pipe6[4]), .CO(n23263), .S(n23219)
         );
  NAND2XL U29753 ( .A(n23264), .B(n23282), .Y(n23265) );
  NOR2XL U29754 ( .A(n23268), .B(n23271), .Y(n23273) );
  OAI21XL U29755 ( .A0(n23271), .A1(n23270), .B0(n23269), .Y(n23272) );
  CMPR32X1 U29756 ( .A(n23276), .B(n23275), .C(U2_A_i_d[3]), .CO(n23277), .S(
        n23227) );
  NOR2XL U29757 ( .A(n23278), .B(n23277), .Y(n23360) );
  NAND2XL U29758 ( .A(n23278), .B(n23277), .Y(n23362) );
  OAI21XL U29759 ( .A0(n23284), .A1(n23283), .B0(n23282), .Y(n23378) );
  CMPR22X1 U29760 ( .A(U0_pipe7[5]), .B(U0_pipe6[5]), .CO(n23287), .S(n23262)
         );
  OAI21XL U29761 ( .A0(n23294), .A1(n23293), .B0(n23292), .Y(n23394) );
  CMPR22X1 U29762 ( .A(U0_pipe5[5]), .B(U0_pipe4[5]), .CO(n23297), .S(n23243)
         );
  CMPR22X1 U29763 ( .A(U0_pipe14[5]), .B(n28822), .CO(n23304), .S(n23256) );
  OAI21XL U29764 ( .A0(n23312), .A1(n23311), .B0(n23310), .Y(n23417) );
  CMPR22X1 U29765 ( .A(U0_pipe11[5]), .B(U0_pipe10[5]), .CO(n23315), .S(n23234) );
  CMPR32X1 U29766 ( .A(n23322), .B(n23321), .C(U2_A_i_d[4]), .CO(n23323), .S(
        n23278) );
  INVXL U29767 ( .A(n23363), .Y(n23325) );
  NAND2XL U29768 ( .A(n23324), .B(n23323), .Y(n23361) );
  OAI21XL U29769 ( .A0(n23329), .A1(n23372), .B0(n23375), .Y(n23334) );
  CMPR22X1 U29770 ( .A(U0_pipe7[6]), .B(U0_pipe6[6]), .CO(n23331), .S(n23286)
         );
  OAI21XL U29771 ( .A0(n23336), .A1(n23388), .B0(n23391), .Y(n23341) );
  CMPR22X1 U29772 ( .A(U0_pipe5[6]), .B(U0_pipe4[6]), .CO(n23338), .S(n23296)
         );
  OAI21XL U29773 ( .A0(n23346), .A1(n23345), .B0(n23344), .Y(n23454) );
  CMPR22X1 U29774 ( .A(U0_pipe14[6]), .B(n28726), .CO(n23349), .S(n23303) );
  OAI21XL U29775 ( .A0(n23353), .A1(n23411), .B0(n23414), .Y(n23358) );
  CMPR22X1 U29776 ( .A(U0_pipe11[6]), .B(U0_pipe10[6]), .CO(n23355), .S(n23314) );
  NOR2XL U29777 ( .A(n23360), .B(n23363), .Y(n23471) );
  OAI21XL U29778 ( .A0(n23363), .A1(n23362), .B0(n23361), .Y(n23476) );
  AOI21XL U29779 ( .A0(n23364), .A1(n23471), .B0(n23476), .Y(n23427) );
  CMPR32X1 U29780 ( .A(n23366), .B(n23365), .C(U2_A_i_d[5]), .CO(n23367), .S(
        n23324) );
  OAI21XL U29781 ( .A0(n23376), .A1(n23375), .B0(n23374), .Y(n23377) );
  OAI21XL U29782 ( .A0(n23382), .A1(n23381), .B0(n23380), .Y(n23862) );
  CMPR22X1 U29783 ( .A(U0_pipe7[7]), .B(U0_pipe6[7]), .CO(n23384), .S(n23330)
         );
  OAI21XL U29784 ( .A0(n23392), .A1(n23391), .B0(n23390), .Y(n23393) );
  OAI21XL U29785 ( .A0(n23398), .A1(n23397), .B0(n23396), .Y(n23843) );
  CMPR22X1 U29786 ( .A(U0_pipe5[7]), .B(U0_pipe4[7]), .CO(n23400), .S(n23337)
         );
  OAI21XL U29787 ( .A0(n23404), .A1(n23448), .B0(n23451), .Y(n23409) );
  CMPR22X1 U29788 ( .A(U0_pipe14[7]), .B(n28821), .CO(n23406), .S(n23348) );
  CLKINVX3 U29789 ( .A(n28997), .Y(n23559) );
  OAI21XL U29790 ( .A0(n23415), .A1(n23414), .B0(n23413), .Y(n23416) );
  OAI21XL U29791 ( .A0(n23421), .A1(n23420), .B0(n23419), .Y(n23824) );
  CMPR22X1 U29792 ( .A(U0_pipe11[7]), .B(U0_pipe10[7]), .CO(n23423), .S(n23354) );
  OAI21XL U29793 ( .A0(n23427), .A1(n23470), .B0(n23473), .Y(n23434) );
  CMPR32X1 U29794 ( .A(n23429), .B(n23428), .C(U2_A_i_d[6]), .CO(n23430), .S(
        n23368) );
  INVXL U29795 ( .A(n23474), .Y(n23432) );
  NAND2XL U29796 ( .A(n23431), .B(n23430), .Y(n23472) );
  OAI21XL U29797 ( .A0(n23590), .A1(n23514), .B0(n23516), .Y(n23440) );
  CMPR22X1 U29798 ( .A(U0_pipe11[8]), .B(U0_pipe10[8]), .CO(n23437), .S(n23422) );
  OAI21XL U29799 ( .A0(n23603), .A1(n23498), .B0(n23500), .Y(n23446) );
  CMPR22X1 U29800 ( .A(U0_pipe5[8]), .B(U0_pipe4[8]), .CO(n23443), .S(n23399)
         );
  OAI21XL U29801 ( .A0(n23452), .A1(n23451), .B0(n23450), .Y(n23453) );
  OAI21XL U29802 ( .A0(n23458), .A1(n23457), .B0(n23456), .Y(n23892) );
  CMPR22X1 U29803 ( .A(U0_pipe14[8]), .B(n28820), .CO(n23460), .S(n23405) );
  OAI21XL U29804 ( .A0(n23625), .A1(n23488), .B0(n23490), .Y(n23468) );
  CMPR22X1 U29805 ( .A(U0_pipe7[8]), .B(U0_pipe6[8]), .CO(n23465), .S(n23383)
         );
  NOR2XL U29806 ( .A(n23470), .B(n23474), .Y(n23477) );
  NAND2XL U29807 ( .A(n23471), .B(n23477), .Y(n23479) );
  OAI21XL U29808 ( .A0(n23474), .A1(n23473), .B0(n23472), .Y(n23475) );
  AOI21XL U29809 ( .A0(n23477), .A1(n23476), .B0(n23475), .Y(n23478) );
  CMPR32X1 U29810 ( .A(n23482), .B(n23481), .C(U2_A_i_d[7]), .CO(n23483), .S(
        n23431) );
  NOR2XL U29811 ( .A(n23484), .B(n23483), .Y(n23570) );
  NAND2XL U29812 ( .A(n23485), .B(n23572), .Y(n23486) );
  OAI21XL U29813 ( .A0(n23491), .A1(n23490), .B0(n23489), .Y(n23623) );
  OAI21XL U29814 ( .A0(n23625), .A1(n23493), .B0(n23492), .Y(n23534) );
  CMPR22X1 U29815 ( .A(U0_pipe7[9]), .B(U0_pipe6[9]), .CO(n23495), .S(n23464)
         );
  OAI21XL U29816 ( .A0(n23501), .A1(n23500), .B0(n23499), .Y(n23601) );
  OAI21XL U29817 ( .A0(n23603), .A1(n23503), .B0(n23502), .Y(n23543) );
  CMPR22X1 U29818 ( .A(U0_pipe5[9]), .B(U0_pipe4[9]), .CO(n23505), .S(n23442)
         );
  OAI21XL U29819 ( .A0(n23649), .A1(n23550), .B0(n23552), .Y(n23512) );
  CMPR22X1 U29820 ( .A(U0_pipe14[9]), .B(n28725), .CO(n23509), .S(n23459) );
  OAI21XL U29821 ( .A0(n23517), .A1(n23516), .B0(n23515), .Y(n23588) );
  OAI21XL U29822 ( .A0(n23590), .A1(n23519), .B0(n23518), .Y(n23563) );
  CMPR22X1 U29823 ( .A(U0_pipe11[9]), .B(U0_pipe10[9]), .CO(n23521), .S(n23436) );
  OAI21XL U29824 ( .A0(n23689), .A1(n23570), .B0(n23572), .Y(n23530) );
  CMPR32X1 U29825 ( .A(n23525), .B(n23524), .C(U2_A_i_d[8]), .CO(n23526), .S(
        n23484) );
  NAND2XL U29826 ( .A(n23527), .B(n23526), .Y(n23571) );
  CMPR22X1 U29827 ( .A(U0_pipe7[10]), .B(U0_pipe6[10]), .CO(n23536), .S(n23494) );
  CMPR22X1 U29828 ( .A(U0_pipe5[10]), .B(U0_pipe4[10]), .CO(n23545), .S(n23504) );
  OAI21XL U29829 ( .A0(n23553), .A1(n23552), .B0(n23551), .Y(n23647) );
  OAI21XL U29830 ( .A0(n23649), .A1(n23555), .B0(n23554), .Y(n23610) );
  CMPR22X1 U29831 ( .A(U0_pipe14[10]), .B(n28819), .CO(n23557), .S(n23508) );
  CMPR22X1 U29832 ( .A(U0_pipe11[10]), .B(U0_pipe10[10]), .CO(n23565), .S(
        n23520) );
  NOR2XL U29833 ( .A(n23570), .B(n23573), .Y(n23682) );
  OAI21XL U29834 ( .A0(n23573), .A1(n23572), .B0(n23571), .Y(n23687) );
  INVXL U29835 ( .A(n23687), .Y(n23574) );
  OAI21XL U29836 ( .A0(n23689), .A1(n23575), .B0(n23574), .Y(n23632) );
  NOR2XL U29837 ( .A(n23579), .B(n23578), .Y(n23681) );
  INVXL U29838 ( .A(n23681), .Y(n23631) );
  NAND2XL U29839 ( .A(n23579), .B(n23578), .Y(n23684) );
  NAND2XL U29840 ( .A(n23631), .B(n23684), .Y(n23580) );
  OAI21XL U29841 ( .A0(n23586), .A1(n23585), .B0(n23584), .Y(n23587) );
  OAI21XL U29842 ( .A0(n23590), .A1(n23812), .B0(n23821), .Y(n23656) );
  CMPR22X1 U29843 ( .A(U0_pipe11[11]), .B(U0_pipe10[11]), .CO(n23592), .S(
        n23564) );
  OAI21XL U29844 ( .A0(n23599), .A1(n23598), .B0(n23597), .Y(n23600) );
  OAI21XL U29845 ( .A0(n23603), .A1(n23831), .B0(n23840), .Y(n23665) );
  CMPR22X1 U29846 ( .A(U0_pipe5[11]), .B(U0_pipe4[11]), .CO(n23605), .S(n23544) );
  CMPR22X1 U29847 ( .A(U0_pipe14[11]), .B(n28818), .CO(n23612), .S(n23556) );
  OAI21XL U29848 ( .A0(n23621), .A1(n23620), .B0(n23619), .Y(n23622) );
  OAI21XL U29849 ( .A0(n23625), .A1(n23850), .B0(n23859), .Y(n23674) );
  CMPR22X1 U29850 ( .A(U0_pipe7[11]), .B(U0_pipe6[11]), .CO(n23627), .S(n23535) );
  INVXL U29851 ( .A(n23684), .Y(n23630) );
  AOI21XL U29852 ( .A0(n23632), .A1(n23631), .B0(n23630), .Y(n23639) );
  CMPR32X1 U29853 ( .A(n23634), .B(n23633), .C(U2_A_i_d[10]), .CO(n23635), .S(
        n23579) );
  NAND2XL U29854 ( .A(n23636), .B(n23635), .Y(n23683) );
  OAI21XL U29855 ( .A0(n23645), .A1(n23644), .B0(n23643), .Y(n23646) );
  OAI21XL U29856 ( .A0(n23649), .A1(n23880), .B0(n23889), .Y(n23699) );
  CMPR22X1 U29857 ( .A(U0_pipe14[12]), .B(n28817), .CO(n23651), .S(n23611) );
  CMPR22X1 U29858 ( .A(U0_pipe11[12]), .B(U0_pipe10[12]), .CO(n23658), .S(
        n23591) );
  NAND2XL U29859 ( .A(n23659), .B(n23729), .Y(n23660) );
  CMPR22X1 U29860 ( .A(U0_pipe5[12]), .B(U0_pipe4[12]), .CO(n23667), .S(n23604) );
  CMPR22X1 U29861 ( .A(U0_pipe7[12]), .B(U0_pipe6[12]), .CO(n23676), .S(n23626) );
  NOR2XL U29862 ( .A(n23681), .B(n23685), .Y(n23688) );
  NAND2XL U29863 ( .A(n23682), .B(n23688), .Y(n23924) );
  OAI21XL U29864 ( .A0(n23685), .A1(n23684), .B0(n23683), .Y(n23686) );
  AOI21XL U29865 ( .A0(n23688), .A1(n23687), .B0(n23686), .Y(n23932) );
  CMPR32X1 U29866 ( .A(n23691), .B(n23690), .C(U2_A_i_d[11]), .CO(n23692), .S(
        n23636) );
  NOR2XL U29867 ( .A(n23693), .B(n23692), .Y(n23788) );
  INVXL U29868 ( .A(n23788), .Y(n23740) );
  NAND2XL U29869 ( .A(n23693), .B(n23692), .Y(n23790) );
  NAND2XL U29870 ( .A(n23740), .B(n23790), .Y(n23694) );
  CMPR22X1 U29871 ( .A(U0_pipe14[13]), .B(n28816), .CO(n23701), .S(n23650) );
  OAI21XL U29872 ( .A0(n23709), .A1(n23708), .B0(n23707), .Y(n23855) );
  OAI21XL U29873 ( .A0(n23712), .A1(n23711), .B0(n23710), .Y(n23781) );
  CMPR22X1 U29874 ( .A(U0_pipe7[13]), .B(U0_pipe6[13]), .CO(n23714), .S(n23675) );
  OAI21XL U29875 ( .A0(n23720), .A1(n23719), .B0(n23718), .Y(n23836) );
  OAI21XL U29876 ( .A0(n23723), .A1(n23722), .B0(n23721), .Y(n23772) );
  CMPR22X1 U29877 ( .A(U0_pipe5[13]), .B(U0_pipe4[13]), .CO(n23725), .S(n23666) );
  OAI21XL U29878 ( .A0(n23731), .A1(n23730), .B0(n23729), .Y(n23817) );
  OAI21XL U29879 ( .A0(n23734), .A1(n23733), .B0(n23732), .Y(n23763) );
  CMPR22X1 U29880 ( .A(U0_pipe11[13]), .B(U0_pipe10[13]), .CO(n23736), .S(
        n23657) );
  INVXL U29881 ( .A(n23790), .Y(n23739) );
  AOI21XL U29882 ( .A0(n23741), .A1(n23740), .B0(n23739), .Y(n23748) );
  CMPR32X1 U29883 ( .A(n23743), .B(n23742), .C(U2_A_i_d[12]), .CO(n23744), .S(
        n23693) );
  INVXL U29884 ( .A(n23791), .Y(n23746) );
  NAND2XL U29885 ( .A(n23746), .B(n23789), .Y(n23747) );
  OAI21XL U29886 ( .A0(n23753), .A1(n23752), .B0(n23751), .Y(n23885) );
  OAI21XL U29887 ( .A0(n23756), .A1(n23755), .B0(n23754), .Y(n23803) );
  CMPR22X1 U29888 ( .A(U0_pipe14[14]), .B(n28815), .CO(n23758), .S(n23700) );
  CMPR22X1 U29889 ( .A(U0_pipe11[14]), .B(U0_pipe10[14]), .CO(n23765), .S(
        n23735) );
  CMPR22X1 U29890 ( .A(U0_pipe5[14]), .B(U0_pipe4[14]), .CO(n23774), .S(n23724) );
  CMPR22X1 U29891 ( .A(U0_pipe7[14]), .B(U0_pipe6[14]), .CO(n23783), .S(n23713) );
  NOR2XL U29892 ( .A(n23788), .B(n23791), .Y(n23923) );
  INVXL U29893 ( .A(n23923), .Y(n23793) );
  INVXL U29894 ( .A(n23929), .Y(n23792) );
  CMPR32X1 U29895 ( .A(n23796), .B(n23795), .C(U2_A_i_d[13]), .CO(n23797), .S(
        n23745) );
  INVXL U29896 ( .A(n23922), .Y(n23868) );
  NAND2XL U29897 ( .A(n23868), .B(n23926), .Y(n23799) );
  CMPR22X1 U29898 ( .A(U0_pipe14[15]), .B(n28814), .CO(n23805), .S(n23757) );
  OAI21XL U29899 ( .A0(n23815), .A1(n23814), .B0(n23813), .Y(n23816) );
  OAI21XL U29900 ( .A0(n23821), .A1(n23820), .B0(n23819), .Y(n23822) );
  CMPR22X1 U29901 ( .A(U0_pipe11[15]), .B(U0_pipe10[15]), .CO(n23826), .S(
        n23764) );
  OAI21XL U29902 ( .A0(n23834), .A1(n23833), .B0(n23832), .Y(n23835) );
  OAI21XL U29903 ( .A0(n23840), .A1(n23839), .B0(n23838), .Y(n23841) );
  CMPR22X1 U29904 ( .A(U0_pipe5[15]), .B(U0_pipe4[15]), .CO(n23845), .S(n23773) );
  OAI21XL U29905 ( .A0(n23853), .A1(n23852), .B0(n23851), .Y(n23854) );
  OAI21XL U29906 ( .A0(n23859), .A1(n23858), .B0(n23857), .Y(n23860) );
  CMPR22X1 U29907 ( .A(U0_pipe7[15]), .B(U0_pipe6[15]), .CO(n23864), .S(n23782) );
  NAND2XL U29908 ( .A(n23899), .B(n23951), .Y(n23865) );
  INVXL U29909 ( .A(n23926), .Y(n23867) );
  AOI21XL U29910 ( .A0(n23869), .A1(n23868), .B0(n23867), .Y(n23876) );
  NAND2XL U29911 ( .A(n23873), .B(n23872), .Y(n23925) );
  XOR2X1 U29912 ( .A(n23876), .B(n23875), .Y(n23877) );
  OAI21XL U29913 ( .A0(n23883), .A1(n23882), .B0(n23881), .Y(n23884) );
  OAI21XL U29914 ( .A0(n23889), .A1(n23888), .B0(n23887), .Y(n23890) );
  NAND2XL U29915 ( .A(n23893), .B(n23942), .Y(n23896) );
  CMPR22X1 U29916 ( .A(U0_pipe7[16]), .B(U0_pipe6[16]), .CO(n23901), .S(n23863) );
  CMPR22X1 U29917 ( .A(U0_pipe5[16]), .B(U0_pipe4[16]), .CO(n23909), .S(n23844) );
  CMPR22X1 U29918 ( .A(U0_pipe11[16]), .B(U0_pipe10[16]), .CO(n23917), .S(
        n23825) );
  NOR2XL U29919 ( .A(n23924), .B(n23931), .Y(n23934) );
  OAI21XL U29920 ( .A0(n23927), .A1(n23926), .B0(n23925), .Y(n23928) );
  AOI21X2 U29921 ( .A0(n23935), .A1(n23934), .B0(n23933), .Y(n24205) );
  CMPR32X1 U29922 ( .A(n23937), .B(n23936), .C(U2_A_i_d[15]), .CO(n23938), .S(
        n23873) );
  NOR2XL U29923 ( .A(n23939), .B(n23938), .Y(n24036) );
  NAND2XL U29924 ( .A(n23980), .B(n24038), .Y(n23940) );
  OAI21XL U29925 ( .A0(n23952), .A1(n23951), .B0(n23950), .Y(n24027) );
  OAI21XL U29926 ( .A0(n23962), .A1(n23961), .B0(n23960), .Y(n24015) );
  OAI21XL U29927 ( .A0(n23972), .A1(n23971), .B0(n23970), .Y(n24003) );
  INVXL U29928 ( .A(n24038), .Y(n23979) );
  AOI21XL U29929 ( .A0(n24158), .A1(n23980), .B0(n23979), .Y(n23987) );
  NOR2X2 U29930 ( .A(n23984), .B(n23983), .Y(n24039) );
  NAND2X1 U29931 ( .A(n23984), .B(n23983), .Y(n24037) );
  NAND2XL U29932 ( .A(n23985), .B(n24037), .Y(n23986) );
  CMPR22X1 U29933 ( .A(U0_pipe14[18]), .B(n28811), .CO(n23995), .S(n23944) );
  CMPR22X1 U29934 ( .A(U0_pipe11[18]), .B(U0_pipe10[18]), .CO(n24007), .S(
        n23974) );
  CMPR22X1 U29935 ( .A(U0_pipe5[18]), .B(U0_pipe4[18]), .CO(n24019), .S(n23964) );
  CMPR22X1 U29936 ( .A(U0_pipe7[18]), .B(U0_pipe6[18]), .CO(n24031), .S(n23954) );
  AOI21XL U29937 ( .A0(n24158), .A1(n24091), .B0(n24094), .Y(n24045) );
  NAND2XL U29938 ( .A(n24043), .B(n24042), .Y(n24092) );
  OAI21XL U29939 ( .A0(n24050), .A1(n24049), .B0(n24048), .Y(n24108) );
  OAI21XL U29940 ( .A0(n24061), .A1(n24060), .B0(n24059), .Y(n24145) );
  OAI21XL U29941 ( .A0(n24072), .A1(n24071), .B0(n24070), .Y(n24133) );
  NAND2XL U29942 ( .A(n24074), .B(n24131), .Y(n24077) );
  OAI21XL U29943 ( .A0(n24083), .A1(n24082), .B0(n24081), .Y(n24120) );
  AOI21XL U29944 ( .A0(n24084), .A1(n24117), .B0(n24120), .Y(n24089) );
  NAND2X1 U29945 ( .A(n24091), .B(n6986), .Y(n24154) );
  INVXL U29946 ( .A(n24154), .Y(n24096) );
  INVXL U29947 ( .A(n24092), .Y(n24093) );
  AOI21XL U29948 ( .A0(n24158), .A1(n24096), .B0(n24095), .Y(n24103) );
  INVXL U29949 ( .A(n24156), .Y(n24101) );
  NAND2XL U29950 ( .A(n24100), .B(n24099), .Y(n24155) );
  OAI21XL U29951 ( .A0(n24111), .A1(n24110), .B0(n24109), .Y(n24169) );
  OAI21XL U29952 ( .A0(n24123), .A1(n24122), .B0(n24121), .Y(n24193) );
  OAI21XL U29953 ( .A0(n24136), .A1(n24135), .B0(n24134), .Y(n24185) );
  OAI21XL U29954 ( .A0(n24148), .A1(n24147), .B0(n24146), .Y(n24177) );
  NOR2XL U29955 ( .A(n24154), .B(n24156), .Y(n24199) );
  OAI21X1 U29956 ( .A0(n24157), .A1(n24156), .B0(n24155), .Y(n24202) );
  AOI21XL U29957 ( .A0(n24158), .A1(n24199), .B0(n24202), .Y(n24165) );
  CMPR32X1 U29958 ( .A(n24160), .B(n24159), .C(U2_A_i_d[19]), .CO(n24162), .S(
        n24100) );
  CMPR22X1 U29959 ( .A(U0_pipe14[21]), .B(n28808), .CO(n24171), .S(n24113) );
  CMPR22X1 U29960 ( .A(U0_pipe7[21]), .B(U0_pipe6[21]), .CO(n24179), .S(n24150) );
  CMPR22X1 U29961 ( .A(U0_pipe5[21]), .B(U0_pipe4[21]), .CO(n24187), .S(n24138) );
  CMPR22X1 U29962 ( .A(U0_pipe11[21]), .B(U0_pipe10[21]), .CO(n24195), .S(
        n24125) );
  NAND2X1 U29963 ( .A(n24199), .B(n24161), .Y(n24204) );
  AOI21X1 U29964 ( .A0(n24202), .A1(n24161), .B0(n24201), .Y(n24203) );
  CMPR32X1 U29965 ( .A(n24207), .B(n24206), .C(U2_A_i_d[20]), .CO(n24208), .S(
        n24163) );
  OR2X2 U29966 ( .A(n24209), .B(n24208), .Y(n24246) );
  NAND2XL U29967 ( .A(n24209), .B(n24208), .Y(n24244) );
  OAI21XL U29968 ( .A0(n24214), .A1(n24213), .B0(n24212), .Y(n24256) );
  OAI21XL U29969 ( .A0(n24222), .A1(n24221), .B0(n24220), .Y(n24264) );
  OAI21XL U29970 ( .A0(n24230), .A1(n24229), .B0(n24228), .Y(n24272) );
  OAI21XL U29971 ( .A0(n24238), .A1(n24237), .B0(n24236), .Y(n24280) );
  INVXL U29972 ( .A(n24244), .Y(n24245) );
  CMPR32X1 U29973 ( .A(n24249), .B(n24248), .C(U2_A_i_d[21]), .CO(n24250), .S(
        n24209) );
  CMPR22X1 U29974 ( .A(U0_pipe14[23]), .B(n28937), .CO(n24258), .S(n24216) );
  CMPR22X1 U29975 ( .A(U0_pipe7[23]), .B(U0_pipe6[23]), .CO(n24266), .S(n24224) );
  CMPR22X1 U29976 ( .A(U0_pipe5[23]), .B(U0_pipe4[23]), .CO(n24274), .S(n24232) );
  CMPR22X1 U29977 ( .A(U0_pipe11[23]), .B(U0_pipe10[23]), .CO(n24282), .S(
        n24240) );
  CMPR32X1 U29978 ( .A(n24290), .B(n24289), .C(U2_A_i_d[22]), .CO(n24291), .S(
        n24251) );
  OR2X2 U29979 ( .A(n24292), .B(n24291), .Y(n24329) );
  OAI21XL U29980 ( .A0(n24297), .A1(n24296), .B0(n24295), .Y(n24340) );
  OAI21XL U29981 ( .A0(n24305), .A1(n24304), .B0(n24303), .Y(n24348) );
  OAI21XL U29982 ( .A0(n24313), .A1(n24312), .B0(n24311), .Y(n24356) );
  OAI21XL U29983 ( .A0(n24321), .A1(n24320), .B0(n24319), .Y(n24364) );
  CMPR32X1 U29984 ( .A(n24332), .B(n24331), .C(U2_A_i_d[23]), .CO(n24333), .S(
        n24292) );
  CMPR22X1 U29985 ( .A(U0_pipe14[25]), .B(n28935), .CO(n24342), .S(n24299) );
  CMPR22X1 U29986 ( .A(U0_pipe11[25]), .B(U0_pipe10[25]), .CO(n24350), .S(
        n24307) );
  CMPR22X1 U29987 ( .A(U0_pipe5[25]), .B(U0_pipe4[25]), .CO(n24358), .S(n24315) );
  CMPR22X1 U29988 ( .A(U0_pipe7[25]), .B(U0_pipe6[25]), .CO(n24366), .S(n24323) );
  CMPR32X1 U29989 ( .A(n24373), .B(n24372), .C(U2_A_i_d[24]), .CO(n24374), .S(
        n24334) );
  OR2X2 U29990 ( .A(n24375), .B(n24374), .Y(n24377) );
  MXI2X1 U29991 ( .A(U2_pipe1[25]), .B(n24379), .S0(n21700), .Y(n4145) );
  CMPR22X1 U29992 ( .A(U0_pipe14[26]), .B(n29002), .CO(n24385), .S(n24341) );
  OAI21XL U29993 ( .A0(n24383), .A1(n24382), .B0(n24381), .Y(n24384) );
  CMPR32X1 U29994 ( .A(n24386), .B(n24385), .C(n24384), .S(n24387) );
  CMPR22X1 U29995 ( .A(U0_pipe7[26]), .B(U0_pipe6[26]), .CO(n24392), .S(n24365) );
  OAI21XL U29996 ( .A0(n24390), .A1(n24389), .B0(n24388), .Y(n24391) );
  CMPR32X1 U29997 ( .A(n24393), .B(n24392), .C(n24391), .S(n24394) );
  CMPR22X1 U29998 ( .A(U0_pipe5[26]), .B(U0_pipe4[26]), .CO(n24399), .S(n24357) );
  OAI21XL U29999 ( .A0(n24397), .A1(n24396), .B0(n24395), .Y(n24398) );
  CMPR32X1 U30000 ( .A(n24400), .B(n24399), .C(n24398), .S(n24401) );
  CMPR22X1 U30001 ( .A(U0_pipe11[26]), .B(U0_pipe10[26]), .CO(n24406), .S(
        n24349) );
  OAI21XL U30002 ( .A0(n24404), .A1(n24403), .B0(n24402), .Y(n24405) );
  CMPR32X1 U30003 ( .A(n24407), .B(n24406), .C(n24405), .S(n24408) );
  CMPR32X1 U30004 ( .A(n24414), .B(n29010), .C(n24413), .CO(n24415), .S(n13499) );
  INVXL U30005 ( .A(n24416), .Y(n24418) );
  OAI21XL U30006 ( .A0(n24447), .A1(n24423), .B0(n24422), .Y(n24428) );
  MXI2X1 U30007 ( .A(U0_pipe2[24]), .B(n24429), .S0(n24784), .Y(n4379) );
  INVXL U30008 ( .A(n24431), .Y(n24432) );
  MXI2X1 U30009 ( .A(U0_pipe2[23]), .B(n24438), .S0(n6888), .Y(n4380) );
  OAI21XL U30010 ( .A0(n24447), .A1(n24440), .B0(n24439), .Y(n24443) );
  MXI2X1 U30011 ( .A(U0_pipe2[22]), .B(n24444), .S0(n5812), .Y(n4381) );
  NAND2XL U30012 ( .A(n24445), .B(n24879), .Y(n24884) );
  XOR2X1 U30013 ( .A(n24447), .B(n24446), .Y(n24448) );
  INVXL U30014 ( .A(n24465), .Y(n24475) );
  AOI21XL U30015 ( .A0(n24475), .A1(n24467), .B0(n24466), .Y(n24471) );
  INVXL U30016 ( .A(n24478), .Y(n24479) );
  OAI21XL U30017 ( .A0(n24490), .A1(n24482), .B0(n24481), .Y(n24486) );
  NAND2XL U30018 ( .A(n24488), .B(n24903), .Y(n24908) );
  AOI21XL U30019 ( .A0(n24501), .A1(n24493), .B0(n24492), .Y(n24497) );
  NAND2XL U30020 ( .A(n24912), .B(n24499), .Y(n24916) );
  AOI21XL U30021 ( .A0(n24515), .A1(n24507), .B0(n24506), .Y(n24511) );
  OAI21XL U30022 ( .A0(n24535), .A1(n24518), .B0(n24517), .Y(n24531) );
  INVXL U30023 ( .A(n24519), .Y(n24522) );
  INVXL U30024 ( .A(n24520), .Y(n24521) );
  INVXL U30025 ( .A(n24523), .Y(n24525) );
  INVXL U30026 ( .A(n24529), .Y(n24933) );
  NAND2XL U30027 ( .A(n24933), .B(n24931), .Y(n24937) );
  AOI21XL U30028 ( .A0(n24556), .A1(n24539), .B0(n24538), .Y(n24543) );
  INVXL U30029 ( .A(n24547), .Y(n24549) );
  OAI21XL U30030 ( .A0(n24569), .A1(n24565), .B0(n24566), .Y(n24563) );
  XOR2XL U30031 ( .A(n24575), .B(n24574), .Y(n24576) );
  XOR2XL U30032 ( .A(n24579), .B(n24578), .Y(n24580) );
  XNOR2XL U30033 ( .A(n24581), .B(U2_A_r_d[0]), .Y(n24986) );
  INVXL U30034 ( .A(n24582), .Y(n24609) );
  NOR2XL U30035 ( .A(n24609), .B(n24608), .Y(n24819) );
  INVXL U30036 ( .A(n24583), .Y(n24607) );
  NOR2XL U30037 ( .A(n24607), .B(n24606), .Y(n24817) );
  NOR2XL U30038 ( .A(n24819), .B(n24817), .Y(n24812) );
  INVXL U30039 ( .A(n24584), .Y(n24611) );
  NAND2XL U30040 ( .A(n24812), .B(n24585), .Y(n24614) );
  INVXL U30041 ( .A(n24586), .Y(n24603) );
  NOR2XL U30042 ( .A(n24603), .B(n24602), .Y(n24833) );
  INVXL U30043 ( .A(n24587), .Y(n24601) );
  NOR2XL U30044 ( .A(n24601), .B(n24600), .Y(n24832) );
  NOR2XL U30045 ( .A(n24833), .B(n24832), .Y(n24605) );
  INVXL U30046 ( .A(n25448), .Y(n24852) );
  NOR2XL U30047 ( .A(n24852), .B(n24851), .Y(n24848) );
  INVXL U30048 ( .A(n24848), .Y(n24594) );
  INVXL U30049 ( .A(n24588), .Y(n24591) );
  NOR2XL U30050 ( .A(n24591), .B(n24590), .Y(n24589) );
  INVXL U30051 ( .A(n24589), .Y(n24593) );
  AOI21XL U30052 ( .A0(n24594), .A1(n24593), .B0(n24592), .Y(n24844) );
  INVXL U30053 ( .A(n24595), .Y(n24597) );
  NOR2XL U30054 ( .A(n24597), .B(n24596), .Y(n24599) );
  NAND2XL U30055 ( .A(n24597), .B(n24596), .Y(n24598) );
  OAI21XL U30056 ( .A0(n24844), .A1(n24599), .B0(n24598), .Y(n24830) );
  NAND2XL U30057 ( .A(n24601), .B(n24600), .Y(n24831) );
  NAND2XL U30058 ( .A(n24603), .B(n24602), .Y(n24834) );
  OAI21XL U30059 ( .A0(n24833), .A1(n24831), .B0(n24834), .Y(n24604) );
  AOI21XL U30060 ( .A0(n24605), .A1(n24830), .B0(n24604), .Y(n24810) );
  NAND2XL U30061 ( .A(n24607), .B(n24606), .Y(n24825) );
  NAND2XL U30062 ( .A(n24609), .B(n24608), .Y(n24820) );
  OAI21XL U30063 ( .A0(n24819), .A1(n24825), .B0(n24820), .Y(n24811) );
  OAI21XL U30064 ( .A0(n24614), .A1(n24810), .B0(n24613), .Y(n24775) );
  INVXL U30065 ( .A(n24616), .Y(n24624) );
  NOR2XL U30066 ( .A(n24624), .B(n24623), .Y(n24792) );
  NOR2XL U30067 ( .A(n24627), .B(n24792), .Y(n24630) );
  INVXL U30068 ( .A(n24617), .Y(n24622) );
  NOR2XL U30069 ( .A(n24622), .B(n24621), .Y(n24791) );
  INVXL U30070 ( .A(n24791), .Y(n24618) );
  NAND2XL U30071 ( .A(n24630), .B(n24618), .Y(n24777) );
  INVXL U30072 ( .A(n24620), .Y(n24632) );
  NAND2XL U30073 ( .A(n7999), .B(n24779), .Y(n24637) );
  NOR2XL U30074 ( .A(n24777), .B(n24637), .Y(n24639) );
  NAND2XL U30075 ( .A(n24622), .B(n24621), .Y(n24790) );
  INVXL U30076 ( .A(n24790), .Y(n24629) );
  NAND2XL U30077 ( .A(n24624), .B(n24623), .Y(n24793) );
  OAI21XL U30078 ( .A0(n24627), .A1(n24793), .B0(n24626), .Y(n24628) );
  AOI21XL U30079 ( .A0(n24630), .A1(n24629), .B0(n24628), .Y(n24776) );
  OAI21X1 U30080 ( .A0(n24776), .A1(n24637), .B0(n24636), .Y(n24638) );
  OR2X2 U30081 ( .A(n24664), .B(n24663), .Y(n24739) );
  NAND2X1 U30082 ( .A(n24735), .B(n24739), .Y(n24669) );
  INVXL U30083 ( .A(n24643), .Y(n24660) );
  OR2X2 U30084 ( .A(n24655), .B(n24654), .Y(n24758) );
  INVXL U30085 ( .A(n24645), .Y(n24653) );
  NOR2XL U30086 ( .A(n24653), .B(n24652), .Y(n24756) );
  INVXL U30087 ( .A(n24756), .Y(n24762) );
  INVXL U30088 ( .A(n24647), .Y(n24650) );
  NAND2XL U30089 ( .A(n6984), .B(n24648), .Y(n24752) );
  NOR2XL U30090 ( .A(n24659), .B(n24752), .Y(n24730) );
  NAND2X1 U30091 ( .A(n24671), .B(n24730), .Y(n24673) );
  NAND2XL U30092 ( .A(n24650), .B(n24649), .Y(n24771) );
  NAND2XL U30093 ( .A(n24653), .B(n24652), .Y(n24761) );
  INVXL U30094 ( .A(n24761), .Y(n24657) );
  NAND2XL U30095 ( .A(n24655), .B(n24654), .Y(n24757) );
  INVXL U30096 ( .A(n24757), .Y(n24656) );
  INVXL U30097 ( .A(n24738), .Y(n24733) );
  NAND2XL U30098 ( .A(n24666), .B(n24665), .Y(n24734) );
  INVXL U30099 ( .A(n24734), .Y(n24667) );
  AOI21X2 U30100 ( .A0(n24671), .A1(n24729), .B0(n24670), .Y(n24672) );
  INVXL U30101 ( .A(n24674), .Y(n24678) );
  NOR2XL U30102 ( .A(n24679), .B(n24678), .Y(n24724) );
  INVXL U30103 ( .A(n24676), .Y(n24685) );
  NAND2X1 U30104 ( .A(n24679), .B(n24678), .Y(n24725) );
  NAND2XL U30105 ( .A(n24681), .B(n24680), .Y(n24682) );
  OAI21XL U30106 ( .A0(n24725), .A1(n24683), .B0(n24682), .Y(n24711) );
  NAND2XL U30107 ( .A(n24688), .B(n24687), .Y(n24689) );
  MXI2X1 U30108 ( .A(U0_pipe3[27]), .B(n24695), .S0(n5812), .Y(n4348) );
  MXI2X1 U30109 ( .A(U0_pipe3[26]), .B(n24697), .S0(n5812), .Y(n4349) );
  XOR2X1 U30110 ( .A(n24699), .B(n24698), .Y(n24700) );
  CLKINVX3 U30111 ( .A(n5837), .Y(n25273) );
  MXI2X1 U30112 ( .A(U0_pipe3[25]), .B(n24700), .S0(n25273), .Y(n4350) );
  OAI21XL U30113 ( .A0(n24727), .A1(n24703), .B0(n24702), .Y(n24708) );
  INVXL U30114 ( .A(n24704), .Y(n24706) );
  INVXL U30115 ( .A(n24990), .Y(n24707) );
  INVXL U30116 ( .A(n24710), .Y(n24713) );
  INVXL U30117 ( .A(n24711), .Y(n24712) );
  OAI21XL U30118 ( .A0(n24727), .A1(n24713), .B0(n24712), .Y(n24718) );
  NAND2XL U30119 ( .A(n5849), .B(n24725), .Y(n24726) );
  AOI21X1 U30120 ( .A0(n24773), .A1(n24730), .B0(n24729), .Y(n24742) );
  XOR2X1 U30121 ( .A(n24736), .B(n25012), .Y(n24737) );
  NAND2XL U30122 ( .A(n24739), .B(n24738), .Y(n25014) );
  XNOR2XL U30123 ( .A(n24740), .B(n25014), .Y(n24741) );
  NAND2XL U30124 ( .A(n5794), .B(n24748), .Y(n24749) );
  OAI21XL U30125 ( .A0(n24764), .A1(n24756), .B0(n24761), .Y(n24759) );
  XNOR2X1 U30126 ( .A(n24759), .B(n25032), .Y(n24760) );
  MXI2X1 U30127 ( .A(U0_pipe3[16]), .B(n24760), .S0(n25273), .Y(n4359) );
  NAND2XL U30128 ( .A(n24762), .B(n24761), .Y(n24763) );
  AOI21XL U30129 ( .A0(n24773), .A1(n24648), .B0(n24766), .Y(n24769) );
  CLKINVX3 U30130 ( .A(n5837), .Y(n25091) );
  INVXL U30131 ( .A(n24775), .Y(n24808) );
  OAI21XL U30132 ( .A0(n24808), .A1(n24777), .B0(n24776), .Y(n24788) );
  NAND2XL U30133 ( .A(n9004), .B(n24786), .Y(n25055) );
  OAI21XL U30134 ( .A0(n24808), .A1(n24791), .B0(n24790), .Y(n24804) );
  INVXL U30135 ( .A(n24792), .Y(n24795) );
  INVXL U30136 ( .A(n24793), .Y(n24794) );
  NAND2XL U30137 ( .A(n24806), .B(n25058), .Y(n25069) );
  OAI21XL U30138 ( .A0(n24841), .A1(n24832), .B0(n24831), .Y(n24837) );
  XOR2XL U30139 ( .A(n24845), .B(n24844), .Y(n24846) );
  XOR2XL U30140 ( .A(n24849), .B(n24848), .Y(n24850) );
  XNOR2XL U30141 ( .A(n24852), .B(n24851), .Y(n25114) );
  OAI21XL U30142 ( .A0(n24862), .A1(n24861), .B0(n24860), .Y(n24863) );
  MXI2X1 U30143 ( .A(U0_pipe0[27]), .B(n24864), .S0(n24784), .Y(n4285) );
  XNOR2X1 U30144 ( .A(n24868), .B(n24867), .Y(n24869) );
  MXI2X1 U30145 ( .A(U0_pipe0[25]), .B(n24869), .S0(n24784), .Y(n4287) );
  XOR2X1 U30146 ( .A(n24871), .B(n24870), .Y(n24872) );
  OAI21XL U30147 ( .A0(n24885), .A1(n24875), .B0(n24874), .Y(n24877) );
  XNOR2X1 U30148 ( .A(n24877), .B(n24876), .Y(n24878) );
  MXI2X1 U30149 ( .A(U0_pipe0[23]), .B(n24878), .S0(n24784), .Y(n4289) );
  OAI21XL U30150 ( .A0(n24885), .A1(n24880), .B0(n24879), .Y(n24882) );
  XNOR2X1 U30151 ( .A(n24882), .B(n24881), .Y(n24883) );
  MXI2X1 U30152 ( .A(U0_pipe0[22]), .B(n24883), .S0(n24784), .Y(n4290) );
  XOR2X1 U30153 ( .A(n24885), .B(n24884), .Y(n24886) );
  XOR2X1 U30154 ( .A(n24888), .B(n24887), .Y(n24889) );
  OAI21XL U30155 ( .A0(n24892), .A1(n24891), .B0(n24890), .Y(n24894) );
  XNOR2X1 U30156 ( .A(n24897), .B(n24896), .Y(n24898) );
  INVXL U30157 ( .A(n24900), .Y(n24901) );
  OAI21XL U30158 ( .A0(n24909), .A1(n24904), .B0(n24903), .Y(n24906) );
  XNOR2XL U30159 ( .A(n24906), .B(n24905), .Y(n24907) );
  AOI21XL U30160 ( .A0(n24917), .A1(n24912), .B0(n24911), .Y(n24914) );
  OAI21XL U30161 ( .A0(n24941), .A1(n24921), .B0(n24920), .Y(n24927) );
  AOI21XL U30162 ( .A0(n24927), .A1(n13507), .B0(n24922), .Y(n24924) );
  OAI21XL U30163 ( .A0(n24941), .A1(n24930), .B0(n24929), .Y(n24938) );
  INVXL U30164 ( .A(n24931), .Y(n24932) );
  INVXL U30165 ( .A(n24943), .Y(n24962) );
  AOI21XL U30166 ( .A0(n24962), .A1(n24945), .B0(n24944), .Y(n24949) );
  INVXL U30167 ( .A(n24953), .Y(n24955) );
  OAI21XL U30168 ( .A0(n24975), .A1(n24971), .B0(n24972), .Y(n24969) );
  INVXL U30169 ( .A(n24965), .Y(n24967) );
  XOR2XL U30170 ( .A(n24981), .B(n24980), .Y(n24982) );
  XNOR2XL U30171 ( .A(n24984), .B(n24983), .Y(n24985) );
  OAI21XL U30172 ( .A0(n25004), .A1(n24993), .B0(n24992), .Y(n24995) );
  OAI21XL U30173 ( .A0(n25004), .A1(n24997), .B0(n25001), .Y(n24999) );
  NAND2XL U30174 ( .A(n25002), .B(n25001), .Y(n25003) );
  XNOR2X1 U30175 ( .A(n25022), .B(n25021), .Y(n25023) );
  INVXL U30176 ( .A(n25027), .Y(n25030) );
  INVXL U30177 ( .A(n25028), .Y(n25029) );
  NAND2XL U30178 ( .A(n25034), .B(n25033), .Y(n25035) );
  AOI21XL U30179 ( .A0(n25046), .A1(n9136), .B0(n25038), .Y(n25042) );
  NAND2XL U30180 ( .A(n9136), .B(n25044), .Y(n25045) );
  OAI21XL U30181 ( .A0(n25070), .A1(n25050), .B0(n25049), .Y(n25056) );
  AOI21XL U30182 ( .A0(n25056), .A1(n9004), .B0(n25051), .Y(n25053) );
  INVXL U30183 ( .A(n25060), .Y(n25061) );
  AOI21XL U30184 ( .A0(n25090), .A1(n25074), .B0(n25073), .Y(n25077) );
  INVXL U30185 ( .A(n25081), .Y(n25083) );
  OAI21XL U30186 ( .A0(n25104), .A1(n25095), .B0(n25094), .Y(n25100) );
  INVXL U30187 ( .A(n25096), .Y(n25098) );
  OAI21XL U30188 ( .A0(n25111), .A1(n25107), .B0(n25106), .Y(n25109) );
  XOR2XL U30189 ( .A(n25112), .B(n25111), .Y(n25113) );
  NAND2XL U30190 ( .A(U0_pipe1[0]), .B(U0_pipe0[0]), .Y(n25116) );
  OAI21XL U30191 ( .A0(n25117), .A1(n25116), .B0(n25115), .Y(n25866) );
  CMPR32X1 U30192 ( .A(n25123), .B(n29010), .C(n25122), .CO(n14498), .S(n25124) );
  MXI2X1 U30193 ( .A(U0_pipe12[26]), .B(n25124), .S0(n5810), .Y(n4694) );
  NAND2XL U30194 ( .A(n25125), .B(U2_A_r_d[25]), .Y(n25524) );
  XOR2X1 U30195 ( .A(n25127), .B(n25126), .Y(n25128) );
  OAI21XL U30196 ( .A0(n25153), .A1(n25131), .B0(n25130), .Y(n25135) );
  INVXL U30197 ( .A(n25523), .Y(n25133) );
  INVXL U30198 ( .A(n25533), .Y(n25134) );
  XNOR2X1 U30199 ( .A(n25135), .B(n25134), .Y(n25136) );
  MXI2X1 U30200 ( .A(U0_pipe12[24]), .B(n25136), .S0(n5810), .Y(n4696) );
  OAI21XL U30201 ( .A0(n25153), .A1(n25139), .B0(n25138), .Y(n25143) );
  INVXL U30202 ( .A(n25519), .Y(n25141) );
  NAND2XL U30203 ( .A(n25140), .B(U2_A_r_d[23]), .Y(n25518) );
  XNOR2X1 U30204 ( .A(n25143), .B(n25142), .Y(n25144) );
  MXI2X1 U30205 ( .A(U0_pipe12[23]), .B(n25144), .S0(n5810), .Y(n4697) );
  OAI21XL U30206 ( .A0(n25153), .A1(n25146), .B0(n25145), .Y(n25149) );
  OR2X2 U30207 ( .A(n25147), .B(U2_A_r_d[22]), .Y(n25516) );
  NAND2XL U30208 ( .A(n25147), .B(U2_A_r_d[22]), .Y(n25514) );
  XNOR2X1 U30209 ( .A(n25149), .B(n25148), .Y(n25150) );
  MXI2X1 U30210 ( .A(U0_pipe12[22]), .B(n25150), .S0(n5810), .Y(n4698) );
  NOR2XL U30211 ( .A(n25151), .B(U2_A_r_d[21]), .Y(n25543) );
  INVXL U30212 ( .A(n25543), .Y(n25513) );
  NAND2XL U30213 ( .A(n25151), .B(U2_A_r_d[21]), .Y(n25542) );
  XOR2X1 U30214 ( .A(n25153), .B(n25152), .Y(n25154) );
  AOI21X1 U30215 ( .A0(n25205), .A1(n25157), .B0(n25156), .Y(n25170) );
  NAND2XL U30216 ( .A(n25162), .B(U2_A_r_d[20]), .Y(n25504) );
  NAND2XL U30217 ( .A(n6948), .B(n25504), .Y(n25559) );
  XOR2X1 U30218 ( .A(n25164), .B(n25163), .Y(n25165) );
  MXI2X1 U30219 ( .A(U0_pipe12[20]), .B(n25165), .S0(n5810), .Y(n4700) );
  NOR2XL U30220 ( .A(n25166), .B(U2_A_r_d[19]), .Y(n25558) );
  INVXL U30221 ( .A(n25558), .Y(n25488) );
  NAND2XL U30222 ( .A(n25166), .B(U2_A_r_d[19]), .Y(n25557) );
  NAND2XL U30223 ( .A(n25488), .B(n25557), .Y(n25562) );
  INVXL U30224 ( .A(n25170), .Y(n25180) );
  AOI21XL U30225 ( .A0(n25180), .A1(n25172), .B0(n25171), .Y(n25176) );
  NOR2XL U30226 ( .A(n25174), .B(U2_A_r_d[18]), .Y(n25173) );
  NAND2XL U30227 ( .A(n25174), .B(U2_A_r_d[18]), .Y(n25500) );
  NAND2XL U30228 ( .A(n25503), .B(n25500), .Y(n25568) );
  XOR2X1 U30229 ( .A(n25176), .B(n25175), .Y(n25177) );
  NOR2XL U30230 ( .A(n25178), .B(U2_A_r_d[17]), .Y(n25566) );
  INVXL U30231 ( .A(n25566), .Y(n25489) );
  NAND2XL U30232 ( .A(n25178), .B(U2_A_r_d[17]), .Y(n25565) );
  NAND2XL U30233 ( .A(n25489), .B(n25565), .Y(n25571) );
  OAI21XL U30234 ( .A0(n25195), .A1(n25187), .B0(n25186), .Y(n25191) );
  NOR2XL U30235 ( .A(n25189), .B(U2_A_r_d[16]), .Y(n25188) );
  NAND2XL U30236 ( .A(n25189), .B(U2_A_r_d[16]), .Y(n25494) );
  NAND2XL U30237 ( .A(n25497), .B(n25494), .Y(n25580) );
  XNOR2X1 U30238 ( .A(n25191), .B(n25190), .Y(n25192) );
  NOR2XL U30239 ( .A(n25193), .B(U2_A_r_d[15]), .Y(n25579) );
  INVXL U30240 ( .A(n25579), .Y(n25487) );
  NAND2XL U30241 ( .A(n25193), .B(U2_A_r_d[15]), .Y(n25578) );
  AOI21XL U30242 ( .A0(n25205), .A1(n25198), .B0(n25197), .Y(n25201) );
  NAND2XL U30243 ( .A(n25199), .B(U2_A_r_d[14]), .Y(n25491) );
  OR2X1 U30244 ( .A(n25203), .B(U2_A_r_d[13]), .Y(n25587) );
  NAND2XL U30245 ( .A(n25203), .B(U2_A_r_d[13]), .Y(n25490) );
  OAI21XL U30246 ( .A0(n25237), .A1(n25209), .B0(n25208), .Y(n25218) );
  NAND2XL U30247 ( .A(n25212), .B(U2_A_r_d[12]), .Y(n25481) );
  NAND2XL U30248 ( .A(n5775), .B(n25480), .Y(n25601) );
  OAI21XL U30249 ( .A0(n25237), .A1(n25221), .B0(n25220), .Y(n25233) );
  NOR2X2 U30250 ( .A(n25226), .B(U2_A_r_d[10]), .Y(n25476) );
  INVXL U30251 ( .A(n25476), .Y(n25227) );
  NAND2XL U30252 ( .A(n25226), .B(U2_A_r_d[10]), .Y(n25475) );
  NAND2XL U30253 ( .A(n25227), .B(n25475), .Y(n25609) );
  NOR2XL U30254 ( .A(n25231), .B(U2_A_r_d[9]), .Y(n25473) );
  NAND2XL U30255 ( .A(n25231), .B(U2_A_r_d[9]), .Y(n25606) );
  NOR2XL U30256 ( .A(n25235), .B(U2_A_r_d[8]), .Y(n25605) );
  INVXL U30257 ( .A(n25605), .Y(n25474) );
  NAND2XL U30258 ( .A(n25235), .B(U2_A_r_d[8]), .Y(n25604) );
  NAND2XL U30259 ( .A(n25474), .B(n25604), .Y(n25616) );
  AOI21XL U30260 ( .A0(n25258), .A1(n25241), .B0(n25240), .Y(n25245) );
  NAND2XL U30261 ( .A(n25243), .B(U2_A_r_d[7]), .Y(n25469) );
  INVXL U30262 ( .A(n25468), .Y(n25252) );
  NAND2XL U30263 ( .A(n25251), .B(U2_A_r_d[6]), .Y(n25467) );
  NAND2XL U30264 ( .A(n25252), .B(n25467), .Y(n25628) );
  NOR2XL U30265 ( .A(n25256), .B(U2_A_r_d[5]), .Y(n25457) );
  NAND2XL U30266 ( .A(n25256), .B(U2_A_r_d[5]), .Y(n25625) );
  OAI21XL U30267 ( .A0(n25272), .A1(n25262), .B0(n25261), .Y(n25266) );
  NOR2XL U30268 ( .A(n25263), .B(U2_A_r_d[4]), .Y(n25464) );
  INVXL U30269 ( .A(n25464), .Y(n25264) );
  NAND2XL U30270 ( .A(n25263), .B(U2_A_r_d[4]), .Y(n25463) );
  NOR2XL U30271 ( .A(n25269), .B(U2_A_r_d[3]), .Y(n25636) );
  NAND2XL U30272 ( .A(n25269), .B(U2_A_r_d[3]), .Y(n25635) );
  NOR2XL U30273 ( .A(n25275), .B(U2_A_r_d[2]), .Y(n25462) );
  NAND2XL U30274 ( .A(n25275), .B(U2_A_r_d[2]), .Y(n25461) );
  XOR2XL U30275 ( .A(n25278), .B(n25277), .Y(n25279) );
  NAND2XL U30276 ( .A(n25281), .B(U2_A_r_d[1]), .Y(n25459) );
  XOR2XL U30277 ( .A(n25283), .B(n25282), .Y(n25284) );
  XNOR2XL U30278 ( .A(n25285), .B(U2_A_r_d[0]), .Y(n25649) );
  MXI2X1 U30279 ( .A(U0_pipe13[27]), .B(n25287), .S0(n25318), .Y(n4665) );
  MXI2X1 U30280 ( .A(U0_pipe13[25]), .B(n25288), .S0(n25318), .Y(n4667) );
  OAI21XL U30281 ( .A0(n25317), .A1(n25291), .B0(n25290), .Y(n25296) );
  NAND2X1 U30282 ( .A(n25294), .B(n25293), .Y(n25660) );
  XNOR2X1 U30283 ( .A(n25296), .B(n25295), .Y(n25297) );
  MXI2X1 U30284 ( .A(U0_pipe13[20]), .B(n25331), .S0(U1_valid[0]), .Y(n4672)
         );
  XNOR2X1 U30285 ( .A(n25334), .B(n25333), .Y(n25335) );
  MXI2X1 U30286 ( .A(U0_pipe13[18]), .B(n25342), .S0(U1_valid[0]), .Y(n4674)
         );
  INVXL U30287 ( .A(n25347), .Y(n25350) );
  INVXL U30288 ( .A(n25348), .Y(n25349) );
  OAI21XL U30289 ( .A0(n25360), .A1(n25351), .B0(n25357), .Y(n25355) );
  NAND2XL U30290 ( .A(n25353), .B(n25352), .Y(n25354) );
  XNOR2X1 U30291 ( .A(n25355), .B(n25354), .Y(n25356) );
  NAND2XL U30292 ( .A(n25358), .B(n25357), .Y(n25359) );
  AOI21XL U30293 ( .A0(n25370), .A1(n12385), .B0(n25362), .Y(n25366) );
  NAND2XL U30294 ( .A(n12385), .B(n25368), .Y(n25369) );
  INVXL U30295 ( .A(n25372), .Y(n25402) );
  OAI21XL U30296 ( .A0(n25402), .A1(n25374), .B0(n25373), .Y(n25383) );
  AOI21XL U30297 ( .A0(n25383), .A1(n6992), .B0(n25375), .Y(n25379) );
  NAND2XL U30298 ( .A(n6992), .B(n25381), .Y(n25382) );
  OAI21XL U30299 ( .A0(n25402), .A1(n25386), .B0(n25385), .Y(n25398) );
  AOI21XL U30300 ( .A0(n25398), .A1(n25396), .B0(n25388), .Y(n25393) );
  INVXL U30301 ( .A(n25389), .Y(n25391) );
  NAND2XL U30302 ( .A(n25400), .B(n25737), .Y(n25752) );
  CLKINVX3 U30303 ( .A(n17032), .Y(n25611) );
  OAI21XL U30304 ( .A0(n25435), .A1(n25426), .B0(n25425), .Y(n25431) );
  INVXL U30305 ( .A(n25427), .Y(n25429) );
  XOR2XL U30306 ( .A(n25441), .B(n25440), .Y(n25442) );
  XOR2XL U30307 ( .A(n25446), .B(n25445), .Y(n25447) );
  XNOR2XL U30308 ( .A(n25449), .B(n25448), .Y(n25791) );
  NOR2XL U30309 ( .A(n25468), .B(n25457), .Y(n25621) );
  NAND2XL U30310 ( .A(n25621), .B(n25242), .Y(n25472) );
  NOR2XL U30311 ( .A(n25464), .B(n25636), .Y(n25466) );
  INVXL U30312 ( .A(n25459), .Y(n25460) );
  AOI21XL U30313 ( .A0(n25646), .A1(n25280), .B0(n25460), .Y(n25643) );
  OAI21XL U30314 ( .A0(n25643), .A1(n25462), .B0(n25461), .Y(n25634) );
  OAI21XL U30315 ( .A0(n25464), .A1(n25635), .B0(n25463), .Y(n25465) );
  AOI21XL U30316 ( .A0(n25466), .A1(n25634), .B0(n25465), .Y(n25619) );
  OAI21XL U30317 ( .A0(n25468), .A1(n25625), .B0(n25467), .Y(n25620) );
  INVXL U30318 ( .A(n25469), .Y(n25470) );
  OAI21XL U30319 ( .A0(n25472), .A1(n25619), .B0(n25471), .Y(n25594) );
  NOR2XL U30320 ( .A(n25476), .B(n25473), .Y(n25479) );
  NAND2XL U30321 ( .A(n25479), .B(n25474), .Y(n25596) );
  NOR2XL U30322 ( .A(n25596), .B(n25484), .Y(n25486) );
  INVXL U30323 ( .A(n25604), .Y(n25478) );
  OAI21XL U30324 ( .A0(n25476), .A1(n25606), .B0(n25475), .Y(n25477) );
  AOI21XL U30325 ( .A0(n25479), .A1(n25478), .B0(n25477), .Y(n25595) );
  INVXL U30326 ( .A(n25480), .Y(n25597) );
  INVXL U30327 ( .A(n25481), .Y(n25482) );
  NAND2XL U30328 ( .A(n25497), .B(n25487), .Y(n25499) );
  NAND2XL U30329 ( .A(n25493), .B(n25587), .Y(n25574) );
  NOR2XL U30330 ( .A(n25499), .B(n25574), .Y(n25552) );
  NAND2X1 U30331 ( .A(n25503), .B(n25489), .Y(n25553) );
  NOR2X1 U30332 ( .A(n25508), .B(n25553), .Y(n25510) );
  INVXL U30333 ( .A(n25490), .Y(n25586) );
  INVXL U30334 ( .A(n25491), .Y(n25492) );
  AOI21XL U30335 ( .A0(n25493), .A1(n25586), .B0(n25492), .Y(n25575) );
  INVXL U30336 ( .A(n25578), .Y(n25496) );
  INVXL U30337 ( .A(n25494), .Y(n25495) );
  AOI21XL U30338 ( .A0(n25497), .A1(n25496), .B0(n25495), .Y(n25498) );
  OAI21XL U30339 ( .A0(n25499), .A1(n25575), .B0(n25498), .Y(n25551) );
  INVXL U30340 ( .A(n25565), .Y(n25502) );
  INVXL U30341 ( .A(n25500), .Y(n25501) );
  INVXL U30342 ( .A(n25557), .Y(n25506) );
  INVXL U30343 ( .A(n25504), .Y(n25505) );
  AOI21X1 U30344 ( .A0(n25551), .A1(n25510), .B0(n25509), .Y(n25511) );
  OAI21X2 U30345 ( .A0(n25550), .A1(n25512), .B0(n25511), .Y(n25536) );
  NAND2XL U30346 ( .A(n25513), .B(n25516), .Y(n25538) );
  INVXL U30347 ( .A(n25542), .Y(n25517) );
  INVXL U30348 ( .A(n25514), .Y(n25515) );
  OAI21X1 U30349 ( .A0(n25537), .A1(n25519), .B0(n25518), .Y(n25520) );
  INVXL U30350 ( .A(n25524), .Y(n25525) );
  MXI2X1 U30351 ( .A(U0_pipe8[27]), .B(n25527), .S0(n5812), .Y(n4606) );
  MXI2X1 U30352 ( .A(U0_pipe8[26]), .B(n25529), .S0(n5812), .Y(n4607) );
  XNOR2X1 U30353 ( .A(n25531), .B(n25530), .Y(n25532) );
  MXI2X1 U30354 ( .A(U0_pipe8[24]), .B(n25535), .S0(n5812), .Y(n4410) );
  INVXL U30355 ( .A(n25536), .Y(n25548) );
  OAI21XL U30356 ( .A0(n25548), .A1(n25538), .B0(n25537), .Y(n25540) );
  XNOR2XL U30357 ( .A(n25540), .B(n25539), .Y(n25541) );
  OAI21XL U30358 ( .A0(n25548), .A1(n25543), .B0(n25542), .Y(n25545) );
  XNOR2XL U30359 ( .A(n25545), .B(n25544), .Y(n25546) );
  INVXL U30360 ( .A(n25554), .Y(n25555) );
  OAI21XL U30361 ( .A0(n25567), .A1(n25566), .B0(n25565), .Y(n25569) );
  INVXL U30362 ( .A(n25575), .Y(n25576) );
  OAI21XL U30363 ( .A0(n25584), .A1(n25579), .B0(n25578), .Y(n25581) );
  OAI21XL U30364 ( .A0(n25617), .A1(n25596), .B0(n25595), .Y(n25602) );
  AOI21XL U30365 ( .A0(n25602), .A1(n5775), .B0(n25597), .Y(n25599) );
  OAI21XL U30366 ( .A0(n25617), .A1(n25605), .B0(n25604), .Y(n25614) );
  INVXL U30367 ( .A(n25619), .Y(n25632) );
  AOI21XL U30368 ( .A0(n25632), .A1(n25621), .B0(n25620), .Y(n25623) );
  OAI21XL U30369 ( .A0(n25641), .A1(n25636), .B0(n25635), .Y(n25638) );
  XOR2XL U30370 ( .A(n25644), .B(n25643), .Y(n25645) );
  XNOR2XL U30371 ( .A(n25647), .B(n25646), .Y(n25648) );
  INVXL U30372 ( .A(n25650), .Y(n25651) );
  MXI2X1 U30373 ( .A(U0_pipe9[27]), .B(n25655), .S0(n6888), .Y(n4578) );
  MXI2X1 U30374 ( .A(U0_pipe9[26]), .B(n25659), .S0(n5812), .Y(n4579) );
  XOR2X1 U30375 ( .A(n25661), .B(n25660), .Y(n25662) );
  MXI2X1 U30376 ( .A(U0_pipe9[24]), .B(n25662), .S0(n5812), .Y(n4581) );
  OAI21XL U30377 ( .A0(n25675), .A1(n25665), .B0(n25664), .Y(n25667) );
  XNOR2X1 U30378 ( .A(n25667), .B(n25666), .Y(n25668) );
  MXI2X1 U30379 ( .A(U0_pipe9[23]), .B(n25668), .S0(n6888), .Y(n4582) );
  OAI21XL U30380 ( .A0(n25675), .A1(n25670), .B0(n25669), .Y(n25672) );
  XNOR2X1 U30381 ( .A(n25672), .B(n25671), .Y(n25673) );
  MXI2X1 U30382 ( .A(U0_pipe9[22]), .B(n25673), .S0(n6888), .Y(n4583) );
  XOR2X1 U30383 ( .A(n25675), .B(n25674), .Y(n25676) );
  INVX2 U30384 ( .A(n25677), .Y(n25722) );
  INVXL U30385 ( .A(n25681), .Y(n25682) );
  XNOR2X1 U30386 ( .A(n25686), .B(n25685), .Y(n25687) );
  OAI21XL U30387 ( .A0(n25693), .A1(n25692), .B0(n25691), .Y(n25695) );
  XNOR2XL U30388 ( .A(n25695), .B(n25694), .Y(n25696) );
  INVXL U30389 ( .A(n25699), .Y(n25702) );
  OAI21XL U30390 ( .A0(n25712), .A1(n25703), .B0(n25709), .Y(n25707) );
  NAND2XL U30391 ( .A(n25705), .B(n25704), .Y(n25706) );
  NAND2XL U30392 ( .A(n25710), .B(n25709), .Y(n25711) );
  AOI21XL U30393 ( .A0(n25722), .A1(n12204), .B0(n25714), .Y(n25718) );
  NAND2XL U30394 ( .A(n25716), .B(n25715), .Y(n25717) );
  NAND2XL U30395 ( .A(n12204), .B(n25720), .Y(n25721) );
  OAI21XL U30396 ( .A0(n25753), .A1(n25725), .B0(n25724), .Y(n25735) );
  AOI21XL U30397 ( .A0(n25735), .A1(n25733), .B0(n25726), .Y(n25730) );
  NAND2XL U30398 ( .A(n25733), .B(n25732), .Y(n25734) );
  OAI21XL U30399 ( .A0(n25753), .A1(n25738), .B0(n25737), .Y(n25750) );
  INVXL U30400 ( .A(n25739), .Y(n25748) );
  INVXL U30401 ( .A(n25747), .Y(n25740) );
  AOI21XL U30402 ( .A0(n25750), .A1(n25748), .B0(n25740), .Y(n25745) );
  NAND2XL U30403 ( .A(n25748), .B(n25747), .Y(n25749) );
  AOI21XL U30404 ( .A0(n25773), .A1(n25757), .B0(n25756), .Y(n25760) );
  OAI21XL U30405 ( .A0(n25782), .A1(n25777), .B0(n25776), .Y(n25779) );
  XOR2XL U30406 ( .A(n25785), .B(n25784), .Y(n25786) );
  XNOR2XL U30407 ( .A(n25789), .B(n25788), .Y(n25790) );
  OR2XL U30408 ( .A(n28904), .B(U0_pipe8[0]), .Y(n25795) );
  OAI21XL U30409 ( .A0(n25845), .A1(n25799), .B0(n25838), .Y(n25804) );
  NOR2XL U30410 ( .A(n25802), .B(U2_A_r_d[1]), .Y(n25801) );
  INVXL U30411 ( .A(n25801), .Y(n25842) );
  NAND2XL U30412 ( .A(n25802), .B(U2_A_r_d[1]), .Y(n25839) );
  OAI21XL U30413 ( .A0(n25808), .A1(n25807), .B0(n25806), .Y(n25930) );
  CMPR22X1 U30414 ( .A(U0_pipe2[2]), .B(n28721), .CO(n25810), .S(n24853) );
  OAI21XL U30415 ( .A0(n25814), .A1(n25861), .B0(n25863), .Y(n25819) );
  CMPR22X1 U30416 ( .A(U0_pipe1[2]), .B(U0_pipe0[2]), .CO(n25816), .S(n25118)
         );
  OAI21XL U30417 ( .A0(n25823), .A1(n25822), .B0(n25821), .Y(n25919) );
  CMPR22X1 U30418 ( .A(U0_pipe12[2]), .B(n28745), .CO(n25825), .S(n25450) );
  OAI21XL U30419 ( .A0(n25831), .A1(n25830), .B0(n25829), .Y(n25900) );
  CMPR22X1 U30420 ( .A(U0_pipe8[2]), .B(n28717), .CO(n25833), .S(n25792) );
  NAND2XL U30421 ( .A(n25842), .B(n25837), .Y(n25844) );
  INVXL U30422 ( .A(n25839), .Y(n25840) );
  AOI21XL U30423 ( .A0(n25842), .A1(n25841), .B0(n25840), .Y(n25843) );
  OAI21XL U30424 ( .A0(n25845), .A1(n25844), .B0(n25843), .Y(n25942) );
  CMPR32X1 U30425 ( .A(n25848), .B(n25847), .C(n25846), .CO(n25849), .S(n25802) );
  NOR2XL U30426 ( .A(n25850), .B(n25849), .Y(n25936) );
  OAI21XL U30427 ( .A0(n25854), .A1(n25895), .B0(n25897), .Y(n25859) );
  CMPR22X1 U30428 ( .A(U0_pipe8[3]), .B(n28716), .CO(n25856), .S(n25832) );
  OAI21XL U30429 ( .A0(n25864), .A1(n25863), .B0(n25862), .Y(n25865) );
  CMPR22X1 U30430 ( .A(U0_pipe1[3]), .B(U0_pipe0[3]), .CO(n25869), .S(n25815)
         );
  OAI21XL U30431 ( .A0(n25872), .A1(n25914), .B0(n25916), .Y(n25877) );
  CMPR22X1 U30432 ( .A(U0_pipe12[3]), .B(n28724), .CO(n25874), .S(n25824) );
  OAI21XL U30433 ( .A0(n25879), .A1(n25925), .B0(n25927), .Y(n25884) );
  CMPR22X1 U30434 ( .A(U0_pipe2[3]), .B(n28720), .CO(n25881), .S(n25809) );
  OAI21XL U30435 ( .A0(n25886), .A1(n25936), .B0(n25938), .Y(n25893) );
  CMPR32X1 U30436 ( .A(n25888), .B(n25887), .C(U2_A_r_d[2]), .CO(n25889), .S(
        n25850) );
  OAI21XL U30437 ( .A0(n25898), .A1(n25897), .B0(n25896), .Y(n25899) );
  CMPR22X1 U30438 ( .A(U0_pipe8[4]), .B(n28775), .CO(n25903), .S(n25855) );
  CMPR22X1 U30439 ( .A(U0_pipe1[4]), .B(U0_pipe0[4]), .CO(n25909), .S(n25868)
         );
  OAI21XL U30440 ( .A0(n25917), .A1(n25916), .B0(n25915), .Y(n25918) );
  CMPR22X1 U30441 ( .A(U0_pipe12[4]), .B(n28807), .CO(n25922), .S(n25873) );
  OAI21XL U30442 ( .A0(n25928), .A1(n25927), .B0(n25926), .Y(n25929) );
  CMPR22X1 U30443 ( .A(U0_pipe2[4]), .B(n28791), .CO(n25933), .S(n25880) );
  NOR2XL U30444 ( .A(n25936), .B(n25939), .Y(n25941) );
  OAI21XL U30445 ( .A0(n25939), .A1(n25938), .B0(n25937), .Y(n25940) );
  AOI21XL U30446 ( .A0(n25942), .A1(n25941), .B0(n25940), .Y(n26152) );
  NAND2XL U30447 ( .A(n25946), .B(n25945), .Y(n26032) );
  CMPR22X1 U30448 ( .A(U0_pipe8[5]), .B(n28774), .CO(n25952), .S(n25902) );
  OAI21XL U30449 ( .A0(n25960), .A1(n25959), .B0(n25958), .Y(n26055) );
  CMPR22X1 U30450 ( .A(U0_pipe1[5]), .B(U0_pipe0[5]), .CO(n25963), .S(n25908)
         );
  NAND2XL U30451 ( .A(n25964), .B(n26052), .Y(n25965) );
  CMPR22X1 U30452 ( .A(U0_pipe12[5]), .B(n28806), .CO(n25970), .S(n25921) );
  CMPR22X1 U30453 ( .A(U0_pipe2[5]), .B(n28790), .CO(n25978), .S(n25932) );
  NAND2XL U30454 ( .A(n25988), .B(n25987), .Y(n26031) );
  OAI21XL U30455 ( .A0(n25996), .A1(n25995), .B0(n25994), .Y(n26132) );
  CMPR22X1 U30456 ( .A(U0_pipe2[6]), .B(n28719), .CO(n25999), .S(n25977) );
  OAI21XL U30457 ( .A0(n26003), .A1(n26049), .B0(n26052), .Y(n26008) );
  CMPR22X1 U30458 ( .A(U0_pipe1[6]), .B(U0_pipe0[6]), .CO(n26005), .S(n25962)
         );
  OAI21XL U30459 ( .A0(n26013), .A1(n26012), .B0(n26011), .Y(n26116) );
  CMPR22X1 U30460 ( .A(U0_pipe12[6]), .B(n28723), .CO(n26016), .S(n25969) );
  OAI21XL U30461 ( .A0(n26023), .A1(n26022), .B0(n26021), .Y(n26094) );
  CMPR22X1 U30462 ( .A(U0_pipe8[6]), .B(n28715), .CO(n26026), .S(n25951) );
  NOR2XL U30463 ( .A(n26030), .B(n26033), .Y(n26143) );
  OAI21XL U30464 ( .A0(n26033), .A1(n26032), .B0(n26031), .Y(n26148) );
  CMPR32X1 U30465 ( .A(n26036), .B(n26035), .C(U2_A_r_d[5]), .CO(n26037), .S(
        n25988) );
  NAND2XL U30466 ( .A(n26038), .B(n26037), .Y(n26145) );
  OAI21XL U30467 ( .A0(n26042), .A1(n26126), .B0(n26129), .Y(n26047) );
  CMPR22X1 U30468 ( .A(U0_pipe2[7]), .B(n28789), .CO(n26044), .S(n25998) );
  OAI21XL U30469 ( .A0(n26053), .A1(n26052), .B0(n26051), .Y(n26054) );
  OAI21XL U30470 ( .A0(n26059), .A1(n26058), .B0(n26057), .Y(n26498) );
  CMPR22X1 U30471 ( .A(U0_pipe1[7]), .B(U0_pipe0[7]), .CO(n26061), .S(n26004)
         );
  OAI21XL U30472 ( .A0(n26065), .A1(n26110), .B0(n26113), .Y(n26070) );
  CMPR22X1 U30473 ( .A(U0_pipe12[7]), .B(n28805), .CO(n26067), .S(n26015) );
  OAI21XL U30474 ( .A0(n26072), .A1(n26088), .B0(n26091), .Y(n26077) );
  CMPR22X1 U30475 ( .A(U0_pipe8[7]), .B(n28773), .CO(n26074), .S(n26025) );
  OAI21XL U30476 ( .A0(n26079), .A1(n26142), .B0(n26145), .Y(n26086) );
  CMPR32X1 U30477 ( .A(n26081), .B(n26080), .C(U2_A_r_d[6]), .CO(n26082), .S(
        n26038) );
  INVXL U30478 ( .A(n26146), .Y(n26084) );
  NAND2XL U30479 ( .A(n26083), .B(n26082), .Y(n26144) );
  OAI21XL U30480 ( .A0(n26092), .A1(n26091), .B0(n26090), .Y(n26093) );
  OAI21XL U30481 ( .A0(n26098), .A1(n26097), .B0(n26096), .Y(n26585) );
  CMPR22X1 U30482 ( .A(U0_pipe8[8]), .B(n28772), .CO(n26100), .S(n26073) );
  NAND2XL U30483 ( .A(n26101), .B(n26198), .Y(n26102) );
  OAI21XL U30484 ( .A0(n26264), .A1(n26166), .B0(n26168), .Y(n26108) );
  CMPR22X1 U30485 ( .A(U0_pipe1[8]), .B(U0_pipe0[8]), .CO(n26105), .S(n26060)
         );
  OAI21XL U30486 ( .A0(n26114), .A1(n26113), .B0(n26112), .Y(n26115) );
  OAI21XL U30487 ( .A0(n26120), .A1(n26119), .B0(n26118), .Y(n26537) );
  CMPR22X1 U30488 ( .A(U0_pipe12[8]), .B(n28804), .CO(n26122), .S(n26066) );
  OAI21XL U30489 ( .A0(n26130), .A1(n26129), .B0(n26128), .Y(n26131) );
  OAI21XL U30490 ( .A0(n26136), .A1(n26135), .B0(n26134), .Y(n26557) );
  CMPR22X1 U30491 ( .A(U0_pipe2[8]), .B(n28788), .CO(n26138), .S(n26043) );
  NAND2XL U30492 ( .A(n26143), .B(n26149), .Y(n26151) );
  OAI21XL U30493 ( .A0(n26146), .A1(n26145), .B0(n26144), .Y(n26147) );
  AOI21XL U30494 ( .A0(n26149), .A1(n26148), .B0(n26147), .Y(n26150) );
  OAI21XL U30495 ( .A0(n26152), .A1(n26151), .B0(n26150), .Y(n26605) );
  CMPR32X1 U30496 ( .A(n26154), .B(n26153), .C(U2_A_r_d[7]), .CO(n26155), .S(
        n26083) );
  NOR2XL U30497 ( .A(n26156), .B(n26155), .Y(n26235) );
  NAND2XL U30498 ( .A(n26156), .B(n26155), .Y(n26237) );
  NAND2XL U30499 ( .A(n26157), .B(n26237), .Y(n26158) );
  OAI21XL U30500 ( .A0(n26319), .A1(n26225), .B0(n26227), .Y(n26164) );
  CMPR22X1 U30501 ( .A(U0_pipe2[9]), .B(n28718), .CO(n26161), .S(n26137) );
  OAI21XL U30502 ( .A0(n26169), .A1(n26168), .B0(n26167), .Y(n26262) );
  OAI21XL U30503 ( .A0(n26264), .A1(n26171), .B0(n26170), .Y(n26208) );
  CMPR22X1 U30504 ( .A(U0_pipe1[9]), .B(U0_pipe0[9]), .CO(n26173), .S(n26104)
         );
  OAI21XL U30505 ( .A0(n26306), .A1(n26215), .B0(n26217), .Y(n26180) );
  CMPR22X1 U30506 ( .A(U0_pipe12[9]), .B(n28722), .CO(n26177), .S(n26121) );
  OAI21XL U30507 ( .A0(n26341), .A1(n26196), .B0(n26198), .Y(n26186) );
  CMPR22X1 U30508 ( .A(U0_pipe8[9]), .B(n28714), .CO(n26183), .S(n26099) );
  OAI21XL U30509 ( .A0(n26354), .A1(n26235), .B0(n26237), .Y(n26194) );
  CMPR32X1 U30510 ( .A(n26189), .B(n26188), .C(U2_A_r_d[8]), .CO(n26190), .S(
        n26156) );
  INVXL U30511 ( .A(n26238), .Y(n26192) );
  NAND2XL U30512 ( .A(n26191), .B(n26190), .Y(n26236) );
  NAND2XL U30513 ( .A(n26192), .B(n26236), .Y(n26193) );
  OAI21XL U30514 ( .A0(n26199), .A1(n26198), .B0(n26197), .Y(n26339) );
  OAI21XL U30515 ( .A0(n26341), .A1(n26201), .B0(n26200), .Y(n26249) );
  CMPR22X1 U30516 ( .A(U0_pipe8[10]), .B(n28771), .CO(n26203), .S(n26182) );
  CMPR22X1 U30517 ( .A(U0_pipe1[10]), .B(U0_pipe0[10]), .CO(n26210), .S(n26172) );
  OAI21XL U30518 ( .A0(n26218), .A1(n26217), .B0(n26216), .Y(n26304) );
  OAI21XL U30519 ( .A0(n26306), .A1(n26220), .B0(n26219), .Y(n26271) );
  CMPR22X1 U30520 ( .A(U0_pipe12[10]), .B(n28803), .CO(n26222), .S(n26176) );
  OAI21XL U30521 ( .A0(n26228), .A1(n26227), .B0(n26226), .Y(n26317) );
  OAI21XL U30522 ( .A0(n26319), .A1(n26230), .B0(n26229), .Y(n26280) );
  CMPR22X1 U30523 ( .A(U0_pipe2[10]), .B(n28787), .CO(n26232), .S(n26160) );
  NOR2XL U30524 ( .A(n26235), .B(n26238), .Y(n26347) );
  OAI21XL U30525 ( .A0(n26238), .A1(n26237), .B0(n26236), .Y(n26352) );
  INVXL U30526 ( .A(n26352), .Y(n26239) );
  OAI21XL U30527 ( .A0(n26354), .A1(n26240), .B0(n26239), .Y(n26289) );
  CMPR32X1 U30528 ( .A(n26242), .B(n26241), .C(U2_A_r_d[9]), .CO(n26243), .S(
        n26191) );
  NOR2XL U30529 ( .A(n26244), .B(n26243), .Y(n26346) );
  INVXL U30530 ( .A(n26346), .Y(n26288) );
  NAND2XL U30531 ( .A(n26244), .B(n26243), .Y(n26349) );
  NAND2XL U30532 ( .A(n26288), .B(n26349), .Y(n26245) );
  CMPR22X1 U30533 ( .A(U0_pipe8[11]), .B(n28770), .CO(n26251), .S(n26202) );
  OAI21XL U30534 ( .A0(n26260), .A1(n26259), .B0(n26258), .Y(n26261) );
  OAI21XL U30535 ( .A0(n26264), .A1(n26486), .B0(n26495), .Y(n26326) );
  CMPR22X1 U30536 ( .A(U0_pipe1[11]), .B(U0_pipe0[11]), .CO(n26266), .S(n26209) );
  CMPR22X1 U30537 ( .A(U0_pipe12[11]), .B(n28802), .CO(n26273), .S(n26221) );
  CMPR22X1 U30538 ( .A(U0_pipe2[11]), .B(n28786), .CO(n26282), .S(n26231) );
  INVXL U30539 ( .A(n26349), .Y(n26287) );
  INVXL U30540 ( .A(n26350), .Y(n26294) );
  NAND2XL U30541 ( .A(n26293), .B(n26292), .Y(n26348) );
  OAI21XL U30542 ( .A0(n26302), .A1(n26301), .B0(n26300), .Y(n26303) );
  OAI21XL U30543 ( .A0(n26306), .A1(n26525), .B0(n26534), .Y(n26364) );
  CMPR22X1 U30544 ( .A(U0_pipe12[12]), .B(n28801), .CO(n26308), .S(n26272) );
  OAI21XL U30545 ( .A0(n26315), .A1(n26314), .B0(n26313), .Y(n26316) );
  OAI21XL U30546 ( .A0(n26319), .A1(n26545), .B0(n26554), .Y(n26393) );
  CMPR22X1 U30547 ( .A(U0_pipe2[12]), .B(n28785), .CO(n26321), .S(n26281) );
  CMPR22X1 U30548 ( .A(U0_pipe1[12]), .B(U0_pipe0[12]), .CO(n26328), .S(n26265) );
  OAI21XL U30549 ( .A0(n26337), .A1(n26336), .B0(n26335), .Y(n26338) );
  OAI21XL U30550 ( .A0(n26341), .A1(n26573), .B0(n26582), .Y(n26373) );
  CMPR22X1 U30551 ( .A(U0_pipe8[12]), .B(n28769), .CO(n26343), .S(n26250) );
  NOR2XL U30552 ( .A(n26346), .B(n26350), .Y(n26353) );
  OAI21XL U30553 ( .A0(n26350), .A1(n26349), .B0(n26348), .Y(n26351) );
  OAI21XL U30554 ( .A0(n26354), .A1(n26593), .B0(n26602), .Y(n26402) );
  INVXL U30555 ( .A(n26402), .Y(n26459) );
  CMPR32X1 U30556 ( .A(n26356), .B(n26355), .C(U2_A_r_d[11]), .CO(n26357), .S(
        n26293) );
  NOR2XL U30557 ( .A(n26358), .B(n26357), .Y(n26453) );
  INVXL U30558 ( .A(n26453), .Y(n26401) );
  NAND2XL U30559 ( .A(n26401), .B(n26455), .Y(n26359) );
  CMPR22X1 U30560 ( .A(U0_pipe12[13]), .B(n28800), .CO(n26366), .S(n26307) );
  CMPR22X1 U30561 ( .A(U0_pipe8[13]), .B(n28768), .CO(n26375), .S(n26342) );
  OAI21XL U30562 ( .A0(n26383), .A1(n26382), .B0(n26381), .Y(n26491) );
  OAI21XL U30563 ( .A0(n26386), .A1(n26385), .B0(n26384), .Y(n26435) );
  CMPR22X1 U30564 ( .A(U0_pipe1[13]), .B(U0_pipe0[13]), .CO(n26388), .S(n26327) );
  CMPR22X1 U30565 ( .A(U0_pipe2[13]), .B(n28784), .CO(n26395), .S(n26320) );
  INVXL U30566 ( .A(n26455), .Y(n26400) );
  CMPR32X1 U30567 ( .A(n26404), .B(n26403), .C(U2_A_r_d[12]), .CO(n26405), .S(
        n26358) );
  INVXL U30568 ( .A(n26456), .Y(n26407) );
  NAND2XL U30569 ( .A(n26406), .B(n26405), .Y(n26454) );
  NAND2XL U30570 ( .A(n26407), .B(n26454), .Y(n26408) );
  OAI21XL U30571 ( .A0(n26414), .A1(n26413), .B0(n26412), .Y(n26530) );
  OAI21XL U30572 ( .A0(n26417), .A1(n26416), .B0(n26415), .Y(n26468) );
  CMPR22X1 U30573 ( .A(U0_pipe12[14]), .B(n28799), .CO(n26419), .S(n26365) );
  OAI21XL U30574 ( .A0(n26425), .A1(n26424), .B0(n26423), .Y(n26578) );
  OAI21XL U30575 ( .A0(n26428), .A1(n26427), .B0(n26426), .Y(n26505) );
  CMPR22X1 U30576 ( .A(U0_pipe8[14]), .B(n28767), .CO(n26430), .S(n26374) );
  CMPR22X1 U30577 ( .A(U0_pipe1[14]), .B(U0_pipe0[14]), .CO(n26437), .S(n26387) );
  OAI21XL U30578 ( .A0(n26445), .A1(n26444), .B0(n26443), .Y(n26550) );
  OAI21XL U30579 ( .A0(n26448), .A1(n26447), .B0(n26446), .Y(n26477) );
  CMPR22X1 U30580 ( .A(U0_pipe2[14]), .B(n28783), .CO(n26450), .S(n26394) );
  NOR2XL U30581 ( .A(n26453), .B(n26456), .Y(n26592) );
  INVXL U30582 ( .A(n26592), .Y(n26458) );
  INVXL U30583 ( .A(n26598), .Y(n26457) );
  OAI21XL U30584 ( .A0(n26459), .A1(n26458), .B0(n26457), .Y(n26514) );
  INVXL U30585 ( .A(n26591), .Y(n26513) );
  NAND2XL U30586 ( .A(n26513), .B(n26595), .Y(n26464) );
  CMPR22X1 U30587 ( .A(U0_pipe12[15]), .B(n28798), .CO(n26470), .S(n26418) );
  CMPR22X1 U30588 ( .A(U0_pipe2[15]), .B(n28782), .CO(n26479), .S(n26449) );
  OAI21XL U30589 ( .A0(n26489), .A1(n26488), .B0(n26487), .Y(n26490) );
  OAI21XL U30590 ( .A0(n26495), .A1(n26494), .B0(n26493), .Y(n26496) );
  CMPR22X1 U30591 ( .A(U0_pipe1[15]), .B(U0_pipe0[15]), .CO(n26500), .S(n26436) );
  CMPR22X1 U30592 ( .A(U0_pipe8[15]), .B(n28766), .CO(n26507), .S(n26429) );
  INVXL U30593 ( .A(n26595), .Y(n26512) );
  AOI21XL U30594 ( .A0(n26514), .A1(n26513), .B0(n26512), .Y(n26521) );
  NOR2X2 U30595 ( .A(n26518), .B(n26517), .Y(n26596) );
  INVXL U30596 ( .A(n26596), .Y(n26519) );
  NAND2XL U30597 ( .A(n26518), .B(n26517), .Y(n26594) );
  XOR2X1 U30598 ( .A(n26521), .B(n26520), .Y(n26522) );
  OAI21XL U30599 ( .A0(n26528), .A1(n26527), .B0(n26526), .Y(n26529) );
  OAI21XL U30600 ( .A0(n26534), .A1(n26533), .B0(n26532), .Y(n26535) );
  OAI21XL U30601 ( .A0(n26548), .A1(n26547), .B0(n26546), .Y(n26549) );
  OAI21XL U30602 ( .A0(n26554), .A1(n26553), .B0(n26552), .Y(n26555) );
  CMPR22X1 U30603 ( .A(U0_pipe1[16]), .B(U0_pipe0[16]), .CO(n26566), .S(n26499) );
  OAI21XL U30604 ( .A0(n26576), .A1(n26575), .B0(n26574), .Y(n26577) );
  OAI21XL U30605 ( .A0(n26582), .A1(n26581), .B0(n26580), .Y(n26583) );
  NOR2XL U30606 ( .A(n26591), .B(n26596), .Y(n26599) );
  NAND2XL U30607 ( .A(n26592), .B(n26599), .Y(n26601) );
  NOR2XL U30608 ( .A(n26593), .B(n26601), .Y(n26604) );
  OAI21XL U30609 ( .A0(n26596), .A1(n26595), .B0(n26594), .Y(n26597) );
  AOI21X1 U30610 ( .A0(n26599), .A1(n26598), .B0(n26597), .Y(n26600) );
  OAI21X1 U30611 ( .A0(n26602), .A1(n26601), .B0(n26600), .Y(n26603) );
  AOI21X1 U30612 ( .A0(n26605), .A1(n26604), .B0(n26603), .Y(n26865) );
  INVXL U30613 ( .A(n26865), .Y(n26818) );
  CMPR32X1 U30614 ( .A(n26607), .B(n26606), .C(U2_A_r_d[15]), .CO(n26608), .S(
        n26518) );
  NOR2XL U30615 ( .A(n26609), .B(n26608), .Y(n26698) );
  INVXL U30616 ( .A(n26698), .Y(n26644) );
  NAND2XL U30617 ( .A(n26644), .B(n26700), .Y(n26610) );
  OAI21XL U30618 ( .A0(n26629), .A1(n26628), .B0(n26627), .Y(n26678) );
  INVXL U30619 ( .A(n26700), .Y(n26643) );
  AOI21XL U30620 ( .A0(n26818), .A1(n26644), .B0(n26643), .Y(n26651) );
  CMPR32X1 U30621 ( .A(n26646), .B(n26645), .C(U2_A_r_d[16]), .CO(n26647), .S(
        n26609) );
  INVXL U30622 ( .A(n26701), .Y(n26649) );
  NAND2XL U30623 ( .A(n26648), .B(n26647), .Y(n26699) );
  NAND2XL U30624 ( .A(n26649), .B(n26699), .Y(n26650) );
  CMPR22X1 U30625 ( .A(U0_pipe12[18]), .B(n28795), .CO(n26659), .S(n26614) );
  CMPR22X1 U30626 ( .A(U0_pipe8[18]), .B(n28763), .CO(n26670), .S(n26621) );
  CMPR22X1 U30627 ( .A(U0_pipe1[18]), .B(U0_pipe0[18]), .CO(n26682), .S(n26631) );
  CMPR22X1 U30628 ( .A(U0_pipe2[18]), .B(n28779), .CO(n26693), .S(n26638) );
  AOI21XL U30629 ( .A0(n26818), .A1(n26753), .B0(n26756), .Y(n26707) );
  ADDFHX1 U30630 ( .A(n26703), .B(n26702), .CI(U2_A_r_d[17]), .CO(n26704), .S(
        n26648) );
  OR2X2 U30631 ( .A(n26705), .B(n26704), .Y(n26755) );
  NAND2XL U30632 ( .A(n26705), .B(n26704), .Y(n26754) );
  NAND2XL U30633 ( .A(n26755), .B(n26754), .Y(n26706) );
  OAI21XL U30634 ( .A0(n26712), .A1(n26711), .B0(n26710), .Y(n26770) );
  OAI21XL U30635 ( .A0(n26723), .A1(n26722), .B0(n26721), .Y(n26806) );
  OAI21XL U30636 ( .A0(n26734), .A1(n26733), .B0(n26732), .Y(n26794) );
  OAI21XL U30637 ( .A0(n26745), .A1(n26744), .B0(n26743), .Y(n26782) );
  NAND2X1 U30638 ( .A(n26753), .B(n26755), .Y(n26815) );
  INVXL U30639 ( .A(n26815), .Y(n26758) );
  AOI21XL U30640 ( .A0(n26818), .A1(n26758), .B0(n26757), .Y(n26765) );
  NAND2XL U30641 ( .A(n26762), .B(n26761), .Y(n26816) );
  OAI21XL U30642 ( .A0(n26773), .A1(n26772), .B0(n26771), .Y(n26829) );
  OAI21XL U30643 ( .A0(n26785), .A1(n26784), .B0(n26783), .Y(n26837) );
  OAI21XL U30644 ( .A0(n26797), .A1(n26796), .B0(n26795), .Y(n26845) );
  NAND2XL U30645 ( .A(n26798), .B(n26843), .Y(n26801) );
  OAI21XL U30646 ( .A0(n26809), .A1(n26808), .B0(n26807), .Y(n26853) );
  NOR2X1 U30647 ( .A(n26815), .B(n26817), .Y(n26859) );
  AOI21XL U30648 ( .A0(n26818), .A1(n26859), .B0(n26862), .Y(n26825) );
  NAND2XL U30649 ( .A(n26823), .B(n26822), .Y(n26860) );
  CMPR22X1 U30650 ( .A(U0_pipe12[21]), .B(n28792), .CO(n26831), .S(n26775) );
  CMPR22X1 U30651 ( .A(U0_pipe8[21]), .B(n28760), .CO(n26839), .S(n26787) );
  CMPR22X1 U30652 ( .A(U0_pipe1[21]), .B(U0_pipe0[21]), .CO(n26847), .S(n26799) );
  CMPR22X1 U30653 ( .A(U0_pipe2[21]), .B(n28776), .CO(n26855), .S(n26811) );
  NAND2X1 U30654 ( .A(n26859), .B(n26821), .Y(n26864) );
  INVXL U30655 ( .A(n26860), .Y(n26861) );
  AOI21X1 U30656 ( .A0(n26862), .A1(n26821), .B0(n26861), .Y(n26863) );
  OAI21X1 U30657 ( .A0(n26865), .A1(n26864), .B0(n26863), .Y(n26907) );
  CMPR32X1 U30658 ( .A(n26867), .B(n26866), .C(U2_A_r_d[20]), .CO(n26868), .S(
        n26823) );
  OR2X2 U30659 ( .A(n26869), .B(n26868), .Y(n26906) );
  NAND2X1 U30660 ( .A(n26869), .B(n26868), .Y(n26904) );
  XNOR2X1 U30661 ( .A(n26907), .B(n26870), .Y(n26871) );
  OAI21XL U30662 ( .A0(n26874), .A1(n26873), .B0(n26872), .Y(n26916) );
  OAI21XL U30663 ( .A0(n26882), .A1(n26881), .B0(n26880), .Y(n26924) );
  OAI21XL U30664 ( .A0(n26890), .A1(n26889), .B0(n26888), .Y(n26932) );
  OAI21XL U30665 ( .A0(n26898), .A1(n26897), .B0(n26896), .Y(n26940) );
  CMPR32X1 U30666 ( .A(n26909), .B(n26908), .C(U2_A_r_d[21]), .CO(n26910), .S(
        n26869) );
  NOR2X1 U30667 ( .A(n26911), .B(n26910), .Y(n26947) );
  CMPR22X1 U30668 ( .A(U0_pipe12[23]), .B(n28933), .CO(n26918), .S(n26876) );
  CMPR22X1 U30669 ( .A(U0_pipe8[23]), .B(n28925), .CO(n26926), .S(n26884) );
  CMPR22X1 U30670 ( .A(U0_pipe1[23]), .B(U0_pipe0[23]), .CO(n26934), .S(n26892) );
  CMPR22X1 U30671 ( .A(U0_pipe2[23]), .B(n28929), .CO(n26942), .S(n26900) );
  CMPR32X1 U30672 ( .A(n26949), .B(n26948), .C(U2_A_r_d[22]), .CO(n26950), .S(
        n26911) );
  OR2X2 U30673 ( .A(n26951), .B(n26950), .Y(n26988) );
  OAI21XL U30674 ( .A0(n26956), .A1(n26955), .B0(n26954), .Y(n26999) );
  OAI21XL U30675 ( .A0(n26964), .A1(n26963), .B0(n26962), .Y(n27007) );
  OAI21XL U30676 ( .A0(n26972), .A1(n26971), .B0(n26970), .Y(n27015) );
  OAI21XL U30677 ( .A0(n26980), .A1(n26979), .B0(n26978), .Y(n27023) );
  CMPR32X1 U30678 ( .A(n26991), .B(n26990), .C(U2_A_r_d[23]), .CO(n26992), .S(
        n26951) );
  CMPR22X1 U30679 ( .A(U0_pipe12[25]), .B(n28931), .CO(n27001), .S(n26958) );
  CMPR22X1 U30680 ( .A(U0_pipe2[25]), .B(n28927), .CO(n27009), .S(n26966) );
  CMPR22X1 U30681 ( .A(U0_pipe1[25]), .B(U0_pipe0[25]), .CO(n27017), .S(n26974) );
  CMPR22X1 U30682 ( .A(U0_pipe8[25]), .B(n28923), .CO(n27025), .S(n26982) );
  CMPR32X1 U30683 ( .A(n27033), .B(n27032), .C(U2_A_r_d[24]), .CO(n27034), .S(
        n26993) );
  MXI2X1 U30684 ( .A(U2_pipe0[25]), .B(n27041), .S0(n27040), .Y(n4093) );
  CMPR22X1 U30685 ( .A(U0_pipe12[26]), .B(n29001), .CO(n27047), .S(n27000) );
  OAI21XL U30686 ( .A0(n27045), .A1(n27044), .B0(n27043), .Y(n27046) );
  CMPR32X1 U30687 ( .A(n27048), .B(n27047), .C(n27046), .S(n27049) );
  CMPR22X1 U30688 ( .A(U0_pipe2[26]), .B(n29000), .CO(n27054), .S(n27008) );
  OAI21XL U30689 ( .A0(n27052), .A1(n27051), .B0(n27050), .Y(n27053) );
  CMPR32X1 U30690 ( .A(n27055), .B(n27054), .C(n27053), .S(n27056) );
  CMPR22X1 U30691 ( .A(U0_pipe1[26]), .B(U0_pipe0[26]), .CO(n27061), .S(n27016) );
  OAI21XL U30692 ( .A0(n27059), .A1(n27058), .B0(n27057), .Y(n27060) );
  CMPR32X1 U30693 ( .A(n27062), .B(n27061), .C(n27060), .S(n27063) );
  CMPR22X1 U30694 ( .A(U0_pipe8[26]), .B(n28999), .CO(n27068), .S(n27024) );
  OAI21XL U30695 ( .A0(n27066), .A1(n27065), .B0(n27064), .Y(n27067) );
  CMPR32X1 U30696 ( .A(n27069), .B(n27068), .C(n27067), .S(n27070) );
  AOI21XL U30697 ( .A0(n5921), .A1(Q0_addr[0]), .B0(n27081), .Y(n27072) );
  AOI21XL U30698 ( .A0(n5921), .A1(Q0_addr[1]), .B0(n27073), .Y(n27075) );
  AOI21XL U30699 ( .A0(n5921), .A1(Q0_addr[2]), .B0(n27084), .Y(n27077) );
  AOI21XL U30700 ( .A0(n5798), .A1(Q0_addr[0]), .B0(n27081), .Y(n27083) );
  AOI22XL U30701 ( .A0(Q3_addr[0]), .A1(n27497), .B0(Q2_addr[0]), .B1(n27496), 
        .Y(n27082) );
  AOI21XL U30702 ( .A0(n5918), .A1(Q0_addr[2]), .B0(n27084), .Y(n27086) );
  AOI22XL U30703 ( .A0(Q3_addr[2]), .A1(n27497), .B0(Q2_addr[2]), .B1(n27496), 
        .Y(n27085) );
  AOI22X1 U30704 ( .A0(n7123), .A1(CQ1[0]), .B0(Q6[0]), .B1(n27211), .Y(n27503) );
  AOI22X1 U30705 ( .A0(n7123), .A1(CQ1[0]), .B0(Q7[0]), .B1(n28922), .Y(n27499) );
  OAI21XL U30706 ( .A0(n5823), .A1(n27503), .B0(n27090), .Y(A7_d[0]) );
  AOI22X1 U30707 ( .A0(n7123), .A1(CQ1[1]), .B0(Q6[1]), .B1(n28922), .Y(n27504) );
  NOR2BX1 U30708 ( .AN(buffer[1]), .B(n27122), .Y(n28291) );
  AOI22X1 U30709 ( .A0(n7123), .A1(CQ1[1]), .B0(Q7[1]), .B1(n28922), .Y(n27505) );
  AOI22X1 U30710 ( .A0(n7123), .A1(CQ1[1]), .B0(Q5[1]), .B1(n28922), .Y(n27509) );
  OAI21XL U30711 ( .A0(n5823), .A1(n27504), .B0(n27093), .Y(A7_d[1]) );
  AOI22X1 U30712 ( .A0(n7123), .A1(CQ1[2]), .B0(Q6[2]), .B1(n28922), .Y(n27510) );
  NOR2BX1 U30713 ( .AN(buffer[2]), .B(n27122), .Y(n28299) );
  AOI22X1 U30714 ( .A0(n7123), .A1(CQ1[2]), .B0(Q7[2]), .B1(n28922), .Y(n27511) );
  AOI22X1 U30715 ( .A0(n7123), .A1(CQ1[2]), .B0(Q5[2]), .B1(n28922), .Y(n27515) );
  OAI21XL U30716 ( .A0(n5823), .A1(n27510), .B0(n27096), .Y(A7_d[2]) );
  AOI22X1 U30717 ( .A0(n7123), .A1(CQ1[3]), .B0(Q7[3]), .B1(n28922), .Y(n27517) );
  AOI22X1 U30718 ( .A0(n7123), .A1(CQ1[3]), .B0(Q5[3]), .B1(n28922), .Y(n27521) );
  OAI21XL U30719 ( .A0(n5823), .A1(n27516), .B0(n27099), .Y(A7_d[3]) );
  AOI22X1 U30720 ( .A0(n7123), .A1(CQ1[4]), .B0(Q5[4]), .B1(n28922), .Y(n27527) );
  NOR2BX1 U30721 ( .AN(buffer[4]), .B(n27122), .Y(n28313) );
  AOI22X1 U30722 ( .A0(n7123), .A1(CQ1[4]), .B0(Q7[4]), .B1(n28922), .Y(n27523) );
  OAI21XL U30723 ( .A0(n7140), .A1(n27527), .B0(n27102), .Y(A7_d[4]) );
  CLKINVX3 U30724 ( .A(n27205), .Y(n27264) );
  AOI22X1 U30725 ( .A0(n7123), .A1(CQ1[5]), .B0(Q6[5]), .B1(n28922), .Y(n27533) );
  NOR2BX1 U30726 ( .AN(buffer[5]), .B(n27122), .Y(n28320) );
  AOI22X1 U30727 ( .A0(n5840), .A1(CQ1[5]), .B0(Q7[5]), .B1(n28922), .Y(n27529) );
  AOI22X1 U30728 ( .A0(n5840), .A1(CQ1[5]), .B0(Q5[5]), .B1(n28922), .Y(n27528) );
  OAI21XL U30729 ( .A0(n27264), .A1(n27533), .B0(n27105), .Y(A7_d[5]) );
  AOI22X1 U30730 ( .A0(n5927), .A1(CQ1[6]), .B0(Q6[6]), .B1(n28922), .Y(n27539) );
  AOI22X1 U30731 ( .A0(n5927), .A1(CQ1[6]), .B0(Q7[6]), .B1(n27211), .Y(n27535) );
  OAI21XL U30732 ( .A0(n5823), .A1(n27539), .B0(n27108), .Y(A7_d[6]) );
  AOI22X1 U30733 ( .A0(n5927), .A1(CQ1[7]), .B0(Q5[7]), .B1(n28922), .Y(n27545) );
  AOI22X1 U30734 ( .A0(n5927), .A1(CQ1[7]), .B0(Q7[7]), .B1(n27211), .Y(n27541) );
  AOI22X1 U30735 ( .A0(n5927), .A1(CQ1[7]), .B0(Q6[7]), .B1(n27211), .Y(n27540) );
  OAI21XL U30736 ( .A0(n7140), .A1(n27545), .B0(n27111), .Y(A7_d[7]) );
  AOI22X1 U30737 ( .A0(n5927), .A1(CQ1[8]), .B0(Q6[8]), .B1(n28922), .Y(n27551) );
  AOI22X1 U30738 ( .A0(n5927), .A1(CQ1[8]), .B0(Q7[8]), .B1(n27211), .Y(n27547) );
  OAI21XL U30739 ( .A0(n27264), .A1(n27551), .B0(n27114), .Y(A7_d[8]) );
  AOI22X1 U30740 ( .A0(n5927), .A1(CQ1[9]), .B0(Q6[9]), .B1(n27213), .Y(n27557) );
  AOI22X1 U30741 ( .A0(n5927), .A1(CQ1[9]), .B0(Q7[9]), .B1(n27213), .Y(n27553) );
  OAI21XL U30742 ( .A0(n5823), .A1(n27557), .B0(n27117), .Y(A7_d[9]) );
  AOI22X1 U30743 ( .A0(n5927), .A1(CQ1[10]), .B0(Q5[10]), .B1(n27211), .Y(
        n27558) );
  AOI22X1 U30744 ( .A0(n5927), .A1(CQ1[10]), .B0(Q7[10]), .B1(n28922), .Y(
        n27559) );
  OAI21XL U30745 ( .A0(n7140), .A1(n27558), .B0(n27120), .Y(A7_d[10]) );
  OAI21XL U30746 ( .A0(Q5[11]), .A1(n5927), .B0(n27123), .Y(n27570) );
  OAI21X1 U30747 ( .A0(n28955), .A1(n27976), .B0(n27121), .Y(n27568) );
  OAI21XL U30748 ( .A0(n7140), .A1(n7098), .B0(n27125), .Y(A7_d[11]) );
  OAI21XL U30749 ( .A0(Q5[12]), .A1(n5927), .B0(n27127), .Y(n27576) );
  NOR2BX1 U30750 ( .AN(buffer[12]), .B(n5922), .Y(n28371) );
  OAI21XL U30751 ( .A0(n7140), .A1(n7106), .B0(n27129), .Y(A7_d[12]) );
  NOR2BX1 U30752 ( .AN(buffer[13]), .B(n5922), .Y(n28378) );
  OAI21XL U30753 ( .A0(n27264), .A1(n27577), .B0(n27133), .Y(A7_d[13]) );
  NOR2BX1 U30754 ( .AN(buffer[14]), .B(n5922), .Y(n28385) );
  OAI21XL U30755 ( .A0(Q6[14]), .A1(n5840), .B0(n27135), .Y(n27588) );
  OAI21XL U30756 ( .A0(n7140), .A1(n27583), .B0(n27137), .Y(A7_d[14]) );
  OAI21XL U30757 ( .A0(Q5[15]), .A1(n5840), .B0(n27139), .Y(n27594) );
  OAI21X1 U30758 ( .A0(n28959), .A1(n27976), .B0(n27138), .Y(n27592) );
  OAI21XL U30759 ( .A0(n7140), .A1(n7100), .B0(n27141), .Y(A7_d[15]) );
  OAI21X1 U30760 ( .A0(n28960), .A1(n27976), .B0(n27142), .Y(n27598) );
  OAI21XL U30761 ( .A0(Q5[16]), .A1(n5840), .B0(n27143), .Y(n27600) );
  OAI21XL U30762 ( .A0(n27264), .A1(n27595), .B0(n27145), .Y(A7_d[16]) );
  OAI21X1 U30763 ( .A0(n28961), .A1(OP2_done0), .B0(n27146), .Y(n27604) );
  OAI21XL U30764 ( .A0(Q6[17]), .A1(n5840), .B0(n27147), .Y(n27606) );
  OAI21XL U30765 ( .A0(n7140), .A1(n27601), .B0(n27149), .Y(A7_d[17]) );
  OAI21X1 U30766 ( .A0(n28962), .A1(n27976), .B0(n27150), .Y(n27610) );
  OAI21X1 U30767 ( .A0(Q7[18]), .A1(OP_done1), .B0(n27151), .Y(n27608) );
  OAI21XL U30768 ( .A0(Q5[18]), .A1(OP_done1), .B0(n27151), .Y(n27612) );
  OAI21XL U30769 ( .A0(n27264), .A1(n27607), .B0(n27153), .Y(A7_d[18]) );
  OAI21XL U30770 ( .A0(Q6[19]), .A1(OP_done1), .B0(n27155), .Y(n27618) );
  OAI21X1 U30771 ( .A0(n28963), .A1(n27976), .B0(n27154), .Y(n27616) );
  OAI21X1 U30772 ( .A0(Q7[19]), .A1(OP_done1), .B0(n27155), .Y(n27614) );
  OAI21XL U30773 ( .A0(n5823), .A1(n7090), .B0(n27157), .Y(A7_d[19]) );
  OAI21XL U30774 ( .A0(Q5[20]), .A1(OP_done1), .B0(n27159), .Y(n27624) );
  OAI21X1 U30775 ( .A0(n28964), .A1(OP2_done0), .B0(n27158), .Y(n27622) );
  OAI21X1 U30776 ( .A0(Q7[20]), .A1(OP_done1), .B0(n27159), .Y(n27620) );
  OAI21XL U30777 ( .A0(n7140), .A1(n7108), .B0(n27161), .Y(A7_d[20]) );
  OAI21XL U30778 ( .A0(Q6[21]), .A1(n5927), .B0(n27164), .Y(n27630) );
  OAI21X1 U30779 ( .A0(n28965), .A1(n27976), .B0(n27163), .Y(n27628) );
  OAI21XL U30780 ( .A0(Q5[21]), .A1(n5927), .B0(n27164), .Y(n27625) );
  OAI21XL U30781 ( .A0(n27264), .A1(n27630), .B0(n27166), .Y(A7_d[21]) );
  OAI21X1 U30782 ( .A0(n28966), .A1(n27976), .B0(n27167), .Y(n27635) );
  OAI21XL U30783 ( .A0(Q5[22]), .A1(OP_done1), .B0(n27168), .Y(n27632) );
  OAI21XL U30784 ( .A0(n27264), .A1(n27637), .B0(n27170), .Y(A7_d[22]) );
  OAI21X1 U30785 ( .A0(n28967), .A1(n27976), .B0(n27171), .Y(n27641) );
  OAI21X1 U30786 ( .A0(Q7[23]), .A1(OP_done1), .B0(n27172), .Y(n27639) );
  OAI21XL U30787 ( .A0(n27264), .A1(n27638), .B0(n27174), .Y(A7_d[23]) );
  OAI21XL U30788 ( .A0(Q6[24]), .A1(n5927), .B0(n27176), .Y(n27649) );
  OAI21X1 U30789 ( .A0(n28968), .A1(n27976), .B0(n27175), .Y(n27647) );
  OAI21XL U30790 ( .A0(n27264), .A1(n7092), .B0(n27178), .Y(A7_d[24]) );
  OAI21XL U30791 ( .A0(Q5[25]), .A1(n5840), .B0(n27180), .Y(n27655) );
  OAI21X1 U30792 ( .A0(n28969), .A1(n27976), .B0(n27179), .Y(n27653) );
  OAI21XL U30793 ( .A0(n7140), .A1(n7094), .B0(n27182), .Y(A7_d[25]) );
  AOI22X1 U30794 ( .A0(n5840), .A1(CQ1[26]), .B0(Q6[28]), .B1(n28922), .Y(
        n27661) );
  NOR2BX1 U30795 ( .AN(buffer[16]), .B(n5922), .Y(n28459) );
  AOI22X1 U30796 ( .A0(n5840), .A1(CQ1[26]), .B0(Q7[28]), .B1(n27211), .Y(
        n27657) );
  OAI21XL U30797 ( .A0(n27264), .A1(n27661), .B0(n27185), .Y(A7_d[26]) );
  NOR2BX1 U30798 ( .AN(buffer[17]), .B(n5922), .Y(n28466) );
  AOI22X1 U30799 ( .A0(n5840), .A1(CQ1[27]), .B0(Q7[29]), .B1(n28922), .Y(
        n27663) );
  AOI22X1 U30800 ( .A0(n5840), .A1(CQ1[27]), .B0(Q5[29]), .B1(n28922), .Y(
        n27667) );
  OAI21XL U30801 ( .A0(n5823), .A1(n27662), .B0(n27188), .Y(A7_d[27]) );
  AOI22X1 U30802 ( .A0(OP_done1), .A1(CQ1[28]), .B0(Q6[30]), .B1(n28922), .Y(
        n27668) );
  AOI22X1 U30803 ( .A0(n5927), .A1(CQ1[28]), .B0(Q7[30]), .B1(n28922), .Y(
        n27669) );
  AOI22X1 U30804 ( .A0(n5927), .A1(CQ1[28]), .B0(Q5[30]), .B1(n28922), .Y(
        n27673) );
  OAI21XL U30805 ( .A0(n27264), .A1(n27668), .B0(n27191), .Y(A7_d[28]) );
  AOI22X1 U30806 ( .A0(OP_done1), .A1(CQ1[29]), .B0(Q5[31]), .B1(n28922), .Y(
        n27674) );
  AOI22X1 U30807 ( .A0(n5927), .A1(CQ1[29]), .B0(Q7[31]), .B1(n28922), .Y(
        n27675) );
  AOI22X1 U30808 ( .A0(OP_done1), .A1(CQ1[29]), .B0(Q6[31]), .B1(n28922), .Y(
        n27679) );
  OAI21XL U30809 ( .A0(n7140), .A1(n27674), .B0(n27194), .Y(A7_d[29]) );
  AOI22X1 U30810 ( .A0(OP_done1), .A1(CQ1[30]), .B0(Q6[32]), .B1(n28922), .Y(
        n27685) );
  AOI22X1 U30811 ( .A0(n5927), .A1(CQ1[30]), .B0(Q7[32]), .B1(n27213), .Y(
        n27681) );
  OAI21XL U30812 ( .A0(n5823), .A1(n27685), .B0(n27197), .Y(A7_d[30]) );
  AOI22X1 U30813 ( .A0(n5927), .A1(CQ1[31]), .B0(Q6[33]), .B1(n27213), .Y(
        n27687) );
  AOI22X1 U30814 ( .A0(n5927), .A1(CQ1[31]), .B0(Q7[33]), .B1(n27213), .Y(
        n27688) );
  AOI22X1 U30815 ( .A0(n5927), .A1(CQ1[31]), .B0(Q5[33]), .B1(n27211), .Y(
        n27692) );
  OAI21XL U30816 ( .A0(n27264), .A1(n27687), .B0(n27200), .Y(A7_d[31]) );
  AOI22X1 U30817 ( .A0(n5840), .A1(CQ1[32]), .B0(Q5[34]), .B1(n28922), .Y(
        n27698) );
  NOR2BX1 U30818 ( .AN(buffer[22]), .B(n5922), .Y(n28501) );
  AOI22X1 U30819 ( .A0(n5840), .A1(CQ1[32]), .B0(Q7[34]), .B1(n27211), .Y(
        n27694) );
  OAI21XL U30820 ( .A0(n7140), .A1(n27698), .B0(n27203), .Y(A7_d[32]) );
  AOI22X1 U30821 ( .A0(n5840), .A1(CQ1[33]), .B0(Q5[35]), .B1(n28922), .Y(
        n27699) );
  NOR2BX1 U30822 ( .AN(buffer[23]), .B(n5922), .Y(n28508) );
  AOI22X1 U30823 ( .A0(n5840), .A1(CQ1[33]), .B0(Q7[35]), .B1(n28922), .Y(
        n27700) );
  OAI21XL U30824 ( .A0(n7140), .A1(n27699), .B0(n27207), .Y(A7_d[33]) );
  AOI22X1 U30825 ( .A0(n5927), .A1(CQ1[34]), .B0(Q6[36]), .B1(n27211), .Y(
        n27705) );
  AOI22X1 U30826 ( .A0(n5927), .A1(CQ1[34]), .B0(Q7[36]), .B1(n27213), .Y(
        n27706) );
  AOI22X1 U30827 ( .A0(n5927), .A1(CQ1[34]), .B0(Q5[36]), .B1(n27213), .Y(
        n27710) );
  OAI21XL U30828 ( .A0(n5823), .A1(n27705), .B0(n27210), .Y(A7_d[34]) );
  AOI22X1 U30829 ( .A0(n5840), .A1(CQ1[35]), .B0(Q6[37]), .B1(n27211), .Y(
        n27711) );
  NOR2BX1 U30830 ( .AN(buffer[25]), .B(n5922), .Y(n28522) );
  AOI22X1 U30831 ( .A0(n5840), .A1(CQ1[35]), .B0(Q7[37]), .B1(n27211), .Y(
        n27712) );
  AOI22X1 U30832 ( .A0(n5840), .A1(CQ1[35]), .B0(Q5[37]), .B1(n27211), .Y(
        n27716) );
  OAI21XL U30833 ( .A0(n27264), .A1(n27711), .B0(n27215), .Y(A7_d[35]) );
  AOI22X1 U30834 ( .A0(n7123), .A1(CQ1[36]), .B0(Q6[38]), .B1(n27211), .Y(
        n27722) );
  AOI22X1 U30835 ( .A0(n5840), .A1(CQ1[36]), .B0(Q7[38]), .B1(n27213), .Y(
        n27718) );
  OAI21XL U30836 ( .A0(n5823), .A1(n27722), .B0(n27218), .Y(A7_d[36]) );
  OAI21X1 U30837 ( .A0(n28970), .A1(n27976), .B0(n27219), .Y(n27726) );
  OAI21XL U30838 ( .A0(Q5[39]), .A1(n5840), .B0(n27220), .Y(n27728) );
  OAI21XL U30839 ( .A0(n27264), .A1(n27723), .B0(n27222), .Y(A7_d[37]) );
  OAI21X1 U30840 ( .A0(n28971), .A1(n27976), .B0(n27223), .Y(n27732) );
  OAI21XL U30841 ( .A0(Q5[40]), .A1(n5840), .B0(n27224), .Y(n27734) );
  OAI21XL U30842 ( .A0(n5823), .A1(n27729), .B0(n27226), .Y(A7_d[38]) );
  OAI21XL U30843 ( .A0(Q6[41]), .A1(n5840), .B0(n27228), .Y(n27740) );
  OAI21X1 U30844 ( .A0(n28972), .A1(n27976), .B0(n27227), .Y(n27738) );
  OAI21XL U30845 ( .A0(n27264), .A1(n7116), .B0(n27230), .Y(A7_d[39]) );
  OAI21X1 U30846 ( .A0(n28973), .A1(n27976), .B0(n27231), .Y(n27744) );
  OAI21XL U30847 ( .A0(n28054), .A1(n27741), .B0(n27234), .Y(A7_d[40]) );
  OAI21X1 U30848 ( .A0(n28974), .A1(n27976), .B0(n27235), .Y(n27750) );
  OAI21X1 U30849 ( .A0(Q7[43]), .A1(n7123), .B0(n27237), .Y(n27748) );
  OAI21XL U30850 ( .A0(n7140), .A1(n27752), .B0(n27239), .Y(A7_d[41]) );
  OAI21X1 U30851 ( .A0(n28975), .A1(n27976), .B0(n27240), .Y(n27756) );
  OAI21X1 U30852 ( .A0(Q7[44]), .A1(n7123), .B0(n27241), .Y(n27754) );
  OAI21XL U30853 ( .A0(n28054), .A1(n27753), .B0(n27243), .Y(A7_d[42]) );
  OAI21X1 U30854 ( .A0(n28976), .A1(n27976), .B0(n27244), .Y(n27762) );
  OAI21X1 U30855 ( .A0(Q7[45]), .A1(n7123), .B0(n27245), .Y(n27760) );
  OAI21XL U30856 ( .A0(n7140), .A1(n27764), .B0(n27247), .Y(A7_d[43]) );
  OAI21XL U30857 ( .A0(Q5[46]), .A1(n5927), .B0(n27249), .Y(n27770) );
  OAI21X1 U30858 ( .A0(n28977), .A1(n27976), .B0(n27248), .Y(n27768) );
  OAI21X1 U30859 ( .A0(Q7[46]), .A1(OP_done1), .B0(n27249), .Y(n27766) );
  OAI21XL U30860 ( .A0(n7140), .A1(n7110), .B0(n27251), .Y(A7_d[44]) );
  OAI21XL U30861 ( .A0(Q5[47]), .A1(n5927), .B0(n27253), .Y(n27771) );
  OAI21X1 U30862 ( .A0(n28978), .A1(n27976), .B0(n27252), .Y(n27775) );
  OAI21XL U30863 ( .A0(n7140), .A1(n7086), .B0(n27255), .Y(A7_d[45]) );
  OAI21X1 U30864 ( .A0(n28979), .A1(n27976), .B0(n27256), .Y(n27781) );
  OAI21XL U30865 ( .A0(Q5[48]), .A1(n5927), .B0(n27257), .Y(n27783) );
  OAI21XL U30866 ( .A0(n28054), .A1(n27778), .B0(n27259), .Y(A7_d[46]) );
  OAI21X1 U30867 ( .A0(n28980), .A1(n27976), .B0(n27260), .Y(n27787) );
  OAI21XL U30868 ( .A0(n27264), .A1(n27789), .B0(n27263), .Y(A7_d[47]) );
  OAI21X1 U30869 ( .A0(Q7[50]), .A1(OP_done1), .B0(n27266), .Y(n27791) );
  OAI21XL U30870 ( .A0(n28054), .A1(n27790), .B0(n27268), .Y(A7_d[48]) );
  OAI21X1 U30871 ( .A0(n28982), .A1(n27976), .B0(n27269), .Y(n27799) );
  OAI21X1 U30872 ( .A0(Q7[51]), .A1(OP_done1), .B0(n27270), .Y(n27797) );
  OAI21XL U30873 ( .A0(n7140), .A1(n27796), .B0(n27272), .Y(A7_d[49]) );
  OAI21X1 U30874 ( .A0(n28983), .A1(n27976), .B0(n27273), .Y(n27805) );
  OAI21X1 U30875 ( .A0(Q7[52]), .A1(OP_done1), .B0(n27274), .Y(n27803) );
  OAI21XL U30876 ( .A0(n7140), .A1(n27802), .B0(n27276), .Y(A7_d[50]) );
  OAI21X1 U30877 ( .A0(n28984), .A1(n27976), .B0(n27277), .Y(n27811) );
  OAI21X1 U30878 ( .A0(Q7[53]), .A1(OP_done1), .B0(n27278), .Y(n27809) );
  OAI21XL U30879 ( .A0(n7140), .A1(n27808), .B0(n27280), .Y(A7_d[51]) );
  OAI21XL U30880 ( .A0(n28158), .A1(n27503), .B0(n27283), .Y(A6_d[0]) );
  OAI21XL U30881 ( .A0(n28138), .A1(n27504), .B0(n27285), .Y(A6_d[1]) );
  OAI21XL U30882 ( .A0(n28118), .A1(n27510), .B0(n27287), .Y(A6_d[2]) );
  CLKINVX3 U30883 ( .A(n5904), .Y(n28093) );
  OAI21XL U30884 ( .A0(n28068), .A1(n27521), .B0(n27289), .Y(A6_d[3]) );
  OAI21XL U30885 ( .A0(n28118), .A1(n27522), .B0(n27291), .Y(A6_d[4]) );
  OAI21XL U30886 ( .A0(n28068), .A1(n27528), .B0(n27293), .Y(A6_d[5]) );
  OAI21XL U30887 ( .A0(n28138), .A1(n27539), .B0(n27295), .Y(A6_d[6]) );
  OAI21XL U30888 ( .A0(n28138), .A1(n27540), .B0(n27297), .Y(A6_d[7]) );
  CLKINVX3 U30889 ( .A(n5904), .Y(n28138) );
  OAI21XL U30890 ( .A0(n28068), .A1(n27546), .B0(n27300), .Y(A6_d[8]) );
  OAI21XL U30891 ( .A0(n28165), .A1(n27557), .B0(n27302), .Y(A6_d[9]) );
  OAI21XL U30892 ( .A0(n28068), .A1(n27558), .B0(n27304), .Y(A6_d[10]) );
  CLKINVX3 U30893 ( .A(n5904), .Y(n28158) );
  OAI21XL U30894 ( .A0(n28158), .A1(n27565), .B0(n27306), .Y(A6_d[11]) );
  OAI21XL U30895 ( .A0(n28068), .A1(n7106), .B0(n27308), .Y(A6_d[12]) );
  OAI21XL U30896 ( .A0(n28068), .A1(n27582), .B0(n27310), .Y(A6_d[13]) );
  OAI21XL U30897 ( .A0(n28158), .A1(n7112), .B0(n27312), .Y(A6_d[14]) );
  OAI21XL U30898 ( .A0(n28165), .A1(n27589), .B0(n27314), .Y(A6_d[15]) );
  OAI21XL U30899 ( .A0(n28158), .A1(n27595), .B0(n27316), .Y(A6_d[16]) );
  OAI21XL U30900 ( .A0(n28158), .A1(n7114), .B0(n27318), .Y(A6_d[17]) );
  OAI21XL U30901 ( .A0(n28068), .A1(n7102), .B0(n27320), .Y(A6_d[18]) );
  OAI21XL U30902 ( .A0(n28158), .A1(n7090), .B0(n27322), .Y(A6_d[19]) );
  OAI21XL U30903 ( .A0(n28068), .A1(n7108), .B0(n27324), .Y(A6_d[20]) );
  OAI21XL U30904 ( .A0(n28068), .A1(n27625), .B0(n27326), .Y(A6_d[21]) );
  OAI21XL U30905 ( .A0(n28068), .A1(n27632), .B0(n27328), .Y(A6_d[22]) );
  OAI21XL U30906 ( .A0(n28158), .A1(n27638), .B0(n27330), .Y(A6_d[23]) );
  OAI21XL U30907 ( .A0(n28158), .A1(n7092), .B0(n27332), .Y(A6_d[24]) );
  OAI21XL U30908 ( .A0(n28068), .A1(n7094), .B0(n27334), .Y(A6_d[25]) );
  OAI21XL U30909 ( .A0(n28068), .A1(n27656), .B0(n27336), .Y(A6_d[26]) );
  OAI21XL U30910 ( .A0(n28068), .A1(n27667), .B0(n27338), .Y(A6_d[27]) );
  OAI21XL U30911 ( .A0(n28158), .A1(n27668), .B0(n27340), .Y(A6_d[28]) );
  OAI21XL U30912 ( .A0(n28068), .A1(n27674), .B0(n27342), .Y(A6_d[29]) );
  OAI21XL U30913 ( .A0(n28158), .A1(n27685), .B0(n27344), .Y(A6_d[30]) );
  OAI21XL U30914 ( .A0(n28068), .A1(n27692), .B0(n27346), .Y(A6_d[31]) );
  OAI21XL U30915 ( .A0(n28068), .A1(n27698), .B0(n27348), .Y(A6_d[32]) );
  OAI21XL U30916 ( .A0(n28068), .A1(n27699), .B0(n27350), .Y(A6_d[33]) );
  OAI21XL U30917 ( .A0(n28068), .A1(n27710), .B0(n27352), .Y(A6_d[34]) );
  OAI21XL U30918 ( .A0(n28158), .A1(n27711), .B0(n27354), .Y(A6_d[35]) );
  OAI21XL U30919 ( .A0(n28158), .A1(n27722), .B0(n27356), .Y(A6_d[36]) );
  OAI21XL U30920 ( .A0(n28068), .A1(n27728), .B0(n27358), .Y(A6_d[37]) );
  OAI21XL U30921 ( .A0(n28068), .A1(n7104), .B0(n27360), .Y(A6_d[38]) );
  OAI21XL U30922 ( .A0(n28158), .A1(n7116), .B0(n27362), .Y(A6_d[39]) );
  OAI21XL U30923 ( .A0(n28158), .A1(n27741), .B0(n27364), .Y(A6_d[40]) );
  OAI21XL U30924 ( .A0(n28068), .A1(n27752), .B0(n27366), .Y(A6_d[41]) );
  OAI21XL U30925 ( .A0(n28068), .A1(n27758), .B0(n27368), .Y(A6_d[42]) );
  OAI21XL U30926 ( .A0(n28068), .A1(n27764), .B0(n27370), .Y(A6_d[43]) );
  OAI21XL U30927 ( .A0(n28068), .A1(n7110), .B0(n27372), .Y(A6_d[44]) );
  OAI21XL U30928 ( .A0(n28068), .A1(n7086), .B0(n27374), .Y(A6_d[45]) );
  OAI21XL U30929 ( .A0(n28068), .A1(n27783), .B0(n27376), .Y(A6_d[46]) );
  OAI21XL U30930 ( .A0(n28068), .A1(n27784), .B0(n27378), .Y(A6_d[47]) );
  OAI21XL U30931 ( .A0(n28118), .A1(n27790), .B0(n27381), .Y(A6_d[48]) );
  OAI21XL U30932 ( .A0(n28158), .A1(n27801), .B0(n27383), .Y(A6_d[49]) );
  OAI21XL U30933 ( .A0(n28068), .A1(n27802), .B0(n27385), .Y(A6_d[50]) );
  OAI21XL U30934 ( .A0(n28068), .A1(n27808), .B0(n27388), .Y(A6_d[51]) );
  INVX4 U30935 ( .A(n27389), .Y(n28186) );
  OAI21XL U30936 ( .A0(n28271), .A1(n27498), .B0(n27392), .Y(A5_d[0]) );
  OAI21XL U30937 ( .A0(n28278), .A1(n27509), .B0(n27394), .Y(A5_d[1]) );
  OAI21XL U30938 ( .A0(n28271), .A1(n27515), .B0(n27396), .Y(A5_d[2]) );
  OAI21XL U30939 ( .A0(n28271), .A1(n27521), .B0(n27398), .Y(A5_d[3]) );
  OAI21XL U30940 ( .A0(n28278), .A1(n27527), .B0(n27400), .Y(A5_d[4]) );
  OAI21XL U30941 ( .A0(n28278), .A1(n27528), .B0(n27402), .Y(A5_d[5]) );
  OAI21XL U30942 ( .A0(n28179), .A1(n27539), .B0(n27404), .Y(A5_d[6]) );
  OAI21XL U30943 ( .A0(n27431), .A1(n27540), .B0(n27406), .Y(A5_d[7]) );
  OAI21XL U30944 ( .A0(n27431), .A1(n27551), .B0(n27408), .Y(A5_d[8]) );
  OAI21XL U30945 ( .A0(n28278), .A1(n27552), .B0(n27410), .Y(A5_d[9]) );
  OAI21XL U30946 ( .A0(n28278), .A1(n27558), .B0(n27412), .Y(A5_d[10]) );
  CLKINVX3 U30947 ( .A(n11891), .Y(n28278) );
  OAI21XL U30948 ( .A0(n28278), .A1(n7098), .B0(n27414), .Y(A5_d[11]) );
  OAI21XL U30949 ( .A0(n28179), .A1(n27571), .B0(n27416), .Y(A5_d[12]) );
  OAI21XL U30950 ( .A0(n28179), .A1(n27577), .B0(n27418), .Y(A5_d[13]) );
  OAI21XL U30951 ( .A0(n27431), .A1(n7112), .B0(n27420), .Y(A5_d[14]) );
  OAI21XL U30952 ( .A0(n28278), .A1(n7100), .B0(n27422), .Y(A5_d[15]) );
  OAI21XL U30953 ( .A0(n28271), .A1(n27600), .B0(n27424), .Y(A5_d[16]) );
  OAI21XL U30954 ( .A0(n27431), .A1(n7114), .B0(n27426), .Y(A5_d[17]) );
  OAI21XL U30955 ( .A0(n28271), .A1(n7102), .B0(n27428), .Y(A5_d[18]) );
  OAI21XL U30956 ( .A0(n27431), .A1(n7090), .B0(n27430), .Y(A5_d[19]) );
  OAI21XL U30957 ( .A0(n28179), .A1(n27619), .B0(n27433), .Y(A5_d[20]) );
  OAI21XL U30958 ( .A0(n28278), .A1(n27625), .B0(n27435), .Y(A5_d[21]) );
  OAI21XL U30959 ( .A0(n28278), .A1(n27632), .B0(n27437), .Y(A5_d[22]) );
  OAI21XL U30960 ( .A0(n28179), .A1(n27638), .B0(n27439), .Y(A5_d[23]) );
  OAI21XL U30961 ( .A0(n28179), .A1(n7092), .B0(n27441), .Y(A5_d[24]) );
  OAI21XL U30962 ( .A0(n28278), .A1(n7094), .B0(n27443), .Y(A5_d[25]) );
  OAI21XL U30963 ( .A0(n28179), .A1(n27661), .B0(n27445), .Y(A5_d[26]) );
  OAI21XL U30964 ( .A0(n28278), .A1(n27667), .B0(n27447), .Y(A5_d[27]) );
  OAI21XL U30965 ( .A0(n28278), .A1(n27673), .B0(n27449), .Y(A5_d[28]) );
  OAI21XL U30966 ( .A0(n28179), .A1(n27679), .B0(n27451), .Y(A5_d[29]) );
  OAI21XL U30967 ( .A0(n28278), .A1(n27680), .B0(n27453), .Y(A5_d[30]) );
  OAI21XL U30968 ( .A0(n28179), .A1(n27687), .B0(n27455), .Y(A5_d[31]) );
  OAI21XL U30969 ( .A0(n28179), .A1(n27693), .B0(n27457), .Y(A5_d[32]) );
  OAI21XL U30970 ( .A0(n28278), .A1(n27699), .B0(n27459), .Y(A5_d[33]) );
  OAI21XL U30971 ( .A0(n28179), .A1(n27705), .B0(n27461), .Y(A5_d[34]) );
  OAI21XL U30972 ( .A0(n28278), .A1(n27716), .B0(n27463), .Y(A5_d[35]) );
  OAI21XL U30973 ( .A0(n28179), .A1(n27722), .B0(n27465), .Y(A5_d[36]) );
  OAI21XL U30974 ( .A0(n28179), .A1(n27723), .B0(n27467), .Y(A5_d[37]) );
  OAI21XL U30975 ( .A0(n28278), .A1(n7104), .B0(n27469), .Y(A5_d[38]) );
  OAI21XL U30976 ( .A0(n28278), .A1(n27735), .B0(n27471), .Y(A5_d[39]) );
  OAI21XL U30977 ( .A0(n28179), .A1(n27741), .B0(n27473), .Y(A5_d[40]) );
  OAI21XL U30978 ( .A0(n28278), .A1(n27752), .B0(n27475), .Y(A5_d[41]) );
  OAI21XL U30979 ( .A0(n28179), .A1(n27753), .B0(n27477), .Y(A5_d[42]) );
  OAI21XL U30980 ( .A0(n28179), .A1(n27759), .B0(n27479), .Y(A5_d[43]) );
  OAI21XL U30981 ( .A0(n28179), .A1(n27765), .B0(n27481), .Y(A5_d[44]) );
  OAI21XL U30982 ( .A0(n28278), .A1(n7086), .B0(n27483), .Y(A5_d[45]) );
  OAI21XL U30983 ( .A0(n28179), .A1(n27778), .B0(n27485), .Y(A5_d[46]) );
  OAI21XL U30984 ( .A0(n28179), .A1(n27789), .B0(n27487), .Y(A5_d[47]) );
  OAI21XL U30985 ( .A0(n28179), .A1(n27790), .B0(n27489), .Y(A5_d[48]) );
  OAI21XL U30986 ( .A0(n28179), .A1(n27801), .B0(n27491), .Y(A5_d[49]) );
  OAI21XL U30987 ( .A0(n28179), .A1(n27807), .B0(n27493), .Y(A5_d[50]) );
  OAI21XL U30988 ( .A0(n28278), .A1(n27808), .B0(n27495), .Y(A5_d[51]) );
  OAI22XL U30989 ( .A0(n28579), .A1(n27499), .B0(n27772), .B1(n27498), .Y(
        n27500) );
  OAI21XL U30990 ( .A0(n28353), .A1(n27503), .B0(n27502), .Y(A4_d[0]) );
  OAI21XL U30991 ( .A0(n28295), .A1(n27509), .B0(n27508), .Y(A4_d[1]) );
  OAI21XL U30992 ( .A0(n28295), .A1(n27515), .B0(n27514), .Y(A4_d[2]) );
  OAI21XL U30993 ( .A0(n28295), .A1(n27521), .B0(n27520), .Y(A4_d[3]) );
  OAI21XL U30994 ( .A0(n28295), .A1(n27527), .B0(n27526), .Y(A4_d[4]) );
  OAI21XL U30995 ( .A0(n28353), .A1(n27533), .B0(n27532), .Y(A4_d[5]) );
  OAI22XL U30996 ( .A0(n27560), .A1(n27535), .B0(n27772), .B1(n27534), .Y(
        n27536) );
  OAI21XL U30997 ( .A0(n28353), .A1(n27539), .B0(n27538), .Y(A4_d[6]) );
  OAI21XL U30998 ( .A0(n28295), .A1(n27545), .B0(n27544), .Y(A4_d[7]) );
  OAI21XL U30999 ( .A0(n28353), .A1(n27551), .B0(n27550), .Y(A4_d[8]) );
  OAI21XL U31000 ( .A0(n28353), .A1(n27557), .B0(n27556), .Y(A4_d[9]) );
  OAI21XL U31001 ( .A0(n27686), .A1(n27564), .B0(n27563), .Y(A4_d[10]) );
  OAI21XL U31002 ( .A0(n28295), .A1(n7098), .B0(n27569), .Y(A4_d[11]) );
  OAI21XL U31003 ( .A0(n28295), .A1(n7106), .B0(n27575), .Y(A4_d[12]) );
  OAI21XL U31004 ( .A0(n28295), .A1(n27582), .B0(n27581), .Y(A4_d[13]) );
  OAI21XL U31005 ( .A0(n28353), .A1(n7112), .B0(n27587), .Y(A4_d[14]) );
  OAI21XL U31006 ( .A0(n28295), .A1(n7100), .B0(n27593), .Y(A4_d[15]) );
  OAI21XL U31007 ( .A0(n28295), .A1(n27600), .B0(n27599), .Y(A4_d[16]) );
  OAI22XL U31008 ( .A0(n28579), .A1(n27602), .B0(n27772), .B1(n27601), .Y(
        n27603) );
  OAI21XL U31009 ( .A0(n27686), .A1(n7114), .B0(n27605), .Y(A4_d[17]) );
  OAI21XL U31010 ( .A0(n28295), .A1(n7102), .B0(n27611), .Y(A4_d[18]) );
  OAI22XL U31011 ( .A0(n28579), .A1(n27614), .B0(n27772), .B1(n27613), .Y(
        n27615) );
  OAI21XL U31012 ( .A0(n28353), .A1(n7090), .B0(n27617), .Y(A4_d[19]) );
  OAI21XL U31013 ( .A0(n28295), .A1(n7108), .B0(n27623), .Y(A4_d[20]) );
  OAI22XL U31014 ( .A0(n28579), .A1(n27626), .B0(n27772), .B1(n27625), .Y(
        n27627) );
  OAI21XL U31015 ( .A0(n28353), .A1(n27630), .B0(n27629), .Y(A4_d[21]) );
  OAI22XL U31016 ( .A0(n28579), .A1(n27633), .B0(n27772), .B1(n27632), .Y(
        n27634) );
  OAI21XL U31017 ( .A0(n28353), .A1(n27637), .B0(n27636), .Y(A4_d[22]) );
  OAI21XL U31018 ( .A0(n28295), .A1(n27643), .B0(n27642), .Y(A4_d[23]) );
  OAI22XL U31019 ( .A0(n28579), .A1(n27645), .B0(n27772), .B1(n27644), .Y(
        n27646) );
  OAI21XL U31020 ( .A0(n27686), .A1(n7092), .B0(n27648), .Y(A4_d[24]) );
  OAI21XL U31021 ( .A0(n28295), .A1(n7094), .B0(n27654), .Y(A4_d[25]) );
  OAI22XL U31022 ( .A0(n28579), .A1(n27657), .B0(n27772), .B1(n27656), .Y(
        n27658) );
  OAI21XL U31023 ( .A0(n27686), .A1(n27661), .B0(n27660), .Y(A4_d[26]) );
  OAI21XL U31024 ( .A0(n28295), .A1(n27667), .B0(n27666), .Y(A4_d[27]) );
  OAI21XL U31025 ( .A0(n28295), .A1(n27673), .B0(n27672), .Y(A4_d[28]) );
  OAI22XL U31026 ( .A0(n28579), .A1(n27675), .B0(n27772), .B1(n27674), .Y(
        n27676) );
  OAI21XL U31027 ( .A0(n27686), .A1(n27679), .B0(n27678), .Y(A4_d[29]) );
  OAI22XL U31028 ( .A0(n28579), .A1(n27681), .B0(n27772), .B1(n27680), .Y(
        n27682) );
  OAI21XL U31029 ( .A0(n28353), .A1(n27685), .B0(n27684), .Y(A4_d[30]) );
  OAI21XL U31030 ( .A0(n28295), .A1(n27692), .B0(n27691), .Y(A4_d[31]) );
  OAI21XL U31031 ( .A0(n28295), .A1(n27698), .B0(n27697), .Y(A4_d[32]) );
  OAI22XL U31032 ( .A0(n28579), .A1(n27700), .B0(n27772), .B1(n27699), .Y(
        n27701) );
  OAI21XL U31033 ( .A0(n27686), .A1(n27704), .B0(n27703), .Y(A4_d[33]) );
  OAI21XL U31034 ( .A0(n28295), .A1(n27710), .B0(n27709), .Y(A4_d[34]) );
  OAI21XL U31035 ( .A0(n28295), .A1(n27716), .B0(n27715), .Y(A4_d[35]) );
  OAI22XL U31036 ( .A0(n28579), .A1(n27718), .B0(n27772), .B1(n27717), .Y(
        n27719) );
  OAI21XL U31037 ( .A0(n28353), .A1(n27722), .B0(n27721), .Y(A4_d[36]) );
  OAI21XL U31038 ( .A0(n28295), .A1(n27728), .B0(n27727), .Y(A4_d[37]) );
  OAI21XL U31039 ( .A0(n28295), .A1(n7104), .B0(n27733), .Y(A4_d[38]) );
  OAI22XL U31040 ( .A0(n28579), .A1(n27736), .B0(n27772), .B1(n27735), .Y(
        n27737) );
  OAI21XL U31041 ( .A0(n27686), .A1(n7116), .B0(n27739), .Y(A4_d[39]) );
  OAI21XL U31042 ( .A0(n28295), .A1(n27746), .B0(n27745), .Y(A4_d[40]) );
  OAI21XL U31043 ( .A0(n28295), .A1(n27752), .B0(n27751), .Y(A4_d[41]) );
  OAI21XL U31044 ( .A0(n28295), .A1(n27758), .B0(n27757), .Y(A4_d[42]) );
  OAI21XL U31045 ( .A0(n28295), .A1(n27764), .B0(n27763), .Y(A4_d[43]) );
  OAI21XL U31046 ( .A0(n28295), .A1(n7110), .B0(n27769), .Y(A4_d[44]) );
  OAI22XL U31047 ( .A0(n28579), .A1(n27773), .B0(n27772), .B1(n7086), .Y(
        n27774) );
  OAI21XL U31048 ( .A0(n27686), .A1(n27777), .B0(n27776), .Y(A4_d[45]) );
  OAI21XL U31049 ( .A0(n28295), .A1(n27783), .B0(n27782), .Y(A4_d[46]) );
  OAI22XL U31050 ( .A0(n28579), .A1(n27785), .B0(n27772), .B1(n27784), .Y(
        n27786) );
  OAI21XL U31051 ( .A0(n28353), .A1(n27789), .B0(n27788), .Y(A4_d[47]) );
  OAI21XL U31052 ( .A0(n28295), .A1(n27795), .B0(n27794), .Y(A4_d[48]) );
  OAI22XL U31053 ( .A0(n28579), .A1(n27797), .B0(n27772), .B1(n27796), .Y(
        n27798) );
  OAI21XL U31054 ( .A0(n28353), .A1(n27801), .B0(n27800), .Y(A4_d[49]) );
  OAI22XL U31055 ( .A0(n28579), .A1(n27803), .B0(n27772), .B1(n27802), .Y(
        n27804) );
  OAI21XL U31056 ( .A0(n28353), .A1(n27807), .B0(n27806), .Y(A4_d[50]) );
  OAI22XL U31057 ( .A0(n28579), .A1(n27809), .B0(n27772), .B1(n27808), .Y(
        n27810) );
  OAI21XL U31058 ( .A0(n28353), .A1(n27813), .B0(n27812), .Y(A4_d[51]) );
  AOI21XL U31059 ( .A0(OP2_done0), .A1(Q2[0]), .B0(n27816), .Y(n28287) );
  AOI21XL U31060 ( .A0(OP2_done0), .A1(Q1[0]), .B0(n27816), .Y(n28281) );
  OAI21XL U31061 ( .A0(n28287), .A1(n27264), .B0(n27818), .Y(A3_d[0]) );
  AOI21XL U31062 ( .A0(n27976), .A1(Q1[1]), .B0(n27820), .Y(n28288) );
  AOI21XL U31063 ( .A0(n27976), .A1(Q2[1]), .B0(n27820), .Y(n28294) );
  OAI21XL U31064 ( .A0(n28288), .A1(n7140), .B0(n27822), .Y(A3_d[1]) );
  AOI21XL U31065 ( .A0(n27976), .A1(Q1[2]), .B0(n27824), .Y(n28302) );
  AOI21XL U31066 ( .A0(OP2_done0), .A1(Q2[2]), .B0(n27824), .Y(n28296) );
  OAI21XL U31067 ( .A0(n28302), .A1(n7140), .B0(n27826), .Y(A3_d[2]) );
  AOI21XL U31068 ( .A0(OP2_done0), .A1(Q1[3]), .B0(n27828), .Y(n28309) );
  AOI21XL U31069 ( .A0(OP2_done0), .A1(Q2[3]), .B0(n27828), .Y(n28303) );
  OAI21XL U31070 ( .A0(n28309), .A1(n7140), .B0(n27830), .Y(A3_d[3]) );
  AOI21XL U31071 ( .A0(n27976), .A1(Q2[4]), .B0(n27832), .Y(n28310) );
  AOI21XL U31072 ( .A0(OP2_done0), .A1(Q1[4]), .B0(n27832), .Y(n28316) );
  OAI21XL U31073 ( .A0(n28310), .A1(n27264), .B0(n27834), .Y(A3_d[4]) );
  AOI21XL U31074 ( .A0(OP2_done0), .A1(Q2[5]), .B0(n27836), .Y(n28317) );
  AOI21XL U31075 ( .A0(n27976), .A1(Q1[5]), .B0(n27836), .Y(n28324) );
  OAI21XL U31076 ( .A0(n28317), .A1(n5823), .B0(n27838), .Y(A3_d[5]) );
  AOI21XL U31077 ( .A0(n27976), .A1(Q2[6]), .B0(n27840), .Y(n28325) );
  AOI21XL U31078 ( .A0(n27976), .A1(Q1[6]), .B0(n27840), .Y(n28331) );
  OAI21XL U31079 ( .A0(n28325), .A1(n27264), .B0(n27842), .Y(A3_d[6]) );
  AOI21XL U31080 ( .A0(OP2_done0), .A1(Q1[7]), .B0(n27844), .Y(n28332) );
  AOI21XL U31081 ( .A0(n27976), .A1(Q2[7]), .B0(n27844), .Y(n28338) );
  OAI21XL U31082 ( .A0(n28332), .A1(n7140), .B0(n27846), .Y(A3_d[7]) );
  AOI21XL U31083 ( .A0(n27976), .A1(Q2[8]), .B0(n27848), .Y(n28339) );
  AOI21XL U31084 ( .A0(n27976), .A1(Q1[8]), .B0(n27848), .Y(n28345) );
  OAI21XL U31085 ( .A0(n28339), .A1(n5823), .B0(n27850), .Y(A3_d[8]) );
  AOI21XL U31086 ( .A0(n27976), .A1(Q2[9]), .B0(n27852), .Y(n28346) );
  OAI21XL U31087 ( .A0(n28346), .A1(n5823), .B0(n27854), .Y(A3_d[9]) );
  AOI21XL U31088 ( .A0(OP2_done0), .A1(Q2[10]), .B0(n27856), .Y(n28354) );
  OAI21XL U31089 ( .A0(n28360), .A1(n7140), .B0(n27858), .Y(A3_d[10]) );
  OAI21X1 U31090 ( .A0(Q3[11]), .A1(n27861), .B0(n27860), .Y(n28362) );
  OAI21XL U31091 ( .A0(n28361), .A1(n27264), .B0(n27863), .Y(A3_d[11]) );
  OAI21X1 U31092 ( .A0(Q3[12]), .A1(n27866), .B0(n27865), .Y(n28369) );
  OAI21XL U31093 ( .A0(n28374), .A1(n7140), .B0(n27868), .Y(A3_d[12]) );
  OAI21X1 U31094 ( .A0(Q3[13]), .A1(n27871), .B0(n27870), .Y(n28376) );
  OAI21XL U31095 ( .A0(n28375), .A1(n5823), .B0(n27873), .Y(A3_d[13]) );
  OAI21X1 U31096 ( .A0(Q3[14]), .A1(n27876), .B0(n27875), .Y(n28383) );
  OAI21XL U31097 ( .A0(n28382), .A1(n5823), .B0(n27878), .Y(A3_d[14]) );
  OAI21XL U31098 ( .A0(Q1[15]), .A1(n27881), .B0(n27880), .Y(n28394) );
  OAI21X1 U31099 ( .A0(Q3[15]), .A1(n27881), .B0(n27880), .Y(n28390) );
  OAI21XL U31100 ( .A0(n28394), .A1(n7140), .B0(n27883), .Y(A3_d[15]) );
  OAI21X1 U31101 ( .A0(Q3[16]), .A1(n27886), .B0(n27885), .Y(n28396) );
  OAI21XL U31102 ( .A0(n28395), .A1(n7140), .B0(n27888), .Y(A3_d[16]) );
  OAI21X1 U31103 ( .A0(Q3[17]), .A1(n27891), .B0(n27890), .Y(n28402) );
  OAI21XL U31104 ( .A0(n28406), .A1(n27264), .B0(n27893), .Y(A3_d[17]) );
  OAI21X1 U31105 ( .A0(Q3[18]), .A1(n27896), .B0(n27895), .Y(n28408) );
  OAI21XL U31106 ( .A0(n28407), .A1(n7140), .B0(n27898), .Y(A3_d[18]) );
  OAI21X1 U31107 ( .A0(Q3[19]), .A1(n27901), .B0(n27900), .Y(n28414) );
  OAI21XL U31108 ( .A0(n28413), .A1(n27264), .B0(n27903), .Y(A3_d[19]) );
  OAI21X1 U31109 ( .A0(Q3[20]), .A1(n27906), .B0(n27905), .Y(n28420) );
  OAI21XL U31110 ( .A0(n28424), .A1(n7140), .B0(n27908), .Y(A3_d[20]) );
  OAI21X1 U31111 ( .A0(Q3[21]), .A1(n27911), .B0(n27910), .Y(n28426) );
  OAI21XL U31112 ( .A0(n28430), .A1(n7140), .B0(n27913), .Y(A3_d[21]) );
  OAI21X1 U31113 ( .A0(Q3[22]), .A1(n27916), .B0(n27915), .Y(n28432) );
  OAI21XL U31114 ( .A0(n28431), .A1(n7140), .B0(n27918), .Y(A3_d[22]) );
  OAI21X1 U31115 ( .A0(Q3[23]), .A1(n27921), .B0(n27920), .Y(n28438) );
  OAI21XL U31116 ( .A0(n28442), .A1(n5823), .B0(n27923), .Y(A3_d[23]) );
  OAI21X1 U31117 ( .A0(Q3[24]), .A1(n27926), .B0(n27925), .Y(n28444) );
  OAI21XL U31118 ( .A0(n28448), .A1(n5823), .B0(n27928), .Y(A3_d[24]) );
  OAI21X1 U31119 ( .A0(Q3[25]), .A1(n27931), .B0(n27930), .Y(n28450) );
  OAI21XL U31120 ( .A0(n28455), .A1(n7140), .B0(n27933), .Y(A3_d[25]) );
  AOI21XL U31121 ( .A0(OP2_done0), .A1(Q2[28]), .B0(n27935), .Y(n28456) );
  AOI21XL U31122 ( .A0(n27976), .A1(Q1[28]), .B0(n27935), .Y(n28462) );
  OAI21XL U31123 ( .A0(n28456), .A1(n5823), .B0(n27937), .Y(A3_d[26]) );
  AOI21XL U31124 ( .A0(n27976), .A1(Q2[29]), .B0(n27939), .Y(n28463) );
  AOI21XL U31125 ( .A0(n27976), .A1(Q1[29]), .B0(n27939), .Y(n28469) );
  OAI21XL U31126 ( .A0(n28463), .A1(n5823), .B0(n27941), .Y(A3_d[27]) );
  AOI21XL U31127 ( .A0(n27976), .A1(Q2[30]), .B0(n27943), .Y(n28470) );
  OAI21XL U31128 ( .A0(n28476), .A1(n7140), .B0(n27945), .Y(A3_d[28]) );
  AOI21XL U31129 ( .A0(n27976), .A1(Q2[31]), .B0(n27947), .Y(n28477) );
  OAI21XL U31130 ( .A0(n28483), .A1(n7140), .B0(n27949), .Y(A3_d[29]) );
  AOI21XL U31131 ( .A0(n27976), .A1(Q2[32]), .B0(n27951), .Y(n28484) );
  OAI21XL U31132 ( .A0(n28490), .A1(n7140), .B0(n27953), .Y(A3_d[30]) );
  AOI21XL U31133 ( .A0(OP2_done0), .A1(Q2[33]), .B0(n27955), .Y(n28491) );
  AOI21XL U31134 ( .A0(n27976), .A1(Q1[33]), .B0(n27955), .Y(n28497) );
  OAI21XL U31135 ( .A0(n28491), .A1(n5823), .B0(n27957), .Y(A3_d[31]) );
  AOI21XL U31136 ( .A0(n27976), .A1(Q2[34]), .B0(n27960), .Y(n28498) );
  AOI21XL U31137 ( .A0(n27976), .A1(Q1[34]), .B0(n27960), .Y(n28504) );
  OAI21XL U31138 ( .A0(n28498), .A1(n5823), .B0(n27962), .Y(A3_d[32]) );
  AOI21XL U31139 ( .A0(n27976), .A1(Q1[35]), .B0(n27964), .Y(n28511) );
  AOI21XL U31140 ( .A0(OP2_done0), .A1(Q2[35]), .B0(n27964), .Y(n28505) );
  OAI21XL U31141 ( .A0(n28511), .A1(n7140), .B0(n27966), .Y(A3_d[33]) );
  AOI21XL U31142 ( .A0(OP2_done0), .A1(Q2[36]), .B0(n27968), .Y(n28518) );
  AOI21XL U31143 ( .A0(OP2_done0), .A1(Q1[36]), .B0(n27968), .Y(n28512) );
  OAI21XL U31144 ( .A0(n28518), .A1(n5823), .B0(n27970), .Y(A3_d[34]) );
  AOI21XL U31145 ( .A0(n27976), .A1(Q2[37]), .B0(n27972), .Y(n28519) );
  OAI21XL U31146 ( .A0(n28525), .A1(n7140), .B0(n27974), .Y(A3_d[35]) );
  AOI21XL U31147 ( .A0(n27976), .A1(Q1[38]), .B0(n27977), .Y(n28532) );
  AOI21XL U31148 ( .A0(n27976), .A1(Q2[38]), .B0(n27977), .Y(n28526) );
  OAI21XL U31149 ( .A0(n28532), .A1(n7140), .B0(n27979), .Y(A3_d[36]) );
  OAI21X1 U31150 ( .A0(Q3[39]), .A1(n27982), .B0(n27981), .Y(n28534) );
  OAI21XL U31151 ( .A0(n28539), .A1(n7140), .B0(n27984), .Y(A3_d[37]) );
  OAI21X1 U31152 ( .A0(Q3[40]), .A1(n27987), .B0(n27986), .Y(n28541) );
  OAI21XL U31153 ( .A0(n28540), .A1(n5823), .B0(n27989), .Y(A3_d[38]) );
  OAI21X1 U31154 ( .A0(Q3[41]), .A1(n27992), .B0(n27991), .Y(n28548) );
  OAI21XL U31155 ( .A0(n28553), .A1(n5823), .B0(n27994), .Y(A3_d[39]) );
  OAI21X1 U31156 ( .A0(Q3[42]), .A1(n27997), .B0(n27996), .Y(n28555) );
  OAI21XL U31157 ( .A0(n28554), .A1(n7140), .B0(n27999), .Y(A3_d[40]) );
  OAI21X1 U31158 ( .A0(Q3[43]), .A1(n28002), .B0(n28001), .Y(n28562) );
  OAI21XL U31159 ( .A0(n28561), .A1(n7140), .B0(n28004), .Y(A3_d[41]) );
  OAI21X1 U31160 ( .A0(Q3[44]), .A1(n28007), .B0(n28006), .Y(n28568) );
  OAI21XL U31161 ( .A0(n28572), .A1(n5823), .B0(n28009), .Y(A3_d[42]) );
  OAI21X1 U31162 ( .A0(Q3[45]), .A1(n28012), .B0(n28011), .Y(n28574) );
  OAI21XL U31163 ( .A0(n28578), .A1(n5823), .B0(n28014), .Y(A3_d[43]) );
  OAI21X1 U31164 ( .A0(Q3[46]), .A1(n28017), .B0(n28016), .Y(n28581) );
  OAI21XL U31165 ( .A0(n28585), .A1(n7140), .B0(n28019), .Y(A3_d[44]) );
  OAI21X1 U31166 ( .A0(Q3[47]), .A1(n28022), .B0(n28021), .Y(n28587) );
  OAI21XL U31167 ( .A0(n28586), .A1(n5823), .B0(n28024), .Y(A3_d[45]) );
  OAI21X1 U31168 ( .A0(Q3[48]), .A1(n28027), .B0(n28026), .Y(n28593) );
  OAI21XL U31169 ( .A0(n28597), .A1(n5823), .B0(n28029), .Y(A3_d[46]) );
  OAI21X1 U31170 ( .A0(Q3[49]), .A1(n28032), .B0(n28031), .Y(n28599) );
  OAI21XL U31171 ( .A0(n28603), .A1(n27264), .B0(n28034), .Y(A3_d[47]) );
  OAI21X1 U31172 ( .A0(Q3[50]), .A1(n28037), .B0(n28036), .Y(n28605) );
  OAI21XL U31173 ( .A0(n28609), .A1(n5823), .B0(n28039), .Y(A3_d[48]) );
  OAI21X1 U31174 ( .A0(Q3[51]), .A1(n28042), .B0(n28041), .Y(n28611) );
  OAI21XL U31175 ( .A0(n28610), .A1(n7140), .B0(n28044), .Y(A3_d[49]) );
  OAI21X1 U31176 ( .A0(Q3[52]), .A1(n28047), .B0(n28046), .Y(n28617) );
  OAI21XL U31177 ( .A0(n28616), .A1(n7140), .B0(n28049), .Y(A3_d[50]) );
  OAI21X1 U31178 ( .A0(Q3[53]), .A1(n28053), .B0(n28052), .Y(n28623) );
  OAI21XL U31179 ( .A0(n28628), .A1(n7140), .B0(n28057), .Y(A3_d[51]) );
  OAI21XL U31180 ( .A0(n28281), .A1(n28068), .B0(n28059), .Y(A2_d[0]) );
  OAI21XL U31181 ( .A0(n28294), .A1(n28093), .B0(n28061), .Y(A2_d[1]) );
  CLKINVX3 U31182 ( .A(n5904), .Y(n28165) );
  OAI21XL U31183 ( .A0(n28302), .A1(n28068), .B0(n28063), .Y(A2_d[2]) );
  OAI21XL U31184 ( .A0(n28303), .A1(n28093), .B0(n28065), .Y(A2_d[3]) );
  OAI21XL U31185 ( .A0(n28310), .A1(n28093), .B0(n28067), .Y(A2_d[4]) );
  OAI21XL U31186 ( .A0(n28317), .A1(n28093), .B0(n28070), .Y(A2_d[5]) );
  CLKINVX3 U31187 ( .A(n5904), .Y(n28118) );
  OAI21XL U31188 ( .A0(n28331), .A1(n28068), .B0(n28072), .Y(A2_d[6]) );
  OAI21XL U31189 ( .A0(n28338), .A1(n28165), .B0(n28074), .Y(A2_d[7]) );
  OAI21XL U31190 ( .A0(n28345), .A1(n28068), .B0(n28076), .Y(A2_d[8]) );
  OAI21XL U31191 ( .A0(n28352), .A1(n28068), .B0(n28078), .Y(A2_d[9]) );
  OAI21XL U31192 ( .A0(n28360), .A1(n28068), .B0(n28080), .Y(A2_d[10]) );
  OAI21XL U31193 ( .A0(n28361), .A1(n28093), .B0(n28082), .Y(A2_d[11]) );
  OAI21XL U31194 ( .A0(n28368), .A1(n28165), .B0(n28084), .Y(A2_d[12]) );
  OAI21XL U31195 ( .A0(n28375), .A1(n28165), .B0(n28086), .Y(A2_d[13]) );
  OAI21XL U31196 ( .A0(n28382), .A1(n28165), .B0(n28088), .Y(A2_d[14]) );
  OAI21XL U31197 ( .A0(n28394), .A1(n27379), .B0(n28090), .Y(A2_d[15]) );
  OAI21XL U31198 ( .A0(n28400), .A1(n28093), .B0(n28092), .Y(A2_d[16]) );
  OAI21XL U31199 ( .A0(n28401), .A1(n28068), .B0(n28095), .Y(A2_d[17]) );
  OAI21XL U31200 ( .A0(n28407), .A1(n28068), .B0(n28097), .Y(A2_d[18]) );
  OAI21XL U31201 ( .A0(n28413), .A1(n28165), .B0(n28099), .Y(A2_d[19]) );
  OAI21XL U31202 ( .A0(n28424), .A1(n28068), .B0(n28101), .Y(A2_d[20]) );
  OAI21XL U31203 ( .A0(n28425), .A1(n28165), .B0(n28103), .Y(A2_d[21]) );
  OAI21XL U31204 ( .A0(n28436), .A1(n28165), .B0(n28105), .Y(A2_d[22]) );
  OAI21XL U31205 ( .A0(n28437), .A1(n28068), .B0(n28107), .Y(A2_d[23]) );
  OAI21XL U31206 ( .A0(n28448), .A1(n28165), .B0(n28109), .Y(A2_d[24]) );
  OAI21XL U31207 ( .A0(n28449), .A1(n28165), .B0(n28111), .Y(A2_d[25]) );
  OAI21XL U31208 ( .A0(n28456), .A1(n28165), .B0(n28113), .Y(A2_d[26]) );
  OAI21XL U31209 ( .A0(n28469), .A1(n28068), .B0(n28115), .Y(A2_d[27]) );
  OAI21XL U31210 ( .A0(n28476), .A1(n28068), .B0(n28117), .Y(A2_d[28]) );
  OAI21XL U31211 ( .A0(n28483), .A1(n28068), .B0(n28120), .Y(A2_d[29]) );
  OAI21XL U31212 ( .A0(n28490), .A1(n28068), .B0(n28122), .Y(A2_d[30]) );
  OAI21XL U31213 ( .A0(n28491), .A1(n28165), .B0(n28124), .Y(A2_d[31]) );
  OAI21XL U31214 ( .A0(n28504), .A1(n28068), .B0(n28127), .Y(A2_d[32]) );
  OAI21XL U31215 ( .A0(n28505), .A1(n28165), .B0(n28129), .Y(A2_d[33]) );
  OAI21XL U31216 ( .A0(n28512), .A1(n28068), .B0(n28131), .Y(A2_d[34]) );
  OAI21XL U31217 ( .A0(n28525), .A1(n28068), .B0(n28133), .Y(A2_d[35]) );
  OAI21XL U31218 ( .A0(n28526), .A1(n28165), .B0(n28135), .Y(A2_d[36]) );
  OAI21XL U31219 ( .A0(n28533), .A1(n28165), .B0(n28137), .Y(A2_d[37]) );
  OAI21XL U31220 ( .A0(n28546), .A1(n28068), .B0(n28140), .Y(A2_d[38]) );
  OAI21XL U31221 ( .A0(n28547), .A1(n28068), .B0(n28142), .Y(A2_d[39]) );
  OAI21XL U31222 ( .A0(n28554), .A1(n28068), .B0(n28145), .Y(A2_d[40]) );
  OAI21XL U31223 ( .A0(n28566), .A1(n28165), .B0(n28147), .Y(A2_d[41]) );
  OAI21XL U31224 ( .A0(n28572), .A1(n28158), .B0(n28149), .Y(A2_d[42]) );
  OAI21XL U31225 ( .A0(n28573), .A1(n28068), .B0(n28151), .Y(A2_d[43]) );
  OAI21XL U31226 ( .A0(n28580), .A1(n28158), .B0(n28153), .Y(A2_d[44]) );
  OAI21XL U31227 ( .A0(n28591), .A1(n27379), .B0(n28155), .Y(A2_d[45]) );
  OAI21XL U31228 ( .A0(n28597), .A1(n28158), .B0(n28157), .Y(A2_d[46]) );
  OAI21XL U31229 ( .A0(n28598), .A1(n28068), .B0(n28160), .Y(A2_d[47]) );
  OAI21XL U31230 ( .A0(n28604), .A1(n28068), .B0(n28162), .Y(A2_d[48]) );
  OAI21XL U31231 ( .A0(n28615), .A1(n28165), .B0(n28164), .Y(A2_d[49]) );
  OAI21XL U31232 ( .A0(n28616), .A1(n28068), .B0(n28167), .Y(A2_d[50]) );
  OAI21XL U31233 ( .A0(n28628), .A1(n28068), .B0(n28170), .Y(A2_d[51]) );
  OAI21XL U31234 ( .A0(n28287), .A1(n28179), .B0(n28172), .Y(A1_d[0]) );
  OAI21XL U31235 ( .A0(n28288), .A1(n5825), .B0(n28174), .Y(A1_d[1]) );
  OAI21XL U31236 ( .A0(n28302), .A1(n5825), .B0(n28176), .Y(A1_d[2]) );
  OAI21XL U31237 ( .A0(n28303), .A1(n28179), .B0(n28178), .Y(A1_d[3]) );
  OAI21XL U31238 ( .A0(n28316), .A1(n5825), .B0(n28181), .Y(A1_d[4]) );
  OAI21XL U31239 ( .A0(n28317), .A1(n28179), .B0(n28183), .Y(A1_d[5]) );
  OAI21XL U31240 ( .A0(n28325), .A1(n28179), .B0(n28185), .Y(A1_d[6]) );
  OAI21XL U31241 ( .A0(n28332), .A1(n5825), .B0(n28188), .Y(A1_d[7]) );
  OAI21XL U31242 ( .A0(n28339), .A1(n28179), .B0(n28190), .Y(A1_d[8]) );
  OAI21XL U31243 ( .A0(n28352), .A1(n5825), .B0(n28192), .Y(A1_d[9]) );
  OAI21XL U31244 ( .A0(n28354), .A1(n28179), .B0(n28194), .Y(A1_d[10]) );
  OAI21XL U31245 ( .A0(n28361), .A1(n28179), .B0(n28196), .Y(A1_d[11]) );
  CLKINVX3 U31246 ( .A(n11891), .Y(n28271) );
  OAI21XL U31247 ( .A0(n28374), .A1(n28271), .B0(n28198), .Y(A1_d[12]) );
  OAI21XL U31248 ( .A0(n28375), .A1(n28179), .B0(n28200), .Y(A1_d[13]) );
  OAI21XL U31249 ( .A0(n28388), .A1(n28271), .B0(n28202), .Y(A1_d[14]) );
  OAI21XL U31250 ( .A0(n28394), .A1(n5825), .B0(n28204), .Y(A1_d[15]) );
  OAI21XL U31251 ( .A0(n28395), .A1(n28271), .B0(n28206), .Y(A1_d[16]) );
  OAI21XL U31252 ( .A0(n28406), .A1(n28179), .B0(n28208), .Y(A1_d[17]) );
  OAI21XL U31253 ( .A0(n28412), .A1(n28179), .B0(n28210), .Y(A1_d[18]) );
  OAI21XL U31254 ( .A0(n28418), .A1(n28271), .B0(n28212), .Y(A1_d[19]) );
  OAI21XL U31255 ( .A0(n28419), .A1(n28179), .B0(n28214), .Y(A1_d[20]) );
  OAI21XL U31256 ( .A0(n28425), .A1(n28179), .B0(n28216), .Y(A1_d[21]) );
  OAI21XL U31257 ( .A0(n28436), .A1(n28179), .B0(n28218), .Y(A1_d[22]) );
  OAI21XL U31258 ( .A0(n28442), .A1(n28179), .B0(n28220), .Y(A1_d[23]) );
  OAI21XL U31259 ( .A0(n28443), .A1(n28271), .B0(n28222), .Y(A1_d[24]) );
  OAI21XL U31260 ( .A0(n28455), .A1(n28271), .B0(n28224), .Y(A1_d[25]) );
  OAI21XL U31261 ( .A0(n28462), .A1(n28271), .B0(n28226), .Y(A1_d[26]) );
  OAI21XL U31262 ( .A0(n28463), .A1(n28179), .B0(n28228), .Y(A1_d[27]) );
  OAI21XL U31263 ( .A0(n28476), .A1(n5825), .B0(n28230), .Y(A1_d[28]) );
  OAI21XL U31264 ( .A0(n28483), .A1(n28271), .B0(n28232), .Y(A1_d[29]) );
  OAI21XL U31265 ( .A0(n28490), .A1(n28271), .B0(n28234), .Y(A1_d[30]) );
  OAI21XL U31266 ( .A0(n28491), .A1(n28179), .B0(n28236), .Y(A1_d[31]) );
  OAI21XL U31267 ( .A0(n28498), .A1(n28179), .B0(n28239), .Y(A1_d[32]) );
  OAI21XL U31268 ( .A0(n28505), .A1(n28179), .B0(n28241), .Y(A1_d[33]) );
  OAI21XL U31269 ( .A0(n28512), .A1(n28271), .B0(n28243), .Y(A1_d[34]) );
  OAI21XL U31270 ( .A0(n28525), .A1(n28271), .B0(n28245), .Y(A1_d[35]) );
  OAI21XL U31271 ( .A0(n28526), .A1(n28179), .B0(n28247), .Y(A1_d[36]) );
  OAI21XL U31272 ( .A0(n28539), .A1(n28271), .B0(n28249), .Y(A1_d[37]) );
  OAI21XL U31273 ( .A0(n28540), .A1(n28179), .B0(n28251), .Y(A1_d[38]) );
  OAI21XL U31274 ( .A0(n28547), .A1(n28271), .B0(n28254), .Y(A1_d[39]) );
  OAI21XL U31275 ( .A0(n28554), .A1(n28271), .B0(n28256), .Y(A1_d[40]) );
  OAI21XL U31276 ( .A0(n28566), .A1(n28179), .B0(n28258), .Y(A1_d[41]) );
  OAI21XL U31277 ( .A0(n28567), .A1(n28271), .B0(n28260), .Y(A1_d[42]) );
  OAI21XL U31278 ( .A0(n28578), .A1(n28179), .B0(n28262), .Y(A1_d[43]) );
  OAI21XL U31279 ( .A0(n28585), .A1(n28271), .B0(n28264), .Y(A1_d[44]) );
  OAI21XL U31280 ( .A0(n28591), .A1(n28278), .B0(n28266), .Y(A1_d[45]) );
  OAI21XL U31281 ( .A0(n28592), .A1(n28278), .B0(n28268), .Y(A1_d[46]) );
  OAI21XL U31282 ( .A0(n28598), .A1(n28271), .B0(n28270), .Y(A1_d[47]) );
  OAI21XL U31283 ( .A0(n28609), .A1(n28179), .B0(n28273), .Y(A1_d[48]) );
  OAI21XL U31284 ( .A0(n28615), .A1(n28179), .B0(n28275), .Y(A1_d[49]) );
  OAI21XL U31285 ( .A0(n28616), .A1(n28278), .B0(n28277), .Y(A1_d[50]) );
  OAI21XL U31286 ( .A0(n28622), .A1(n28179), .B0(n28280), .Y(A1_d[51]) );
  OAI21XL U31287 ( .A0(n28287), .A1(n28353), .B0(n28286), .Y(A0_d[0]) );
  OAI21XL U31288 ( .A0(n28294), .A1(n28353), .B0(n28293), .Y(A0_d[1]) );
  OAI21XL U31289 ( .A0(n28302), .A1(n28295), .B0(n28301), .Y(A0_d[2]) );
  OAI21XL U31290 ( .A0(n28309), .A1(n28295), .B0(n28308), .Y(A0_d[3]) );
  OAI21XL U31291 ( .A0(n28316), .A1(n28295), .B0(n28315), .Y(A0_d[4]) );
  OAI21XL U31292 ( .A0(n28324), .A1(n28295), .B0(n28323), .Y(A0_d[5]) );
  OAI21XL U31293 ( .A0(n28331), .A1(n28295), .B0(n28330), .Y(A0_d[6]) );
  OAI21XL U31294 ( .A0(n28338), .A1(n28353), .B0(n28337), .Y(A0_d[7]) );
  OAI21XL U31295 ( .A0(n28345), .A1(n28295), .B0(n28344), .Y(A0_d[8]) );
  OAI21XL U31296 ( .A0(n28352), .A1(n28295), .B0(n28351), .Y(A0_d[9]) );
  OAI21XL U31297 ( .A0(n28360), .A1(n28295), .B0(n28359), .Y(A0_d[10]) );
  OAI21XL U31298 ( .A0(n28367), .A1(n28295), .B0(n28366), .Y(A0_d[11]) );
  OAI21XL U31299 ( .A0(n28374), .A1(n28295), .B0(n28373), .Y(A0_d[12]) );
  OAI21XL U31300 ( .A0(n28381), .A1(n28295), .B0(n28380), .Y(A0_d[13]) );
  OAI21XL U31301 ( .A0(n28388), .A1(n28295), .B0(n28387), .Y(A0_d[14]) );
  OAI21XL U31302 ( .A0(n28394), .A1(n28295), .B0(n28393), .Y(A0_d[15]) );
  OAI21XL U31303 ( .A0(n28400), .A1(n28353), .B0(n28399), .Y(A0_d[16]) );
  OAI21XL U31304 ( .A0(n28406), .A1(n28353), .B0(n28405), .Y(A0_d[17]) );
  OAI21XL U31305 ( .A0(n28412), .A1(n28353), .B0(n28411), .Y(A0_d[18]) );
  OAI21XL U31306 ( .A0(n28418), .A1(n28295), .B0(n28417), .Y(A0_d[19]) );
  OAI21XL U31307 ( .A0(n28424), .A1(n28295), .B0(n28423), .Y(A0_d[20]) );
  OAI21XL U31308 ( .A0(n28430), .A1(n28295), .B0(n28429), .Y(A0_d[21]) );
  OAI21XL U31309 ( .A0(n28436), .A1(n28353), .B0(n28435), .Y(A0_d[22]) );
  OAI21XL U31310 ( .A0(n28442), .A1(n28353), .B0(n28441), .Y(A0_d[23]) );
  OAI21XL U31311 ( .A0(n28448), .A1(n28353), .B0(n28447), .Y(A0_d[24]) );
  OAI21XL U31312 ( .A0(n28455), .A1(n28295), .B0(n28454), .Y(A0_d[25]) );
  OAI21XL U31313 ( .A0(n28462), .A1(n28295), .B0(n28461), .Y(A0_d[26]) );
  OAI21XL U31314 ( .A0(n28469), .A1(n28295), .B0(n28468), .Y(A0_d[27]) );
  OAI21XL U31315 ( .A0(n28476), .A1(n28295), .B0(n28475), .Y(A0_d[28]) );
  OAI21XL U31316 ( .A0(n28483), .A1(n28295), .B0(n28482), .Y(A0_d[29]) );
  OAI21XL U31317 ( .A0(n28490), .A1(n28295), .B0(n28489), .Y(A0_d[30]) );
  OAI21XL U31318 ( .A0(n28497), .A1(n28295), .B0(n28496), .Y(A0_d[31]) );
  OAI21XL U31319 ( .A0(n28504), .A1(n28295), .B0(n28503), .Y(A0_d[32]) );
  OAI21XL U31320 ( .A0(n28511), .A1(n28295), .B0(n28510), .Y(A0_d[33]) );
  OAI21XL U31321 ( .A0(n28518), .A1(n28353), .B0(n28517), .Y(A0_d[34]) );
  OAI21XL U31322 ( .A0(n28525), .A1(n28295), .B0(n28524), .Y(A0_d[35]) );
  OAI21XL U31323 ( .A0(n28532), .A1(n28295), .B0(n28531), .Y(A0_d[36]) );
  OAI21XL U31324 ( .A0(n28539), .A1(n28295), .B0(n28538), .Y(A0_d[37]) );
  OAI21XL U31325 ( .A0(n28546), .A1(n28295), .B0(n28545), .Y(A0_d[38]) );
  OAI21XL U31326 ( .A0(n28553), .A1(n28353), .B0(n28552), .Y(A0_d[39]) );
  OAI21XL U31327 ( .A0(n28560), .A1(n28353), .B0(n28559), .Y(A0_d[40]) );
  OAI21XL U31328 ( .A0(n28566), .A1(n28353), .B0(n28565), .Y(A0_d[41]) );
  OAI21XL U31329 ( .A0(n28572), .A1(n28353), .B0(n28571), .Y(A0_d[42]) );
  OAI21XL U31330 ( .A0(n28578), .A1(n28353), .B0(n28577), .Y(A0_d[43]) );
  OAI21XL U31331 ( .A0(n28585), .A1(n28295), .B0(n28584), .Y(A0_d[44]) );
  OAI21XL U31332 ( .A0(n28591), .A1(n28295), .B0(n28590), .Y(A0_d[45]) );
  OAI21XL U31333 ( .A0(n28597), .A1(n28353), .B0(n28596), .Y(A0_d[46]) );
  OAI21XL U31334 ( .A0(n28603), .A1(n28353), .B0(n28602), .Y(A0_d[47]) );
  OAI21XL U31335 ( .A0(n28609), .A1(n28353), .B0(n28608), .Y(A0_d[48]) );
  OAI21XL U31336 ( .A0(n28615), .A1(n28353), .B0(n28614), .Y(A0_d[49]) );
  OAI21XL U31337 ( .A0(n28621), .A1(n28353), .B0(n28620), .Y(A0_d[50]) );
  OAI21XL U31338 ( .A0(n28628), .A1(n28295), .B0(n28627), .Y(A0_d[51]) );
  OAI21XL U31341 ( .A0(n28630), .A1(cnt[0]), .B0(n28629), .Y(n5679) );
  AOI21XL U31342 ( .A0(n28674), .A1(n28633), .B0(n28631), .Y(n28632) );
  OAI21XL U31343 ( .A0(n28674), .A1(n28633), .B0(n28632), .Y(n5677) );
  OAI21XL U31344 ( .A0(n11956), .A1(Q3_addr[32]), .B0(n28644), .Y(n5536) );
  OAI21XL U31345 ( .A0(n11956), .A1(Q3_addr[33]), .B0(n28653), .Y(n5535) );
  OAI21XL U31346 ( .A0(n11956), .A1(Q3_addr[34]), .B0(n28646), .Y(n5534) );
  OAI21XL U31347 ( .A0(n11956), .A1(Q3_addr[35]), .B0(n28655), .Y(n5533) );
  OAI21XL U31348 ( .A0(n11956), .A1(Q3_addr[36]), .B0(n28647), .Y(n5532) );
  OAI21XL U31349 ( .A0(n11956), .A1(Q3_addr[37]), .B0(n28656), .Y(n5531) );
  OAI21XL U31350 ( .A0(n11956), .A1(Q1_addr[32]), .B0(n28644), .Y(n5530) );
  OAI21XL U31351 ( .A0(n11956), .A1(Q1_addr[33]), .B0(n28649), .Y(n5525) );
  OAI21XL U31352 ( .A0(n11956), .A1(Q1_addr[34]), .B0(n28646), .Y(n5520) );
  OAI21XL U31353 ( .A0(n11956), .A1(Q1_addr[35]), .B0(n28651), .Y(n5515) );
  OAI21XL U31354 ( .A0(n11956), .A1(Q1_addr[36]), .B0(n28647), .Y(n5510) );
  OAI21XL U31355 ( .A0(n11956), .A1(Q0_addr[32]), .B0(n28652), .Y(n5505) );
  OAI21XL U31356 ( .A0(n5834), .A1(Q0_addr[33]), .B0(n28649), .Y(n5503) );
  OAI21XL U31357 ( .A0(n11956), .A1(Q0_addr[34]), .B0(n28654), .Y(n5501) );
  OAI21XL U31358 ( .A0(n11956), .A1(Q0_addr[35]), .B0(n28651), .Y(n5499) );
  OAI21XL U31359 ( .A0(n11956), .A1(Q2_addr[32]), .B0(n28652), .Y(n5473) );
  OAI21XL U31360 ( .A0(n11956), .A1(Q2_addr[33]), .B0(n28653), .Y(n5468) );
  OAI21XL U31361 ( .A0(n11956), .A1(Q2_addr[34]), .B0(n28654), .Y(n5463) );
  OAI21XL U31362 ( .A0(n11956), .A1(Q2_addr[35]), .B0(n28655), .Y(n5458) );
  OAI21XL U31363 ( .A0(n11956), .A1(Q2_addr[37]), .B0(n28656), .Y(n5453) );
  OAI21XL U31364 ( .A0(n11956), .A1(Q3_addr[38]), .B0(n28658), .Y(n5404) );
  OAI21XL U31365 ( .A0(n5834), .A1(Q1_addr[38]), .B0(n28658), .Y(n5399) );
  OAI21XL U31366 ( .A0(n11956), .A1(Q1_addr[39]), .B0(n28660), .Y(n5394) );
  OAI21XL U31367 ( .A0(n11956), .A1(Q0_addr[39]), .B0(n28660), .Y(n5389) );
  OAI21XL U31368 ( .A0(n11956), .A1(Q1_addr[37]), .B0(n28662), .Y(n5384) );
  OAI21XL U31369 ( .A0(n11956), .A1(Q0_addr[37]), .B0(n28662), .Y(n5379) );
  OAI21XL U31370 ( .A0(n11956), .A1(Q0_addr[36]), .B0(n28664), .Y(n5374) );
  OAI21XL U31371 ( .A0(n11956), .A1(Q2_addr[36]), .B0(n28664), .Y(n5369) );
  OAI21XL U31372 ( .A0(n11956), .A1(Q0_addr[38]), .B0(n28668), .Y(n5364) );
  OAI21XL U31373 ( .A0(n11956), .A1(Q2_addr[38]), .B0(n28668), .Y(n5359) );
  OAI21XL U31374 ( .A0(n11956), .A1(Q3_addr[39]), .B0(n28670), .Y(n5354) );
  OAI21XL U31375 ( .A0(n11956), .A1(Q2_addr[39]), .B0(n28670), .Y(n5349) );
endmodule


module FFT2048_DW02_mult_2_stage_J1_20 ( A, B, TC, CLK, PRODUCT );
  input [15:0] A;
  input [26:0] B;
  output [42:0] PRODUCT;
  input TC, CLK;
  wire   n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, mult_x_1_n327, mult_x_1_n320, mult_x_1_n315,
         mult_x_1_n313, mult_x_1_n312, mult_x_1_n306, mult_x_1_n305,
         mult_x_1_n303, mult_x_1_n302, mult_x_1_n300, mult_x_1_n299,
         mult_x_1_n297, mult_x_1_n292, mult_x_1_n291, mult_x_1_n289,
         mult_x_1_n288, mult_x_1_n278, mult_x_1_n277, mult_x_1_n271,
         mult_x_1_n270, mult_x_1_n260, mult_x_1_n259, mult_x_1_n253,
         mult_x_1_n252, mult_x_1_n242, mult_x_1_n241, mult_x_1_n233,
         mult_x_1_n232, mult_x_1_n224, mult_x_1_n223, mult_x_1_n221,
         mult_x_1_n220, mult_x_1_n210, mult_x_1_n209, mult_x_1_n203,
         mult_x_1_n202, mult_x_1_n192, mult_x_1_n191, mult_x_1_n185,
         mult_x_1_n184, mult_x_1_n174, mult_x_1_n173, mult_x_1_n163,
         mult_x_1_n162, mult_x_1_n150, mult_x_1_n149, mult_x_1_n135,
         mult_x_1_n134, mult_x_1_n126, mult_x_1_n125, mult_x_1_n115,
         mult_x_1_n114, mult_x_1_n106, mult_x_1_n105, mult_x_1_n81,
         mult_x_1_n80, mult_x_1_n78, mult_x_1_n54, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238;

  DFFHQXL mult_x_1_clk_r_REG40_S1 ( .D(mult_x_1_n173), .CK(CLK), .Q(n1194) );
  DFFHQX1 mult_x_1_clk_r_REG6_S1 ( .D(mult_x_1_n302), .CK(CLK), .Q(n1227) );
  DFFHQXL mult_x_1_clk_r_REG42_S1 ( .D(mult_x_1_n162), .CK(CLK), .Q(n1192) );
  DFFHQXL mult_x_1_clk_r_REG36_S1 ( .D(mult_x_1_n191), .CK(CLK), .Q(n1198) );
  DFFHQX4 mult_x_1_clk_r_REG54_S1 ( .D(mult_x_1_n315), .CK(CLK), .Q(n1236) );
  DFFHQX4 mult_x_1_clk_r_REG3_S1 ( .D(mult_x_1_n305), .CK(CLK), .Q(n1229) );
  DFFHQX4 mult_x_1_clk_r_REG5_S1 ( .D(mult_x_1_n303), .CK(CLK), .Q(n1228) );
  DFFHQX4 mult_x_1_clk_r_REG7_S1 ( .D(mult_x_1_n297), .CK(CLK), .Q(n1224) );
  DFFHQX4 mult_x_1_clk_r_REG10_S1 ( .D(mult_x_1_n292), .CK(CLK), .Q(n1223) );
  DFFHQX4 mult_x_1_clk_r_REG11_S1 ( .D(mult_x_1_n291), .CK(CLK), .Q(n1222) );
  DFFHQX4 mult_x_1_clk_r_REG32_S1 ( .D(mult_x_1_n288), .CK(CLK), .Q(n1220) );
  DFFHQX4 mult_x_1_clk_r_REG29_S1 ( .D(mult_x_1_n278), .CK(CLK), .Q(n1219) );
  DFFHQX4 mult_x_1_clk_r_REG30_S1 ( .D(mult_x_1_n277), .CK(CLK), .Q(n1218) );
  DFFHQX4 mult_x_1_clk_r_REG28_S1 ( .D(mult_x_1_n270), .CK(CLK), .Q(n1216) );
  DFFHQX4 mult_x_1_clk_r_REG25_S1 ( .D(mult_x_1_n260), .CK(CLK), .Q(n1215) );
  DFFHQX4 mult_x_1_clk_r_REG14_S1 ( .D(mult_x_1_n252), .CK(CLK), .Q(n1212) );
  DFFHQXL clk_r_REG57_S1 ( .D(n1252), .CK(CLK), .Q(PRODUCT[12]) );
  DFFHQX4 mult_x_1_clk_r_REG56_S1 ( .D(mult_x_1_n320), .CK(CLK), .Q(n1237) );
  DFFHQXL mult_x_1_clk_r_REG20_S1 ( .D(mult_x_1_n223), .CK(CLK), .Q(n1206) );
  DFFHQXL clk_r_REG59_S1 ( .D(n1253), .CK(CLK), .Q(PRODUCT[11]) );
  DFFHQXL mult_x_1_clk_r_REG37_S1 ( .D(mult_x_1_n185), .CK(CLK), .Q(n1197) );
  DFFHQXL mult_x_1_clk_r_REG39_S1 ( .D(mult_x_1_n174), .CK(CLK), .Q(n1195) );
  DFFHQX1 mult_x_1_clk_r_REG55_S1 ( .D(mult_x_1_n81), .CK(CLK), .Q(n1234) );
  DFFHQXL clk_r_REG60_S1 ( .D(n1254), .CK(CLK), .Q(PRODUCT[10]) );
  DFFHQXL clk_r_REG61_S1 ( .D(n1255), .CK(CLK), .Q(PRODUCT[9]) );
  DFFHQXL mult_x_1_clk_r_REG38_S1 ( .D(mult_x_1_n184), .CK(CLK), .Q(n1196) );
  DFFHQXL mult_x_1_clk_r_REG41_S1 ( .D(mult_x_1_n163), .CK(CLK), .Q(n1193) );
  DFFHQXL mult_x_1_clk_r_REG23_S1 ( .D(mult_x_1_n210), .CK(CLK), .Q(n1203) );
  DFFHQXL mult_x_1_clk_r_REG24_S1 ( .D(mult_x_1_n209), .CK(CLK), .Q(n1202) );
  DFFHQXL mult_x_1_clk_r_REG12_S1 ( .D(mult_x_1_n54), .CK(CLK), .Q(n1181) );
  DFFHQX4 mult_x_1_clk_r_REG19_S1 ( .D(mult_x_1_n224), .CK(CLK), .Q(n1207) );
  DFFHQXL mult_x_1_clk_r_REG35_S1 ( .D(mult_x_1_n192), .CK(CLK), .Q(n1199) );
  DFFHQX1 mult_x_1_clk_r_REG15_S1 ( .D(mult_x_1_n242), .CK(CLK), .Q(n1211) );
  DFFHQXL clk_r_REG62_S1 ( .D(n1256), .CK(CLK), .Q(PRODUCT[8]) );
  DFFHQXL clk_r_REG63_S1 ( .D(n1257), .CK(CLK), .Q(PRODUCT[7]) );
  DFFHQXL clk_r_REG65_S1 ( .D(n1259), .CK(CLK), .Q(PRODUCT[5]) );
  DFFHQXL clk_r_REG67_S1 ( .D(n1261), .CK(CLK), .Q(PRODUCT[3]) );
  DFFHQXL clk_r_REG68_S1 ( .D(n1262), .CK(CLK), .Q(PRODUCT[2]) );
  DFFHQXL clk_r_REG69_S1 ( .D(n1263), .CK(CLK), .Q(PRODUCT[1]) );
  DFFHQXL clk_r_REG70_S1 ( .D(n1264), .CK(CLK), .Q(PRODUCT[0]) );
  DFFHQXL clk_r_REG64_S1 ( .D(n1258), .CK(CLK), .Q(PRODUCT[6]) );
  DFFHQXL clk_r_REG66_S1 ( .D(n1260), .CK(CLK), .Q(PRODUCT[4]) );
  DFFHQXL mult_x_1_clk_r_REG34_S1 ( .D(mult_x_1_n202), .CK(CLK), .Q(n1200) );
  DFFHQX2 mult_x_1_clk_r_REG16_S1 ( .D(mult_x_1_n241), .CK(CLK), .Q(n1210) );
  DFFHQXL mult_x_1_clk_r_REG4_S1 ( .D(mult_x_1_n78), .CK(CLK), .Q(n1230) );
  DFFHQXL mult_x_1_clk_r_REG17_S1 ( .D(mult_x_1_n233), .CK(CLK), .Q(n1209) );
  DFFHQX2 mult_x_1_clk_r_REG18_S1 ( .D(mult_x_1_n232), .CK(CLK), .Q(n1208) );
  DFFHQX1 mult_x_1_clk_r_REG22_S1 ( .D(mult_x_1_n220), .CK(CLK), .Q(n1204) );
  DFFHQXL mult_x_1_clk_r_REG33_S1 ( .D(mult_x_1_n203), .CK(CLK), .Q(n1201) );
  DFFHQXL mult_x_1_clk_r_REG43_S1 ( .D(mult_x_1_n150), .CK(CLK), .Q(n1191) );
  DFFHQXL mult_x_1_clk_r_REG44_S1 ( .D(mult_x_1_n149), .CK(CLK), .Q(n1190) );
  DFFHQXL mult_x_1_clk_r_REG45_S1 ( .D(mult_x_1_n135), .CK(CLK), .Q(n1189) );
  DFFHQXL mult_x_1_clk_r_REG46_S1 ( .D(mult_x_1_n134), .CK(CLK), .Q(n1188) );
  DFFHQXL mult_x_1_clk_r_REG47_S1 ( .D(mult_x_1_n126), .CK(CLK), .Q(n1187) );
  DFFHQXL mult_x_1_clk_r_REG48_S1 ( .D(mult_x_1_n125), .CK(CLK), .Q(n1186) );
  DFFHQXL mult_x_1_clk_r_REG49_S1 ( .D(mult_x_1_n115), .CK(CLK), .Q(n1185) );
  DFFHQXL mult_x_1_clk_r_REG50_S1 ( .D(mult_x_1_n114), .CK(CLK), .Q(n1184) );
  DFFHQXL mult_x_1_clk_r_REG51_S1 ( .D(mult_x_1_n106), .CK(CLK), .Q(n1183) );
  DFFHQXL mult_x_1_clk_r_REG52_S1 ( .D(mult_x_1_n105), .CK(CLK), .Q(n1182) );
  DFFHQX2 mult_x_1_clk_r_REG8_S1 ( .D(mult_x_1_n300), .CK(CLK), .Q(n1226) );
  DFFHQX2 mult_x_1_clk_r_REG27_S1 ( .D(mult_x_1_n271), .CK(CLK), .Q(n1217) );
  DFFHQX1 mult_x_1_clk_r_REG58_S1 ( .D(mult_x_1_n327), .CK(CLK), .Q(n1238) );
  DFFHQX4 mult_x_1_clk_r_REG31_S1 ( .D(mult_x_1_n289), .CK(CLK), .Q(n1221) );
  DFFHQX4 mult_x_1_clk_r_REG13_S1 ( .D(mult_x_1_n253), .CK(CLK), .Q(n1213) );
  DFFHQX4 mult_x_1_clk_r_REG26_S1 ( .D(mult_x_1_n259), .CK(CLK), .Q(n1214) );
  DFFHQX1 mult_x_1_clk_r_REG21_S1 ( .D(mult_x_1_n221), .CK(CLK), .Q(n1205) );
  DFFHQX1 mult_x_1_clk_r_REG2_S1 ( .D(mult_x_1_n312), .CK(CLK), .Q(n1231) );
  DFFHQX2 mult_x_1_clk_r_REG1_S1 ( .D(mult_x_1_n306), .CK(CLK), .Q(n1235) );
  DFFHQX2 mult_x_1_clk_r_REG9_S1 ( .D(mult_x_1_n299), .CK(CLK), .Q(n1225) );
  DFFHQX1 mult_x_1_clk_r_REG0_S1 ( .D(mult_x_1_n313), .CK(CLK), .Q(n1232) );
  DFFHQX1 mult_x_1_clk_r_REG53_S1 ( .D(mult_x_1_n80), .CK(CLK), .Q(n1233) );
  ADDFHX1 U1 ( .A(n582), .B(n581), .CI(n580), .CO(n569), .S(n611) );
  OAI2BB1X1 U2 ( .A0N(n607), .A1N(n30), .B0(n29), .Y(n581) );
  ADDFHX1 U3 ( .A(n465), .B(n464), .CI(n463), .CO(n439), .S(n470) );
  ADDFHX1 U4 ( .A(n777), .B(n776), .CI(n775), .CO(n778), .S(n790) );
  ADDFX2 U5 ( .A(n152), .B(n151), .CI(n150), .CO(n776), .S(n783) );
  CMPR32X1 U6 ( .A(n1012), .B(n1011), .C(n1010), .CO(n796), .S(n1020) );
  ADDFX2 U7 ( .A(n647), .B(n646), .CI(n645), .CO(n619), .S(n655) );
  ADDFHX1 U8 ( .A(n788), .B(n787), .CI(n786), .CO(n792), .S(n216) );
  ADDFX2 U9 ( .A(n211), .B(n210), .CI(n209), .CO(n784), .S(n786) );
  CMPR32X1 U10 ( .A(n660), .B(n659), .C(n658), .CO(n645), .S(n700) );
  CMPR32X1 U11 ( .A(n492), .B(n491), .C(n490), .CO(n484), .S(n545) );
  ADDFX2 U12 ( .A(n459), .B(n458), .CI(n457), .CO(n451), .S(n507) );
  INVXL U13 ( .A(n5), .Y(n6) );
  ADDFX2 U14 ( .A(n674), .B(n673), .CI(n672), .CO(n688), .S(n724) );
  CMPR32X1 U15 ( .A(n193), .B(n192), .C(n191), .CO(n186), .S(n1005) );
  ADDFX2 U16 ( .A(n603), .B(n602), .CI(n601), .CO(n593), .S(n659) );
  ADDFHX1 U17 ( .A(n943), .B(n942), .CI(n941), .CO(n950), .S(n949) );
  ADDFHX1 U18 ( .A(n972), .B(n971), .CI(n970), .CO(n974), .S(n951) );
  CMPR32X1 U19 ( .A(n176), .B(n175), .C(n174), .CO(n171), .S(n187) );
  ADDFHX1 U20 ( .A(n940), .B(n939), .CI(n938), .CO(n971), .S(n941) );
  CMPR32X1 U21 ( .A(n934), .B(n933), .C(n932), .CO(n959), .S(n943) );
  BUFX3 U22 ( .A(A[7]), .Y(n913) );
  BUFX3 U23 ( .A(A[1]), .Y(n854) );
  BUFX3 U24 ( .A(A[5]), .Y(n894) );
  BUFX3 U25 ( .A(A[3]), .Y(n920) );
  OAI21XL U26 ( .A0(n1179), .A1(n254), .B0(n253), .Y(n257) );
  XNOR2X1 U27 ( .A(n654), .B(n653), .Y(PRODUCT[23]) );
  XNOR2X1 U28 ( .A(n579), .B(n578), .Y(PRODUCT[25]) );
  XNOR2X2 U29 ( .A(n540), .B(n539), .Y(PRODUCT[26]) );
  XOR2X2 U30 ( .A(n1179), .B(n502), .Y(PRODUCT[27]) );
  XOR2X1 U31 ( .A(n791), .B(n33), .Y(PRODUCT[17]) );
  XOR2X1 U32 ( .A(n770), .B(n771), .Y(PRODUCT[19]) );
  OAI21X1 U33 ( .A0(n771), .A1(n1222), .B0(n1223), .Y(n754) );
  INVX4 U34 ( .A(n571), .Y(n771) );
  NOR2X2 U35 ( .A(n1218), .B(n1216), .Y(n218) );
  NAND3BX2 U36 ( .AN(n1236), .B(n1229), .C(n1224), .Y(n39) );
  INVXL U37 ( .A(n518), .Y(n5) );
  XNOR2X2 U38 ( .A(n754), .B(n753), .Y(PRODUCT[20]) );
  XNOR2XL U39 ( .A(n1031), .B(n1030), .Y(PRODUCT[37]) );
  XNOR2XL U40 ( .A(B[5]), .B(n854), .Y(n836) );
  XNOR2XL U41 ( .A(n920), .B(B[7]), .Y(n921) );
  XNOR2XL U42 ( .A(n1130), .B(n893), .Y(n627) );
  XNOR2XL U43 ( .A(n1081), .B(n1080), .Y(PRODUCT[38]) );
  XNOR2XL U44 ( .A(B[7]), .B(n894), .Y(n28) );
  XOR2XL U45 ( .A(n596), .B(n7), .Y(n23) );
  XNOR2XL U46 ( .A(A[13]), .B(n596), .Y(n372) );
  XNOR2XL U47 ( .A(n1043), .B(n893), .Y(n103) );
  XNOR2XL U48 ( .A(A[13]), .B(B[20]), .Y(n265) );
  XNOR2XL U49 ( .A(A[2]), .B(A[1]), .Y(n858) );
  XOR2XL U50 ( .A(n608), .B(n609), .Y(n14) );
  OAI2BB1X1 U51 ( .A0N(n26), .A1N(n25), .B0(n764), .Y(n24) );
  ADDFX2 U52 ( .A(n109), .B(n108), .CI(n107), .CO(n763), .S(n151) );
  ADDFX2 U53 ( .A(n1037), .B(n1036), .CI(n1035), .CO(n1053), .S(n290) );
  XNOR2XL U54 ( .A(n1149), .B(n1148), .Y(n1258) );
  XOR2XL U55 ( .A(n996), .B(n995), .Y(n1256) );
  XOR2XL U56 ( .A(n981), .B(n980), .Y(n1253) );
  NOR2XL U57 ( .A(n611), .B(n610), .Y(mult_x_1_n241) );
  INVX1 U58 ( .A(n977), .Y(n985) );
  INVX1 U59 ( .A(n986), .Y(n996) );
  INVX1 U60 ( .A(n619), .Y(n16) );
  ADDFHX1 U61 ( .A(n386), .B(n385), .CI(n384), .CO(n378), .S(n442) );
  NAND2X1 U62 ( .A(n216), .B(n215), .Y(n799) );
  INVXL U63 ( .A(n620), .Y(n17) );
  INVX1 U64 ( .A(n947), .Y(n983) );
  NAND2X1 U65 ( .A(n975), .B(n974), .Y(n1016) );
  INVXL U66 ( .A(n766), .Y(n25) );
  NAND2BXL U67 ( .AN(n634), .B(n21), .Y(n20) );
  NAND2XL U68 ( .A(n634), .B(n635), .Y(n19) );
  NAND2X1 U69 ( .A(n949), .B(n948), .Y(n982) );
  INVX1 U70 ( .A(n635), .Y(n21) );
  XNOR2X1 U71 ( .A(n913), .B(n1129), .Y(n263) );
  XNOR2X1 U72 ( .A(n894), .B(B[24]), .Y(n344) );
  INVXL U73 ( .A(n208), .Y(n38) );
  XNOR2X1 U74 ( .A(n913), .B(B[7]), .Y(n156) );
  XNOR2X1 U75 ( .A(n1130), .B(n919), .Y(n550) );
  NAND2X1 U76 ( .A(n238), .B(n229), .Y(n231) );
  INVX1 U77 ( .A(n854), .Y(n32) );
  NAND2X1 U78 ( .A(n769), .B(n1223), .Y(n770) );
  INVX1 U79 ( .A(n728), .Y(n729) );
  NAND2X1 U80 ( .A(n1172), .B(n1183), .Y(n1112) );
  INVX1 U81 ( .A(n1202), .Y(n435) );
  INVX1 U82 ( .A(n1182), .Y(n1172) );
  INVX1 U83 ( .A(n1212), .Y(n616) );
  XNOR2X1 U84 ( .A(A[12]), .B(A[11]), .Y(n81) );
  NAND2XL U85 ( .A(n500), .B(n499), .Y(mult_x_1_n221) );
  NOR2XL U86 ( .A(n500), .B(n499), .Y(mult_x_1_n220) );
  OAI21XL U87 ( .A0(n17), .A1(n16), .B0(n15), .Y(n610) );
  ADDFHX1 U88 ( .A(n472), .B(n471), .CI(n470), .CO(n466), .S(n500) );
  XNOR2X1 U89 ( .A(n991), .B(n990), .Y(n1255) );
  OAI21XL U90 ( .A0(n619), .A1(n620), .B0(n18), .Y(n15) );
  XOR2X1 U91 ( .A(n607), .B(n14), .Y(n18) );
  ADDFHX1 U92 ( .A(n443), .B(n442), .CI(n441), .CO(n427), .S(n472) );
  NAND2BXL U93 ( .AN(n609), .B(n31), .Y(n30) );
  NAND2X1 U94 ( .A(n1020), .B(n1019), .Y(n1033) );
  NAND2X1 U95 ( .A(n888), .B(n887), .Y(n993) );
  NOR2X1 U96 ( .A(n888), .B(n887), .Y(n992) );
  XNOR2X1 U97 ( .A(n894), .B(n1129), .Y(n260) );
  OAI22X1 U98 ( .A0(n445), .A1(n997), .B0(n446), .B1(n478), .Y(n477) );
  XNOR2X1 U99 ( .A(B[25]), .B(n854), .Y(n445) );
  ADDFHX1 U100 ( .A(n960), .B(n959), .CI(n958), .CO(n1008), .S(n970) );
  OAI22XL U101 ( .A0(n1094), .A1(n483), .B0(n1123), .B1(n450), .Y(n490) );
  XNOR2X1 U102 ( .A(n1180), .B(n1181), .Y(PRODUCT[40]) );
  OAI22X2 U103 ( .A0(n835), .A1(n931), .B0(n929), .B1(n8), .Y(n71) );
  NOR2X1 U104 ( .A(n237), .B(n231), .Y(n221) );
  OAI21X1 U105 ( .A0(n224), .A1(n231), .B0(n230), .Y(n232) );
  INVXL U106 ( .A(n1063), .Y(n48) );
  INVXL U107 ( .A(n667), .Y(n13) );
  NAND2X1 U108 ( .A(n399), .B(n1201), .Y(n400) );
  INVX1 U109 ( .A(n920), .Y(n7) );
  NAND2X1 U110 ( .A(n435), .B(n1203), .Y(n436) );
  NAND2X1 U111 ( .A(n255), .B(n1193), .Y(n256) );
  INVX1 U112 ( .A(n1186), .Y(n1073) );
  BUFX3 U113 ( .A(A[11]), .Y(n1043) );
  INVX1 U114 ( .A(n1190), .Y(n247) );
  INVX1 U115 ( .A(n1198), .Y(n363) );
  NAND2BX1 U116 ( .AN(n1227), .B(n1228), .Y(n33) );
  ADDFHX2 U117 ( .A(n392), .B(n391), .CI(n390), .CO(n367), .S(n402) );
  XOR3X2 U118 ( .A(n620), .B(n619), .C(n18), .Y(n649) );
  ADDFHX2 U119 ( .A(n429), .B(n428), .CI(n427), .CO(n403), .S(n438) );
  ADDFHX1 U120 ( .A(n505), .B(n504), .CI(n503), .CO(n499), .S(n532) );
  NAND2XL U121 ( .A(n52), .B(n734), .Y(n53) );
  XOR2X1 U122 ( .A(n55), .B(n732), .Y(n751) );
  OR2XL U123 ( .A(n1137), .B(n1136), .Y(n1139) );
  ADDFHX2 U124 ( .A(n688), .B(n687), .CI(n686), .CO(n656), .S(n698) );
  NOR2X1 U125 ( .A(n797), .B(n796), .Y(mult_x_1_n312) );
  XOR2X1 U126 ( .A(n733), .B(n734), .Y(n55) );
  INVX1 U127 ( .A(n608), .Y(n31) );
  NAND2X1 U128 ( .A(n609), .B(n608), .Y(n29) );
  ADDFHX2 U129 ( .A(n568), .B(n567), .CI(n566), .CO(n542), .S(n580) );
  NOR2X1 U130 ( .A(n1020), .B(n1019), .Y(n1032) );
  XOR2X2 U131 ( .A(n633), .B(n22), .Y(n687) );
  OAI2BB1X1 U132 ( .A0N(n20), .A1N(n633), .B0(n19), .Y(n647) );
  AOI21X1 U133 ( .A0(n1143), .A1(n1141), .B0(n884), .Y(n885) );
  XOR2X1 U134 ( .A(n634), .B(n635), .Y(n22) );
  NOR2X1 U135 ( .A(n890), .B(n889), .Y(n987) );
  NAND2BXL U136 ( .AN(n207), .B(n38), .Y(n36) );
  ADDFHX2 U137 ( .A(n202), .B(n201), .CI(n200), .CO(n213), .S(n1010) );
  NAND2XL U138 ( .A(n207), .B(n208), .Y(n35) );
  INVXL U139 ( .A(n882), .Y(n67) );
  ADDFHX1 U140 ( .A(n832), .B(n833), .CI(n834), .CO(n887), .S(n883) );
  ADDFHX1 U141 ( .A(n682), .B(n681), .CI(n680), .CO(n672), .S(n736) );
  OAI22X2 U142 ( .A0(n27), .A1(n929), .B0(n931), .B1(n23), .Y(n718) );
  OAI21X1 U143 ( .A0(n904), .A1(n10), .B0(n9), .Y(n198) );
  OAI22X1 U144 ( .A0(n915), .A1(n895), .B0(n28), .B1(n916), .Y(n966) );
  OAI22XL U145 ( .A0(n181), .A1(n916), .B0(n918), .B1(n28), .Y(n967) );
  NAND2BX1 U146 ( .AN(n588), .B(n13), .Y(n12) );
  XNOR2X1 U147 ( .A(n236), .B(n235), .Y(PRODUCT[36]) );
  OAI22X1 U148 ( .A0(n808), .A1(n929), .B0(n931), .B1(n8), .Y(n822) );
  OR2X2 U149 ( .A(n861), .B(n860), .Y(n859) );
  NAND2XL U150 ( .A(n57), .B(n48), .Y(n56) );
  NAND2BX1 U151 ( .AN(n165), .B(A[0]), .Y(n9) );
  XNOR2X1 U152 ( .A(n1113), .B(n1112), .Y(PRODUCT[39]) );
  OAI22XL U153 ( .A0(n1094), .A1(n592), .B0(n1123), .B1(n553), .Y(n601) );
  AND2XL U154 ( .A(n1165), .B(n1164), .Y(n1263) );
  BUFX3 U155 ( .A(B[11]), .Y(n628) );
  INVXL U156 ( .A(n58), .Y(n57) );
  OR2XL U157 ( .A(n1163), .B(n1162), .Y(n1165) );
  XNOR2X1 U158 ( .A(n249), .B(n248), .Y(PRODUCT[35]) );
  NAND2XL U159 ( .A(n51), .B(n48), .Y(n47) );
  NAND2XL U160 ( .A(n51), .B(n50), .Y(n49) );
  OAI21XL U161 ( .A0(n1179), .A1(n295), .B0(n294), .Y(n298) );
  AND2XL U162 ( .A(n1170), .B(n1172), .Y(n1176) );
  AND2XL U163 ( .A(n536), .B(n650), .Y(n43) );
  INVX1 U164 ( .A(n237), .Y(n362) );
  INVXL U165 ( .A(n926), .Y(n50) );
  NAND2X1 U166 ( .A(n780), .B(n1226), .Y(n781) );
  NAND2X1 U167 ( .A(n577), .B(n1211), .Y(n578) );
  NAND2X1 U168 ( .A(n616), .B(n1213), .Y(n617) );
  NAND2X1 U169 ( .A(n613), .B(n1215), .Y(n653) );
  NAND2X1 U170 ( .A(n695), .B(n1217), .Y(n696) );
  NAND2X1 U171 ( .A(n692), .B(n1219), .Y(n730) );
  INVX1 U172 ( .A(n62), .Y(n61) );
  NAND2X1 U173 ( .A(n74), .B(n1090), .Y(n1089) );
  INVX2 U174 ( .A(n258), .Y(n1118) );
  NAND2X1 U175 ( .A(n72), .B(n73), .Y(n895) );
  NAND2X1 U176 ( .A(n80), .B(n81), .Y(n1122) );
  AND2X2 U177 ( .A(n468), .B(n1205), .Y(n469) );
  INVX1 U178 ( .A(n1043), .Y(n196) );
  INVX1 U179 ( .A(A[15]), .Y(n258) );
  XNOR2X1 U180 ( .A(A[14]), .B(A[13]), .Y(n87) );
  INVX1 U181 ( .A(A[13]), .Y(n149) );
  XNOR2X1 U182 ( .A(n1238), .B(n1234), .Y(PRODUCT[13]) );
  NOR2X1 U183 ( .A(n1225), .B(n1228), .Y(n41) );
  INVX1 U184 ( .A(n1218), .Y(n692) );
  INVX1 U185 ( .A(n1192), .Y(n255) );
  NOR2X1 U186 ( .A(n1198), .B(n1196), .Y(n238) );
  INVX1 U187 ( .A(n1188), .Y(n1071) );
  AOI21X1 U188 ( .A0(n223), .A1(n395), .B0(n222), .Y(n224) );
  OAI21XL U189 ( .A0(n1179), .A1(n325), .B0(n324), .Y(n328) );
  OAI22X1 U190 ( .A0(n1063), .A1(n419), .B0(n1090), .B1(n382), .Y(n425) );
  NAND2X1 U191 ( .A(n1026), .B(n1016), .Y(n976) );
  NOR2X1 U192 ( .A(n975), .B(n974), .Y(n973) );
  XNOR2X1 U193 ( .A(n913), .B(B[4]), .Y(n924) );
  OAI22X1 U194 ( .A0(n1041), .A1(n669), .B0(n1042), .B1(n668), .Y(n719) );
  OAI21X1 U195 ( .A0(n1179), .A1(n434), .B0(n433), .Y(n437) );
  OAI22X1 U196 ( .A0(n931), .A1(n928), .B0(n929), .B1(n179), .Y(n968) );
  OAI22X1 U197 ( .A0(n904), .A1(n836), .B0(n830), .B1(n997), .Y(n840) );
  AOI21X1 U198 ( .A0(n892), .A1(n986), .B0(n891), .Y(n977) );
  AOI21X1 U199 ( .A0(n985), .A1(n983), .B0(n978), .Y(n981) );
  OAI22X1 U200 ( .A0(n1041), .A1(n115), .B0(n1042), .B1(n114), .Y(n125) );
  XNOR2X1 U201 ( .A(B[5]), .B(n920), .Y(n8) );
  XNOR2X1 U202 ( .A(B[5]), .B(n913), .Y(n922) );
  XNOR2X1 U203 ( .A(B[5]), .B(n894), .Y(n917) );
  XNOR2X1 U204 ( .A(B[5]), .B(n480), .Y(n177) );
  XNOR2X1 U205 ( .A(B[5]), .B(n1043), .Y(n104) );
  XNOR2X1 U206 ( .A(B[5]), .B(n1130), .Y(n665) );
  XNOR2X1 U207 ( .A(B[5]), .B(n1092), .Y(n118) );
  OAI22X1 U208 ( .A0(n902), .A1(n904), .B0(n997), .B1(n10), .Y(n899) );
  XNOR2X2 U209 ( .A(n628), .B(n854), .Y(n10) );
  AND2X2 U210 ( .A(n586), .B(n11), .Y(n594) );
  XOR2X1 U211 ( .A(n586), .B(n11), .Y(n635) );
  OAI21XL U212 ( .A0(n550), .A1(n1132), .B0(n12), .Y(n11) );
  OAI22X1 U213 ( .A0(n116), .A1(n931), .B0(n929), .B1(n23), .Y(n709) );
  XNOR2X1 U214 ( .A(B[21]), .B(n854), .Y(n587) );
  OAI2BB1X1 U215 ( .A0N(n766), .A1N(n765), .B0(n24), .Y(n756) );
  XNOR3X2 U216 ( .A(n766), .B(n26), .C(n764), .Y(n772) );
  INVX1 U217 ( .A(n765), .Y(n26) );
  OAI22X2 U218 ( .A0(n631), .A1(n929), .B0(n931), .B1(n27), .Y(n681) );
  XNOR2X4 U219 ( .A(n630), .B(n920), .Y(n27) );
  NOR2X1 U220 ( .A(n689), .B(n690), .Y(mult_x_1_n259) );
  NAND2X1 U221 ( .A(n531), .B(n532), .Y(mult_x_1_n224) );
  XNOR2X1 U222 ( .A(B[24]), .B(n854), .Y(n478) );
  OAI22X1 U223 ( .A0(n587), .A1(n904), .B0(n997), .B1(n549), .Y(n586) );
  XOR2X1 U224 ( .A(B[22]), .B(n32), .Y(n549) );
  AOI21X1 U225 ( .A0(n803), .A1(n1229), .B0(n1235), .Y(n791) );
  INVX1 U226 ( .A(n1236), .Y(n803) );
  NAND2X1 U227 ( .A(n223), .B(n432), .Y(n237) );
  NOR2X1 U228 ( .A(n1206), .B(n1204), .Y(n432) );
  NOR2X1 U229 ( .A(n1202), .B(n1200), .Y(n223) );
  XOR2X4 U230 ( .A(n34), .B(n469), .Y(PRODUCT[28]) );
  OAI21X2 U231 ( .A0(n1179), .A1(n1206), .B0(n1207), .Y(n34) );
  AND3X4 U232 ( .A(n65), .B(n63), .C(n64), .Y(n1179) );
  OAI2BB1X2 U233 ( .A0N(n36), .A1N(n206), .B0(n35), .Y(n787) );
  XOR2X1 U234 ( .A(n206), .B(n37), .Y(n212) );
  XNOR2X1 U235 ( .A(n207), .B(n38), .Y(n37) );
  XNOR2X1 U236 ( .A(B[15]), .B(n854), .Y(n88) );
  NOR2X1 U237 ( .A(n215), .B(n216), .Y(n798) );
  OAI21X1 U238 ( .A0(n771), .A1(n729), .B0(n61), .Y(n731) );
  NAND4BX4 U239 ( .AN(n41), .B(n40), .C(n39), .D(n1226), .Y(n571) );
  NAND2X2 U240 ( .A(n1235), .B(n1224), .Y(n40) );
  AND2X4 U241 ( .A(n728), .B(n218), .Y(n650) );
  NOR2X1 U242 ( .A(n1222), .B(n1220), .Y(n728) );
  XNOR2X1 U243 ( .A(n854), .B(B[10]), .Y(n902) );
  OAI22X1 U244 ( .A0(n925), .A1(n420), .B0(n923), .B1(n373), .Y(n411) );
  XNOR2X1 U245 ( .A(n913), .B(B[21]), .Y(n373) );
  ADDFX2 U246 ( .A(n644), .B(n643), .CI(n642), .CO(n660), .S(n701) );
  XNOR2X1 U247 ( .A(n894), .B(n630), .Y(n597) );
  XNOR2XL U248 ( .A(B[12]), .B(n854), .Y(n165) );
  XNOR2XL U249 ( .A(A[4]), .B(A[3]), .Y(n73) );
  INVXL U250 ( .A(n293), .Y(n250) );
  AOI21XL U251 ( .A0(n232), .A1(n1071), .B0(n1074), .Y(n1028) );
  XOR2XL U252 ( .A(n1043), .B(B[1]), .Y(n51) );
  AOI21XL U253 ( .A0(n232), .A1(n1076), .B0(n1075), .Y(n1077) );
  INVXL U254 ( .A(n1109), .Y(n1075) );
  NAND2XL U255 ( .A(n221), .B(n1076), .Y(n1078) );
  NAND2XL U256 ( .A(n1071), .B(n1189), .Y(n235) );
  INVXL U257 ( .A(n232), .Y(n233) );
  XNOR2XL U258 ( .A(n1130), .B(B[9]), .Y(n512) );
  OAI21XL U259 ( .A0(n771), .A1(n576), .B0(n575), .Y(n579) );
  INVXL U260 ( .A(n1210), .Y(n577) );
  XNOR2XL U261 ( .A(n1092), .B(B[14]), .Y(n414) );
  XNOR2XL U262 ( .A(n480), .B(n1117), .Y(n279) );
  XNOR2XL U263 ( .A(n480), .B(B[24]), .Y(n267) );
  XNOR2XL U264 ( .A(n1043), .B(B[20]), .Y(n300) );
  XNOR2XL U265 ( .A(n854), .B(B[6]), .Y(n830) );
  NAND2XL U266 ( .A(n221), .B(n1170), .Y(n1111) );
  XNOR2XL U267 ( .A(n1118), .B(B[19]), .Y(n278) );
  XNOR2XL U268 ( .A(n1043), .B(B[23]), .Y(n280) );
  XNOR2XL U269 ( .A(n1043), .B(B[24]), .Y(n1044) );
  XNOR2XL U270 ( .A(n480), .B(B[22]), .Y(n304) );
  XNOR2X1 U271 ( .A(n1118), .B(n630), .Y(n259) );
  XNOR2X1 U272 ( .A(n1118), .B(B[18]), .Y(n262) );
  XNOR2X1 U273 ( .A(n1043), .B(B[22]), .Y(n266) );
  XNOR2XL U274 ( .A(A[10]), .B(A[9]), .Y(n1090) );
  NAND2XL U275 ( .A(n221), .B(n1176), .Y(n1178) );
  XNOR2XL U276 ( .A(n1092), .B(n1129), .Y(n1120) );
  XNOR2XL U277 ( .A(n1118), .B(n1117), .Y(n1133) );
  XNOR2XL U278 ( .A(n1118), .B(B[24]), .Y(n1119) );
  XNOR2XL U279 ( .A(n1118), .B(B[23]), .Y(n1091) );
  OAI22XL U280 ( .A0(n895), .A1(n847), .B0(n916), .B1(n846), .Y(n872) );
  OAI22XL U281 ( .A0(n931), .A1(n865), .B0(n929), .B1(n845), .Y(n873) );
  AOI21XL U282 ( .A0(n1168), .A1(n1167), .B0(n879), .Y(n1140) );
  INVXL U283 ( .A(n1166), .Y(n879) );
  AOI21XL U284 ( .A0(n573), .A1(n536), .B0(n535), .Y(n537) );
  INVXL U285 ( .A(n1193), .Y(n239) );
  INVXL U286 ( .A(n1187), .Y(n1072) );
  NAND2XL U287 ( .A(n1073), .B(n1187), .Y(n1030) );
  NAND2XL U288 ( .A(n221), .B(n1071), .Y(n1029) );
  NAND2BXL U289 ( .AN(B[0]), .B(n480), .Y(n809) );
  XNOR2XL U290 ( .A(n1130), .B(B[10]), .Y(n479) );
  NAND2XL U291 ( .A(n247), .B(n1191), .Y(n248) );
  OAI21XL U292 ( .A0(n1179), .A1(n237), .B0(n224), .Y(n365) );
  XNOR2X2 U293 ( .A(n401), .B(n400), .Y(PRODUCT[30]) );
  OAI21XL U294 ( .A0(n1179), .A1(n398), .B0(n397), .Y(n401) );
  INVXL U295 ( .A(n1200), .Y(n399) );
  INVXL U296 ( .A(n395), .Y(n433) );
  INVXL U297 ( .A(n1204), .Y(n468) );
  OAI21XL U298 ( .A0(n771), .A1(n652), .B0(n651), .Y(n654) );
  NAND2XL U299 ( .A(n1079), .B(n1185), .Y(n1080) );
  INVXL U300 ( .A(n1184), .Y(n1079) );
  AOI21XL U301 ( .A0(n247), .A1(n239), .B0(n225), .Y(n226) );
  INVXL U302 ( .A(n1191), .Y(n225) );
  OAI21XL U303 ( .A0(n1208), .A1(n1211), .B0(n1209), .Y(n219) );
  NAND2X1 U304 ( .A(n573), .B(n66), .Y(n64) );
  XNOR2XL U305 ( .A(n480), .B(B[1]), .Y(n906) );
  XNOR2XL U306 ( .A(n913), .B(B[3]), .Y(n914) );
  XNOR2XL U307 ( .A(n920), .B(n919), .Y(n930) );
  XNOR2XL U308 ( .A(n480), .B(B[2]), .Y(n905) );
  XNOR2XL U309 ( .A(n1130), .B(B[12]), .Y(n409) );
  XNOR2XL U310 ( .A(n894), .B(B[23]), .Y(n383) );
  XNOR2XL U311 ( .A(n913), .B(B[20]), .Y(n420) );
  XNOR2XL U312 ( .A(n480), .B(B[14]), .Y(n551) );
  XNOR2XL U313 ( .A(n1092), .B(B[10]), .Y(n553) );
  XNOR2XL U314 ( .A(n1092), .B(B[9]), .Y(n592) );
  XNOR2XL U315 ( .A(n1092), .B(n919), .Y(n632) );
  XNOR2XL U316 ( .A(n1043), .B(B[10]), .Y(n637) );
  XNOR2XL U317 ( .A(n913), .B(B[14]), .Y(n638) );
  XNOR2X1 U318 ( .A(n1092), .B(B[7]), .Y(n670) );
  XNOR2XL U319 ( .A(n1043), .B(B[9]), .Y(n677) );
  XNOR2XL U320 ( .A(n913), .B(B[13]), .Y(n678) );
  XNOR2XL U321 ( .A(n480), .B(B[10]), .Y(n669) );
  XNOR2XL U322 ( .A(n1092), .B(n893), .Y(n671) );
  XNOR2XL U323 ( .A(n894), .B(B[14]), .Y(n676) );
  XOR2XL U324 ( .A(n919), .B(n196), .Y(n59) );
  XNOR2XL U325 ( .A(n913), .B(B[12]), .Y(n679) );
  XNOR2XL U326 ( .A(n1130), .B(B[1]), .Y(n90) );
  XNOR2XL U327 ( .A(B[4]), .B(n1043), .Y(n58) );
  XNOR2XL U328 ( .A(n1092), .B(B[2]), .Y(n136) );
  XNOR2XL U329 ( .A(n894), .B(n919), .Y(n181) );
  XNOR2XL U330 ( .A(n480), .B(B[3]), .Y(n896) );
  XNOR2XL U331 ( .A(n480), .B(B[4]), .Y(n194) );
  NAND2BXL U332 ( .AN(B[0]), .B(n1043), .Y(n195) );
  XNOR2XL U333 ( .A(n1043), .B(B[3]), .Y(n159) );
  XNOR2XL U334 ( .A(n1092), .B(B[1]), .Y(n157) );
  NOR2BXL U335 ( .AN(B[0]), .B(n1123), .Y(n199) );
  OAI21XL U336 ( .A0(n166), .A1(n926), .B0(n47), .Y(n197) );
  XNOR2XL U337 ( .A(n913), .B(B[19]), .Y(n456) );
  XNOR2XL U338 ( .A(n1043), .B(B[14]), .Y(n488) );
  XNOR2X1 U339 ( .A(n913), .B(B[18]), .Y(n489) );
  XNOR2XL U340 ( .A(n1092), .B(B[12]), .Y(n483) );
  XNOR2XL U341 ( .A(n480), .B(B[15]), .Y(n513) );
  XNOR2X1 U342 ( .A(n1092), .B(n628), .Y(n515) );
  XNOR2X1 U343 ( .A(n913), .B(n630), .Y(n521) );
  XNOR2XL U344 ( .A(n913), .B(n596), .Y(n559) );
  XNOR2XL U345 ( .A(n480), .B(B[9]), .Y(n114) );
  XNOR2X1 U346 ( .A(n1043), .B(B[7]), .Y(n83) );
  XNOR2XL U347 ( .A(n894), .B(B[13]), .Y(n82) );
  XNOR2XL U348 ( .A(n913), .B(n628), .Y(n84) );
  XNOR2XL U349 ( .A(n920), .B(B[12]), .Y(n141) );
  XNOR2XL U350 ( .A(n913), .B(n919), .Y(n146) );
  XNOR2XL U351 ( .A(n913), .B(B[10]), .Y(n105) );
  XNOR2XL U352 ( .A(n913), .B(B[9]), .Y(n106) );
  XNOR2XL U353 ( .A(n480), .B(n919), .Y(n115) );
  XNOR2XL U354 ( .A(n1092), .B(B[4]), .Y(n119) );
  XNOR2XL U355 ( .A(n1092), .B(B[3]), .Y(n97) );
  XNOR2XL U356 ( .A(n1130), .B(B[14]), .Y(n346) );
  XNOR2XL U357 ( .A(n913), .B(B[2]), .Y(n813) );
  XNOR2XL U358 ( .A(n854), .B(B[8]), .Y(n811) );
  XNOR2XL U359 ( .A(n894), .B(B[4]), .Y(n805) );
  NAND2BXL U360 ( .AN(B[0]), .B(n913), .Y(n806) );
  XNOR2XL U361 ( .A(n913), .B(B[1]), .Y(n817) );
  XNOR2XL U362 ( .A(n480), .B(n1129), .Y(n1039) );
  CMPR32X1 U363 ( .A(n423), .B(n422), .C(n421), .CO(n415), .S(n474) );
  OAI2BB1XL U364 ( .A0N(n997), .A1N(n904), .B0(n377), .Y(n421) );
  OAI22XL U365 ( .A0(n1134), .A1(n409), .B0(n1132), .B1(n376), .Y(n422) );
  OAI22X1 U366 ( .A0(n1041), .A1(n412), .B0(n1042), .B1(n375), .Y(n423) );
  OAI22XL U367 ( .A0(n1094), .A1(n450), .B0(n1123), .B1(n414), .Y(n457) );
  CMPR32X1 U368 ( .A(n6), .B(n517), .C(n516), .CO(n530), .S(n567) );
  XNOR2XL U369 ( .A(n1118), .B(B[20]), .Y(n1038) );
  XNOR2XL U370 ( .A(n480), .B(B[23]), .Y(n299) );
  XNOR2X1 U371 ( .A(n1043), .B(B[21]), .Y(n270) );
  OAI2BB1XL U372 ( .A0N(n916), .A1N(n918), .B0(n261), .Y(n308) );
  OAI22XL U373 ( .A0(n1134), .A1(n302), .B0(n1132), .B1(n259), .Y(n310) );
  INVXL U374 ( .A(n260), .Y(n261) );
  OAI2BB1XL U375 ( .A0N(n923), .A1N(n600), .B0(n264), .Y(n281) );
  OAI22XL U376 ( .A0(n1134), .A1(n262), .B0(n1132), .B1(n278), .Y(n283) );
  INVXL U377 ( .A(n263), .Y(n264) );
  OAI22XL U378 ( .A0(n1041), .A1(n267), .B0(n1042), .B1(n279), .Y(n284) );
  OAI22XL U379 ( .A0(n1094), .A1(n265), .B0(n1123), .B1(n277), .Y(n286) );
  OAI22X1 U380 ( .A0(n925), .A1(n340), .B0(n923), .B1(n301), .Y(n336) );
  OAI22XL U381 ( .A0(n1041), .A1(n341), .B0(n1042), .B1(n304), .Y(n332) );
  XNOR2XL U382 ( .A(n920), .B(B[4]), .Y(n835) );
  OAI22XL U383 ( .A0(n918), .A1(n838), .B0(n916), .B1(n837), .Y(n848) );
  NOR2BXL U384 ( .AN(B[0]), .B(n923), .Y(n841) );
  OAI22XL U385 ( .A0(n918), .A1(n846), .B0(n916), .B1(n831), .Y(n839) );
  OAI2BB1XL U386 ( .A0N(n1090), .A1N(n1089), .B0(n1088), .Y(n1095) );
  OAI22XL U387 ( .A0(n1134), .A1(n1086), .B0(n1132), .B1(n1091), .Y(n1096) );
  INVXL U388 ( .A(n1087), .Y(n1088) );
  OAI22XL U389 ( .A0(n1094), .A1(n1060), .B0(n1123), .B1(n1082), .Y(n1085) );
  INVXL U390 ( .A(n1097), .Y(n1083) );
  OAI22XL U391 ( .A0(n1134), .A1(n1061), .B0(n1132), .B1(n1086), .Y(n1084) );
  OAI22XL U392 ( .A0(n1094), .A1(n1045), .B0(n1123), .B1(n1060), .Y(n1065) );
  OAI22XL U393 ( .A0(n1063), .A1(n1044), .B0(n1090), .B1(n1062), .Y(n1066) );
  NOR2BXL U394 ( .AN(B[0]), .B(n916), .Y(n876) );
  OAI22XL U395 ( .A0(n931), .A1(n866), .B0(n929), .B1(n865), .Y(n874) );
  OAI22XL U396 ( .A0(n904), .A1(n864), .B0(n863), .B1(n997), .Y(n875) );
  ADDFX2 U397 ( .A(n825), .B(n824), .CI(n823), .CO(n889), .S(n888) );
  OAI21XL U398 ( .A0(n70), .A1(n69), .B0(n68), .Y(n824) );
  INVXL U399 ( .A(n829), .Y(n69) );
  INVXL U400 ( .A(n71), .Y(n70) );
  NAND2XL U401 ( .A(n1143), .B(n1147), .Y(n886) );
  OAI22XL U402 ( .A0(n1134), .A1(n1133), .B0(n1132), .B1(n1131), .Y(n1135) );
  OAI2BB1XL U403 ( .A0N(n1123), .A1N(n1122), .B0(n1121), .Y(n1126) );
  OAI22XL U404 ( .A0(n1134), .A1(n1119), .B0(n1132), .B1(n1133), .Y(n1127) );
  INVXL U405 ( .A(n1120), .Y(n1121) );
  NOR2XL U406 ( .A(n870), .B(n869), .Y(n1150) );
  INVXL U407 ( .A(n1155), .Y(n862) );
  NAND2XL U408 ( .A(n870), .B(n869), .Y(n1151) );
  OAI22XL U409 ( .A0(n904), .A1(B[0]), .B0(n850), .B1(n997), .Y(n1163) );
  NAND2XL U410 ( .A(n851), .B(n904), .Y(n1162) );
  NAND2BXL U411 ( .AN(B[0]), .B(n854), .Y(n851) );
  NAND2XL U412 ( .A(n1163), .B(n1162), .Y(n1164) );
  NAND2XL U413 ( .A(n878), .B(n877), .Y(n1166) );
  INVXL U414 ( .A(n1140), .Y(n1148) );
  INVXL U415 ( .A(n1108), .Y(n1076) );
  INVXL U416 ( .A(n1189), .Y(n1074) );
  INVXL U417 ( .A(n1195), .Y(n240) );
  NAND2XL U418 ( .A(n432), .B(n435), .Y(n398) );
  AOI21XL U419 ( .A0(n323), .A1(n363), .B0(n322), .Y(n324) );
  INVXL U420 ( .A(n1199), .Y(n322) );
  AOI21XL U421 ( .A0(n533), .A1(n573), .B0(n534), .Y(n575) );
  AOI21XL U422 ( .A0(n573), .A1(n613), .B0(n612), .Y(n614) );
  INVXL U423 ( .A(n1215), .Y(n612) );
  INVXL U424 ( .A(n1219), .Y(n691) );
  NAND2XL U425 ( .A(n1071), .B(n1073), .Y(n1108) );
  XNOR2X1 U426 ( .A(n854), .B(B[18]), .Y(n664) );
  XNOR2XL U427 ( .A(n1130), .B(B[4]), .Y(n666) );
  XNOR2X1 U428 ( .A(n1130), .B(B[7]), .Y(n588) );
  XNOR2XL U429 ( .A(n1130), .B(B[3]), .Y(n111) );
  INVXL U430 ( .A(n1208), .Y(n538) );
  XNOR2X2 U431 ( .A(n618), .B(n617), .Y(PRODUCT[24]) );
  OAI21XL U432 ( .A0(n771), .A1(n615), .B0(n614), .Y(n618) );
  NAND2XL U433 ( .A(n801), .B(n1232), .Y(n802) );
  NOR2XL U434 ( .A(n1108), .B(n1184), .Y(n1170) );
  INVXL U435 ( .A(n480), .Y(n810) );
  NOR2BXL U436 ( .AN(B[0]), .B(n926), .Y(n912) );
  OAI22XL U437 ( .A0(n1041), .A1(n906), .B0(n1042), .B1(n905), .Y(n910) );
  OAI22X1 U438 ( .A0(n904), .A1(n903), .B0(n902), .B1(n997), .Y(n911) );
  XNOR2X1 U439 ( .A(n480), .B(B[18]), .Y(n412) );
  XNOR2X1 U440 ( .A(n1043), .B(n628), .Y(n598) );
  XNOR2XL U441 ( .A(n913), .B(B[15]), .Y(n599) );
  XNOR2XL U442 ( .A(n894), .B(B[9]), .Y(n180) );
  OAI21XL U443 ( .A0(n927), .A1(n1063), .B0(n49), .Y(n962) );
  OAI22XL U444 ( .A0(n925), .A1(n922), .B0(n923), .B1(n167), .Y(n969) );
  OAI22XL U445 ( .A0(n1094), .A1(n149), .B0(n1123), .B1(n148), .Y(n163) );
  OAI22XL U446 ( .A0(n904), .A1(n165), .B0(n147), .B1(n997), .Y(n164) );
  NAND2BXL U447 ( .AN(B[0]), .B(n1092), .Y(n148) );
  XNOR2X1 U448 ( .A(n480), .B(n630), .Y(n448) );
  XNOR2XL U449 ( .A(n1092), .B(B[13]), .Y(n450) );
  OAI22X1 U450 ( .A0(n904), .A1(n511), .B0(n478), .B1(n997), .Y(n510) );
  XNOR2XL U451 ( .A(n894), .B(B[10]), .Y(n145) );
  NAND2BXL U452 ( .AN(B[0]), .B(n1130), .Y(n89) );
  XNOR2XL U453 ( .A(n480), .B(B[20]), .Y(n347) );
  XNOR2XL U454 ( .A(n1043), .B(B[19]), .Y(n342) );
  XNOR2X1 U455 ( .A(n480), .B(B[21]), .Y(n341) );
  XNOR2XL U456 ( .A(n1118), .B(n596), .Y(n302) );
  NAND2BXL U457 ( .AN(B[0]), .B(n894), .Y(n837) );
  INVXL U458 ( .A(n1174), .Y(n1175) );
  INVXL U459 ( .A(n1183), .Y(n1171) );
  NAND3X1 U460 ( .A(n650), .B(n66), .C(n571), .Y(n65) );
  NOR2X1 U461 ( .A(n219), .B(n44), .Y(n63) );
  CMPR32X1 U462 ( .A(n909), .B(n908), .C(n907), .CO(n938), .S(n946) );
  OAI22XL U463 ( .A0(n918), .A1(n805), .B0(n916), .B1(n917), .Y(n907) );
  XNOR2XL U464 ( .A(n1043), .B(n1129), .Y(n1087) );
  XNOR2X1 U465 ( .A(n1118), .B(B[22]), .Y(n1086) );
  XNOR2XL U466 ( .A(n1043), .B(n1117), .Y(n1062) );
  XNOR2XL U467 ( .A(A[13]), .B(B[23]), .Y(n1060) );
  CMPR32X1 U468 ( .A(n426), .B(n425), .C(n424), .CO(n443), .S(n473) );
  OAI22X1 U469 ( .A0(n931), .A1(n413), .B0(n858), .B1(n381), .Y(n426) );
  OAI22XL U470 ( .A0(n925), .A1(n456), .B0(n923), .B1(n420), .Y(n460) );
  CMPR32X1 U471 ( .A(n486), .B(n46), .C(n484), .CO(n498), .S(n529) );
  XOR2XL U472 ( .A(n444), .B(n60), .Y(n486) );
  BUFX1 U473 ( .A(n485), .Y(n46) );
  OAI22XL U474 ( .A0(n1094), .A1(n553), .B0(n1123), .B1(n515), .Y(n560) );
  CMPR32X1 U475 ( .A(n606), .B(n605), .C(n604), .CO(n623), .S(n658) );
  OAI22XL U476 ( .A0(n925), .A1(n599), .B0(n923), .B1(n559), .Y(n604) );
  OAI22XL U477 ( .A0(n1063), .A1(n598), .B0(n926), .B1(n558), .Y(n605) );
  OAI22XL U478 ( .A0(n918), .A1(n597), .B0(n916), .B1(n557), .Y(n606) );
  OAI22XL U479 ( .A0(n600), .A1(n638), .B0(n923), .B1(n599), .Y(n642) );
  OAI22X1 U480 ( .A0(n918), .A1(n636), .B0(n916), .B1(n597), .Y(n644) );
  OAI22XL U481 ( .A0(n1063), .A1(n637), .B0(n926), .B1(n598), .Y(n643) );
  OAI22XL U482 ( .A0(n1094), .A1(n632), .B0(n1123), .B1(n592), .Y(n639) );
  ADDFX2 U483 ( .A(n713), .B(n712), .CI(n711), .CO(n725), .S(n748) );
  OAI22XL U484 ( .A0(n1094), .A1(n670), .B0(n1123), .B1(n632), .Y(n680) );
  OAI22XL U485 ( .A0(n925), .A1(n678), .B0(n923), .B1(n638), .Y(n683) );
  OAI22XL U486 ( .A0(n1063), .A1(n677), .B0(n926), .B1(n637), .Y(n684) );
  CMPR32X1 U487 ( .A(n719), .B(n718), .C(n717), .CO(n711), .S(n759) );
  OAI22XL U488 ( .A0(n1094), .A1(n671), .B0(n1123), .B1(n670), .Y(n717) );
  OAI22XL U489 ( .A0(n925), .A1(n679), .B0(n923), .B1(n678), .Y(n720) );
  OAI22X1 U490 ( .A0(n677), .A1(n926), .B0(n1063), .B1(n59), .Y(n721) );
  OAI22XL U491 ( .A0(n1094), .A1(n118), .B0(n1123), .B1(n671), .Y(n708) );
  OAI22XL U492 ( .A0(n1041), .A1(n114), .B0(n1042), .B1(n669), .Y(n710) );
  OAI22XL U493 ( .A0(n925), .A1(n84), .B0(n923), .B1(n679), .Y(n714) );
  OAI22X1 U494 ( .A0(n83), .A1(n1063), .B0(n926), .B1(n59), .Y(n715) );
  OAI22XL U495 ( .A0(n1094), .A1(n136), .B0(n1123), .B1(n97), .Y(n142) );
  OAI22XL U496 ( .A0(n1134), .A1(n91), .B0(n1132), .B1(n90), .Y(n143) );
  OAI22X1 U497 ( .A0(n897), .A1(n140), .B0(n1042), .B1(n96), .Y(n144) );
  ADDFX2 U498 ( .A(n184), .B(n183), .CI(n182), .CO(n155), .S(n185) );
  OAI22X1 U499 ( .A0(n159), .A1(n1063), .B0(n926), .B1(n58), .Y(n183) );
  OAI22XL U500 ( .A0(n897), .A1(n177), .B0(n1042), .B1(n140), .Y(n184) );
  NOR2BXL U501 ( .AN(B[0]), .B(n1132), .Y(n176) );
  OAI22XL U502 ( .A0(n1094), .A1(n157), .B0(n1123), .B1(n136), .Y(n174) );
  OAI22XL U503 ( .A0(n1041), .A1(n896), .B0(n1042), .B1(n194), .Y(n957) );
  OAI22XL U504 ( .A0(n1094), .A1(n158), .B0(n1123), .B1(n157), .Y(n189) );
  OAI22XL U505 ( .A0(n1063), .A1(n166), .B0(n926), .B1(n159), .Y(n188) );
  OAI22XL U506 ( .A0(n925), .A1(n167), .B0(n923), .B1(n156), .Y(n190) );
  CMPR32X1 U507 ( .A(n162), .B(n161), .C(n160), .CO(n153), .S(n201) );
  OAI22XL U508 ( .A0(n918), .A1(n180), .B0(n916), .B1(n145), .Y(n162) );
  OAI22XL U509 ( .A0(n925), .A1(n156), .B0(n923), .B1(n146), .Y(n161) );
  OAI22XL U510 ( .A0(n925), .A1(n489), .B0(n923), .B1(n456), .Y(n493) );
  OAI22XL U511 ( .A0(n918), .A1(n487), .B0(n916), .B1(n454), .Y(n495) );
  CMPR32X1 U512 ( .A(n527), .B(n526), .C(n525), .CO(n546), .S(n583) );
  OAI22XL U513 ( .A0(n1063), .A1(n520), .B0(n1090), .B1(n488), .Y(n526) );
  OAI22XL U514 ( .A0(n918), .A1(n519), .B0(n916), .B1(n487), .Y(n527) );
  OAI22XL U515 ( .A0(n1094), .A1(n515), .B0(n1123), .B1(n483), .Y(n522) );
  CMPR32X1 U516 ( .A(n565), .B(n564), .C(n563), .CO(n585), .S(n621) );
  OAI22XL U517 ( .A0(n1063), .A1(n558), .B0(n926), .B1(n520), .Y(n564) );
  OAI22XL U518 ( .A0(n918), .A1(n557), .B0(n916), .B1(n519), .Y(n565) );
  CMPR32X1 U519 ( .A(n595), .B(n594), .C(n593), .CO(n609), .S(n646) );
  ADDFX2 U520 ( .A(n556), .B(n555), .CI(n554), .CO(n568), .S(n608) );
  OAI22XL U521 ( .A0(n1094), .A1(n119), .B0(n1123), .B1(n118), .Y(n123) );
  OAI22XL U522 ( .A0(n931), .A1(n117), .B0(n929), .B1(n116), .Y(n124) );
  OAI22XL U523 ( .A0(n925), .A1(n105), .B0(n923), .B1(n84), .Y(n126) );
  OAI22XL U524 ( .A0(n925), .A1(n146), .B0(n923), .B1(n106), .Y(n168) );
  OAI21XL U525 ( .A0(n104), .A1(n926), .B0(n56), .Y(n169) );
  OAI22XL U526 ( .A0(n925), .A1(n106), .B0(n923), .B1(n105), .Y(n120) );
  OAI22XL U527 ( .A0(n1094), .A1(n97), .B0(n1123), .B1(n119), .Y(n99) );
  OAI22XL U528 ( .A0(n1089), .A1(n300), .B0(n1090), .B1(n270), .Y(n305) );
  OAI22XL U529 ( .A0(n1122), .A1(n303), .B0(n1123), .B1(n269), .Y(n306) );
  OAI22XL U530 ( .A0(n925), .A1(n301), .B0(n923), .B1(n268), .Y(n307) );
  OAI22XL U531 ( .A0(n1122), .A1(n269), .B0(n1123), .B1(n265), .Y(n273) );
  CMPR32X1 U532 ( .A(n389), .B(n388), .C(n387), .CO(n407), .S(n441) );
  OAI22XL U533 ( .A0(n1041), .A1(n375), .B0(n1042), .B1(n347), .Y(n387) );
  OAI22XL U534 ( .A0(n1134), .A1(n376), .B0(n1132), .B1(n346), .Y(n388) );
  OAI22XL U535 ( .A0(n925), .A1(n373), .B0(n923), .B1(n345), .Y(n389) );
  AND2XL U536 ( .A(n444), .B(n60), .Y(n453) );
  OAI22XL U537 ( .A0(n1122), .A1(n374), .B0(n1123), .B1(n372), .Y(n417) );
  OR2XL U538 ( .A(n411), .B(n410), .Y(n416) );
  OAI22XL U539 ( .A0(n925), .A1(n345), .B0(n923), .B1(n340), .Y(n351) );
  OAI2BB1XL U540 ( .A0N(n858), .A1N(n591), .B0(n331), .Y(n348) );
  XNOR2XL U541 ( .A(n854), .B(B[4]), .Y(n863) );
  NOR2BXL U542 ( .AN(B[0]), .B(n1042), .Y(n816) );
  OAI22XL U543 ( .A0(n925), .A1(n817), .B0(n923), .B1(n813), .Y(n814) );
  OAI22XL U544 ( .A0(n925), .A1(n807), .B0(n923), .B1(n806), .Y(n826) );
  INVXL U545 ( .A(n913), .Y(n807) );
  OAI2BB1XL U546 ( .A0N(n1042), .A1N(n1041), .B0(n1040), .Y(n1057) );
  OAI22XL U547 ( .A0(n1134), .A1(n1038), .B0(n1132), .B1(n1061), .Y(n1059) );
  INVXL U548 ( .A(n1039), .Y(n1040) );
  ADDFX2 U549 ( .A(n498), .B(n497), .CI(n496), .CO(n471), .S(n503) );
  ADDFX2 U550 ( .A(n737), .B(n736), .CI(n735), .CO(n723), .S(n757) );
  ADDFX2 U551 ( .A(n760), .B(n759), .CI(n758), .CO(n747), .S(n774) );
  ADDFX2 U552 ( .A(n1015), .B(n1014), .CI(n1013), .CO(n1019), .S(n1018) );
  OAI22XL U553 ( .A0(n1134), .A1(n278), .B0(n1132), .B1(n1038), .Y(n1047) );
  OAI22XL U554 ( .A0(n1094), .A1(n277), .B0(n1123), .B1(n1045), .Y(n1048) );
  INVXL U555 ( .A(n1058), .Y(n1046) );
  OAI22XL U556 ( .A0(n1063), .A1(n280), .B0(n1090), .B1(n1044), .Y(n1051) );
  OAI22XL U557 ( .A0(n1041), .A1(n304), .B0(n1042), .B1(n299), .Y(n313) );
  OAI22XL U558 ( .A0(n1063), .A1(n270), .B0(n1090), .B1(n266), .Y(n276) );
  OAI22XL U559 ( .A0(n1134), .A1(n259), .B0(n1132), .B1(n262), .Y(n275) );
  CMPR32X1 U560 ( .A(n316), .B(n315), .C(n314), .CO(n317), .S(n357) );
  INVX1 U561 ( .A(A[0]), .Y(n85) );
  OAI22XL U562 ( .A0(n904), .A1(n850), .B0(n855), .B1(n997), .Y(n853) );
  NOR2BXL U563 ( .AN(B[0]), .B(n929), .Y(n852) );
  OAI22XL U564 ( .A0(n931), .A1(n7), .B0(n858), .B1(n857), .Y(n860) );
  NAND2BXL U565 ( .AN(B[0]), .B(n920), .Y(n857) );
  ADDFX2 U566 ( .A(n844), .B(n45), .CI(n842), .CO(n882), .S(n881) );
  OAI22XL U567 ( .A0(n931), .A1(n845), .B0(n929), .B1(n835), .Y(n844) );
  OR2X2 U568 ( .A(n1018), .B(n1017), .Y(n1070) );
  NAND2X1 U569 ( .A(n1018), .B(n1017), .Y(n1069) );
  INVXL U570 ( .A(n973), .Y(n1026) );
  INVX1 U571 ( .A(n1022), .Y(n1027) );
  OAI22XL U572 ( .A0(n1134), .A1(n1091), .B0(n1132), .B1(n1119), .Y(n1116) );
  INVXL U573 ( .A(n1128), .Y(n1115) );
  OAI22XL U574 ( .A0(n1094), .A1(n1082), .B0(n1123), .B1(n1093), .Y(n1105) );
  CMPR32X1 U575 ( .A(n1056), .B(n1055), .C(n1054), .CO(n1068), .S(n1052) );
  NAND2X1 U576 ( .A(n54), .B(n53), .Y(n726) );
  OAI21XL U577 ( .A0(n52), .A1(n734), .B0(n732), .Y(n54) );
  BUFX1 U578 ( .A(n733), .Y(n52) );
  OAI2BB1X1 U579 ( .A0N(n1016), .A1N(n1069), .B0(n1070), .Y(n1024) );
  NOR2XL U580 ( .A(n853), .B(n852), .Y(n1158) );
  NAND2XL U581 ( .A(n853), .B(n852), .Y(n1159) );
  NAND2XL U582 ( .A(n861), .B(n860), .Y(n1155) );
  NAND2BX1 U583 ( .AN(n883), .B(n67), .Y(n1143) );
  NAND2XL U584 ( .A(n1139), .B(n1138), .Y(mult_x_1_n54) );
  NAND2XL U585 ( .A(n1137), .B(n1136), .Y(n1138) );
  INVXL U586 ( .A(n1135), .Y(n1136) );
  NAND2XL U587 ( .A(n989), .B(n988), .Y(n990) );
  XNOR2X1 U588 ( .A(n985), .B(n984), .Y(n1254) );
  OAI21XL U589 ( .A0(n1025), .A1(n1027), .B0(n1024), .Y(mult_x_1_n320) );
  NOR2XL U590 ( .A(n1125), .B(n1124), .Y(mult_x_1_n105) );
  NAND2XL U591 ( .A(n1125), .B(n1124), .Y(mult_x_1_n106) );
  NOR2XL U592 ( .A(n1099), .B(n1098), .Y(mult_x_1_n114) );
  NAND2XL U593 ( .A(n1099), .B(n1098), .Y(mult_x_1_n115) );
  NOR2XL U594 ( .A(n1107), .B(n1106), .Y(mult_x_1_n125) );
  NAND2XL U595 ( .A(n1107), .B(n1106), .Y(mult_x_1_n126) );
  NOR2XL U596 ( .A(n1068), .B(n1067), .Y(mult_x_1_n134) );
  NAND2XL U597 ( .A(n1068), .B(n1067), .Y(mult_x_1_n135) );
  NOR2XL U598 ( .A(n1053), .B(n1052), .Y(mult_x_1_n149) );
  NAND2XL U599 ( .A(n1053), .B(n1052), .Y(mult_x_1_n150) );
  NAND2XL U600 ( .A(n1034), .B(n1033), .Y(mult_x_1_n80) );
  INVXL U601 ( .A(n1032), .Y(n1034) );
  NOR2X1 U602 ( .A(n793), .B(n792), .Y(mult_x_1_n302) );
  XOR2XL U603 ( .A(n1154), .B(n1153), .Y(n1260) );
  NAND2XL U604 ( .A(n1152), .B(n1151), .Y(n1154) );
  INVXL U605 ( .A(n1150), .Y(n1152) );
  NAND2XL U606 ( .A(n1147), .B(n1146), .Y(n1149) );
  NOR2BXL U607 ( .AN(B[0]), .B(n997), .Y(n1264) );
  XOR2XL U608 ( .A(n1161), .B(n1164), .Y(n1262) );
  NAND2XL U609 ( .A(n1160), .B(n1159), .Y(n1161) );
  INVXL U610 ( .A(n1158), .Y(n1160) );
  XNOR2XL U611 ( .A(n1157), .B(n1156), .Y(n1261) );
  NAND2XL U612 ( .A(n859), .B(n1155), .Y(n1157) );
  NAND2XL U613 ( .A(n1167), .B(n1166), .Y(n1169) );
  XOR2XL U614 ( .A(n1145), .B(n1144), .Y(n1257) );
  NAND2XL U615 ( .A(n1143), .B(n1142), .Y(n1144) );
  AOI21XL U616 ( .A0(n1148), .A1(n1147), .B0(n1141), .Y(n1145) );
  NAND2XL U617 ( .A(n994), .B(n993), .Y(n995) );
  INVXL U618 ( .A(n992), .Y(n994) );
  BUFX3 U619 ( .A(A[9]), .Y(n480) );
  OR2X2 U620 ( .A(n951), .B(n950), .Y(n42) );
  OAI21XL U621 ( .A0(n1204), .A1(n1207), .B0(n1205), .Y(n395) );
  AND2X2 U622 ( .A(n534), .B(n220), .Y(n44) );
  XNOR2X2 U623 ( .A(n437), .B(n436), .Y(PRODUCT[29]) );
  OAI22X1 U624 ( .A0(n667), .A1(n512), .B0(n1132), .B1(n479), .Y(n509) );
  OAI22X1 U625 ( .A0(n1041), .A1(n668), .B0(n1042), .B1(n629), .Y(n682) );
  OAI22X1 U626 ( .A0(n446), .A1(n88), .B0(n92), .B1(n997), .Y(n95) );
  OAI22X1 U627 ( .A0(n408), .A1(n997), .B0(n446), .B1(n445), .Y(n60) );
  XNOR2X1 U628 ( .A(n894), .B(B[18]), .Y(n557) );
  OAI22X1 U629 ( .A0(n918), .A1(n338), .B0(n916), .B1(n260), .Y(n309) );
  OAI22X1 U630 ( .A0(n600), .A1(n268), .B0(n923), .B1(n263), .Y(n282) );
  XOR2X1 U631 ( .A(n795), .B(n1230), .Y(PRODUCT[16]) );
  BUFX1 U632 ( .A(n843), .Y(n45) );
  CMPR22X1 U633 ( .A(n707), .B(n706), .CO(n742), .S(n740) );
  OAI22X1 U634 ( .A0(n904), .A1(n811), .B0(n903), .B1(n997), .Y(n901) );
  XNOR2X1 U635 ( .A(n854), .B(B[9]), .Y(n903) );
  OAI22X1 U636 ( .A0(n1134), .A1(n550), .B0(n1132), .B1(n512), .Y(n547) );
  OAI22X1 U637 ( .A0(n1134), .A1(n627), .B0(n1132), .B1(n588), .Y(n624) );
  OAI22X1 U638 ( .A0(n925), .A1(n914), .B0(n923), .B1(n924), .Y(n934) );
  XNOR2X1 U639 ( .A(n1237), .B(n1233), .Y(PRODUCT[14]) );
  XNOR2X2 U640 ( .A(n731), .B(n730), .Y(PRODUCT[21]) );
  OAI21X4 U641 ( .A0(n1220), .A1(n1223), .B0(n1221), .Y(n62) );
  AOI21X4 U642 ( .A0(n62), .A1(n218), .B0(n217), .Y(n651) );
  AOI21X1 U643 ( .A0(n62), .A1(n692), .B0(n691), .Y(n693) );
  AND2X2 U644 ( .A(n533), .B(n220), .Y(n66) );
  OAI21XL U645 ( .A0(n829), .A1(n71), .B0(n828), .Y(n68) );
  XOR3X2 U646 ( .A(n829), .B(n71), .C(n828), .Y(n833) );
  XNOR2X2 U647 ( .A(n854), .B(n630), .Y(n110) );
  OAI21X1 U648 ( .A0(n771), .A1(n694), .B0(n693), .Y(n697) );
  OAI21XL U649 ( .A0(n886), .A1(n1140), .B0(n885), .Y(n986) );
  OAI22X2 U650 ( .A0(n931), .A1(n381), .B0(n929), .B1(n330), .Y(n349) );
  XNOR2X2 U651 ( .A(n920), .B(n1117), .Y(n381) );
  OAI2BB1X1 U652 ( .A0N(n571), .A1N(n43), .B0(n537), .Y(n540) );
  CMPR22X1 U653 ( .A(n113), .B(n112), .CO(n739), .S(n109) );
  OAI21X2 U654 ( .A0(n1216), .A1(n1219), .B0(n1217), .Y(n217) );
  OAI22XL U655 ( .A0(n1041), .A1(n551), .B0(n1042), .B1(n513), .Y(n562) );
  INVX1 U656 ( .A(n224), .Y(n323) );
  OAI22X1 U657 ( .A0(n904), .A1(n147), .B0(n135), .B1(n997), .Y(n175) );
  OAI22X1 U658 ( .A0(n904), .A1(n135), .B0(n88), .B1(n997), .Y(n134) );
  AOI21XL U659 ( .A0(n1074), .A1(n1073), .B0(n1072), .Y(n1109) );
  AOI21XL U660 ( .A0(n1173), .A1(n1172), .B0(n1171), .Y(n1174) );
  AOI21XL U661 ( .A0(n232), .A1(n1170), .B0(n1173), .Y(n1110) );
  OAI22X1 U662 ( .A0(n1041), .A1(n481), .B0(n1042), .B1(n448), .Y(n492) );
  AOI21XL U663 ( .A0(n42), .A1(n978), .B0(n952), .Y(n953) );
  AOI21XL U664 ( .A0(n1156), .A1(n859), .B0(n862), .Y(n1153) );
  XOR2XL U665 ( .A(A[4]), .B(A[5]), .Y(n72) );
  BUFX3 U666 ( .A(n895), .Y(n918) );
  XNOR2X1 U667 ( .A(n894), .B(B[12]), .Y(n102) );
  BUFX3 U668 ( .A(n73), .Y(n916) );
  OAI22XL U669 ( .A0(n918), .A1(n102), .B0(n916), .B1(n82), .Y(n128) );
  XOR2XL U670 ( .A(A[10]), .B(A[11]), .Y(n74) );
  BUFX3 U671 ( .A(n1089), .Y(n1063) );
  BUFX3 U672 ( .A(B[6]), .Y(n893) );
  BUFX3 U673 ( .A(n1090), .Y(n926) );
  OAI22XL U674 ( .A0(n1063), .A1(n103), .B0(n926), .B1(n83), .Y(n127) );
  XOR2XL U675 ( .A(A[6]), .B(A[7]), .Y(n75) );
  XNOR2XL U676 ( .A(A[6]), .B(A[5]), .Y(n76) );
  NAND2X1 U677 ( .A(n75), .B(n76), .Y(n600) );
  BUFX3 U678 ( .A(n600), .Y(n925) );
  BUFX3 U679 ( .A(n76), .Y(n923) );
  XOR2XL U680 ( .A(A[8]), .B(A[9]), .Y(n77) );
  XNOR2XL U681 ( .A(A[8]), .B(A[7]), .Y(n78) );
  NAND2X1 U682 ( .A(n77), .B(n78), .Y(n897) );
  BUFX3 U683 ( .A(n897), .Y(n1041) );
  BUFX3 U684 ( .A(n78), .Y(n1042) );
  XOR2XL U685 ( .A(A[2]), .B(A[3]), .Y(n79) );
  NAND2X1 U686 ( .A(n79), .B(n858), .Y(n591) );
  BUFX3 U687 ( .A(n591), .Y(n931) );
  XNOR2X1 U688 ( .A(n920), .B(B[15]), .Y(n116) );
  BUFX3 U689 ( .A(n858), .Y(n929) );
  BUFX3 U690 ( .A(B[16]), .Y(n596) );
  XOR2XL U691 ( .A(A[12]), .B(A[13]), .Y(n80) );
  BUFX3 U692 ( .A(n1122), .Y(n1094) );
  CLKINVX3 U693 ( .A(n149), .Y(n1092) );
  BUFX3 U694 ( .A(n81), .Y(n1123) );
  OAI22XL U695 ( .A0(n918), .A1(n82), .B0(n916), .B1(n676), .Y(n716) );
  BUFX3 U696 ( .A(B[8]), .Y(n919) );
  NAND2X1 U697 ( .A(A[1]), .B(n85), .Y(n446) );
  XNOR2X1 U698 ( .A(n854), .B(n596), .Y(n92) );
  BUFX3 U699 ( .A(n85), .Y(n997) );
  XOR2XL U700 ( .A(A[14]), .B(A[15]), .Y(n86) );
  NAND2X1 U701 ( .A(n86), .B(n87), .Y(n667) );
  BUFX3 U702 ( .A(n667), .Y(n1134) );
  CLKINVX3 U703 ( .A(n258), .Y(n1130) );
  BUFX3 U704 ( .A(n87), .Y(n1132) );
  XNOR2XL U705 ( .A(n1130), .B(B[2]), .Y(n93) );
  OAI22X1 U706 ( .A0(n1134), .A1(n90), .B0(n1132), .B1(n93), .Y(n94) );
  BUFX3 U707 ( .A(n446), .Y(n904) );
  XNOR2X1 U708 ( .A(n854), .B(B[14]), .Y(n135) );
  OAI22X1 U709 ( .A0(n1134), .A1(n258), .B0(n1132), .B1(n89), .Y(n133) );
  XNOR2X1 U710 ( .A(n480), .B(n893), .Y(n140) );
  XNOR2X1 U711 ( .A(n480), .B(B[7]), .Y(n96) );
  XNOR2XL U712 ( .A(n1130), .B(B[0]), .Y(n91) );
  BUFX8 U713 ( .A(B[17]), .Y(n630) );
  OAI22X1 U714 ( .A0(n446), .A1(n92), .B0(n110), .B1(n997), .Y(n113) );
  OAI22X1 U715 ( .A0(n1134), .A1(n93), .B0(n1132), .B1(n111), .Y(n112) );
  CMPR22X1 U716 ( .A(n95), .B(n94), .CO(n108), .S(n139) );
  OAI22XL U717 ( .A0(n1041), .A1(n96), .B0(n1042), .B1(n115), .Y(n101) );
  XNOR2X1 U718 ( .A(n920), .B(B[13]), .Y(n98) );
  XNOR2X1 U719 ( .A(n920), .B(B[14]), .Y(n117) );
  OAI22XL U720 ( .A0(n931), .A1(n98), .B0(n929), .B1(n117), .Y(n100) );
  OAI22XL U721 ( .A0(n931), .A1(n141), .B0(n929), .B1(n98), .Y(n170) );
  CMPR32X1 U722 ( .A(n101), .B(n100), .C(n99), .CO(n107), .S(n204) );
  XNOR2X1 U723 ( .A(n894), .B(n628), .Y(n132) );
  OAI22XL U724 ( .A0(n918), .A1(n132), .B0(n916), .B1(n102), .Y(n122) );
  OAI22XL U725 ( .A0(n1063), .A1(n104), .B0(n926), .B1(n103), .Y(n121) );
  OAI22X1 U726 ( .A0(n904), .A1(n110), .B0(n664), .B1(n997), .Y(n707) );
  OAI22X1 U727 ( .A0(n1134), .A1(n111), .B0(n1132), .B1(n666), .Y(n706) );
  CMPR32X1 U728 ( .A(n122), .B(n121), .C(n120), .CO(n131), .S(n203) );
  CMPR32X1 U729 ( .A(n125), .B(n124), .C(n123), .CO(n738), .S(n130) );
  CMPR32X1 U730 ( .A(n128), .B(n127), .C(n126), .CO(n746), .S(n129) );
  CMPR32X1 U731 ( .A(n131), .B(n130), .C(n129), .CO(n761), .S(n785) );
  OAI22XL U732 ( .A0(n918), .A1(n145), .B0(n916), .B1(n132), .Y(n173) );
  CMPR22X1 U733 ( .A(n134), .B(n133), .CO(n138), .S(n172) );
  XNOR2X1 U734 ( .A(n854), .B(B[13]), .Y(n147) );
  CMPR32X1 U735 ( .A(n139), .B(n138), .C(n137), .CO(n152), .S(n210) );
  XNOR2X1 U736 ( .A(n920), .B(n628), .Y(n178) );
  OAI22XL U737 ( .A0(n931), .A1(n178), .B0(n929), .B1(n141), .Y(n182) );
  CMPR32X1 U738 ( .A(n144), .B(n143), .C(n142), .CO(n137), .S(n154) );
  NOR2X1 U739 ( .A(n790), .B(n789), .Y(mult_x_1_n299) );
  CMPR32X1 U740 ( .A(n155), .B(n154), .C(n153), .CO(n209), .S(n214) );
  XNOR2X1 U741 ( .A(n913), .B(n893), .Y(n167) );
  XNOR2XL U742 ( .A(n1092), .B(B[0]), .Y(n158) );
  XNOR2XL U743 ( .A(n1043), .B(B[2]), .Y(n166) );
  ADDHXL U744 ( .A(n164), .B(n163), .CO(n160), .S(n1000) );
  XNOR2X1 U745 ( .A(n920), .B(B[9]), .Y(n928) );
  XNOR2X1 U746 ( .A(n920), .B(B[10]), .Y(n179) );
  CMPR32X1 U747 ( .A(n170), .B(n169), .C(n168), .CO(n205), .S(n208) );
  CMPR32X1 U748 ( .A(n173), .B(n172), .C(n171), .CO(n211), .S(n207) );
  OAI22XL U749 ( .A0(n1041), .A1(n194), .B0(n1042), .B1(n177), .Y(n193) );
  OAI22X1 U750 ( .A0(n931), .A1(n179), .B0(n929), .B1(n178), .Y(n192) );
  OAI22XL U751 ( .A0(n895), .A1(n181), .B0(n916), .B1(n180), .Y(n191) );
  CMPR32X1 U752 ( .A(n187), .B(n186), .C(n185), .CO(n206), .S(n1012) );
  CMPR32X1 U753 ( .A(n190), .B(n189), .C(n188), .CO(n202), .S(n1006) );
  OAI22X1 U754 ( .A0(n1063), .A1(n196), .B0(n926), .B1(n195), .Y(n898) );
  ADDFHX1 U755 ( .A(n199), .B(n198), .CI(n197), .CO(n999), .S(n955) );
  NAND2XL U756 ( .A(n797), .B(n796), .Y(mult_x_1_n313) );
  CMPR32X1 U757 ( .A(n205), .B(n204), .C(n203), .CO(n150), .S(n788) );
  CMPR32X1 U758 ( .A(n214), .B(n213), .C(n212), .CO(n215), .S(n797) );
  OAI21XL U759 ( .A0(n798), .A1(mult_x_1_n313), .B0(n799), .Y(mult_x_1_n306)
         );
  NOR2X1 U760 ( .A(n1214), .B(n1212), .Y(n533) );
  NOR2X1 U761 ( .A(n1210), .B(n1208), .Y(n220) );
  OAI21X1 U762 ( .A0(n1212), .A1(n1215), .B0(n1213), .Y(n534) );
  NAND2XL U763 ( .A(n255), .B(n247), .Y(n227) );
  NOR2XL U764 ( .A(n1194), .B(n227), .Y(n229) );
  INVXL U765 ( .A(n221), .Y(n234) );
  OAI21XL U766 ( .A0(n1200), .A1(n1203), .B0(n1201), .Y(n222) );
  OAI21XL U767 ( .A0(n1196), .A1(n1199), .B0(n1197), .Y(n293) );
  OAI21XL U768 ( .A0(n227), .A1(n1195), .B0(n226), .Y(n228) );
  AOI21XL U769 ( .A0(n293), .A1(n229), .B0(n228), .Y(n230) );
  OAI21XL U770 ( .A0(n1179), .A1(n234), .B0(n233), .Y(n236) );
  INVXL U771 ( .A(n238), .Y(n292) );
  INVXL U772 ( .A(n1194), .Y(n296) );
  NAND2XL U773 ( .A(n296), .B(n255), .Y(n242) );
  NOR2XL U774 ( .A(n292), .B(n242), .Y(n244) );
  NAND2XL U775 ( .A(n362), .B(n244), .Y(n246) );
  AOI21XL U776 ( .A0(n240), .A1(n255), .B0(n239), .Y(n241) );
  OAI21XL U777 ( .A0(n250), .A1(n242), .B0(n241), .Y(n243) );
  AOI21XL U778 ( .A0(n323), .A1(n244), .B0(n243), .Y(n245) );
  OAI21XL U779 ( .A0(n1179), .A1(n246), .B0(n245), .Y(n249) );
  NOR2XL U780 ( .A(n292), .B(n1194), .Y(n252) );
  NAND2XL U781 ( .A(n362), .B(n252), .Y(n254) );
  OAI21XL U782 ( .A0(n250), .A1(n1194), .B0(n1195), .Y(n251) );
  AOI21XL U783 ( .A0(n323), .A1(n252), .B0(n251), .Y(n253) );
  XNOR2X2 U784 ( .A(n257), .B(n256), .Y(PRODUCT[34]) );
  INVXL U785 ( .A(n894), .Y(n838) );
  BUFX3 U786 ( .A(B[25]), .Y(n1117) );
  XNOR2X1 U787 ( .A(n894), .B(n1117), .Y(n338) );
  BUFX3 U788 ( .A(B[26]), .Y(n1129) );
  XNOR2X1 U789 ( .A(A[13]), .B(B[19]), .Y(n269) );
  OAI22XL U790 ( .A0(n1041), .A1(n299), .B0(n1042), .B1(n267), .Y(n272) );
  XNOR2X1 U791 ( .A(n913), .B(n1117), .Y(n268) );
  INVXL U792 ( .A(n282), .Y(n271) );
  XNOR2X1 U793 ( .A(A[13]), .B(B[21]), .Y(n277) );
  OAI22XL U794 ( .A0(n1089), .A1(n266), .B0(n1090), .B1(n280), .Y(n285) );
  XNOR2X1 U795 ( .A(n913), .B(B[24]), .Y(n301) );
  XNOR2X1 U796 ( .A(A[13]), .B(B[18]), .Y(n303) );
  CMPR32X1 U797 ( .A(n273), .B(n272), .C(n271), .CO(n289), .S(n315) );
  CMPR32X1 U798 ( .A(n276), .B(n275), .C(n274), .CO(n319), .S(n314) );
  XNOR2X1 U799 ( .A(A[13]), .B(B[22]), .Y(n1045) );
  OAI22X1 U800 ( .A0(n1041), .A1(n279), .B0(n1042), .B1(n1039), .Y(n1058) );
  CMPR32X1 U801 ( .A(n283), .B(n282), .C(n281), .CO(n1050), .S(n288) );
  CMPR32X1 U802 ( .A(n286), .B(n285), .C(n284), .CO(n1049), .S(n287) );
  CMPR32X1 U803 ( .A(n289), .B(n288), .C(n287), .CO(n1035), .S(n318) );
  NOR2XL U804 ( .A(n291), .B(n290), .Y(mult_x_1_n162) );
  NAND2XL U805 ( .A(n291), .B(n290), .Y(mult_x_1_n163) );
  NAND2XL U806 ( .A(n362), .B(n238), .Y(n295) );
  AOI21XL U807 ( .A0(n323), .A1(n238), .B0(n293), .Y(n294) );
  NAND2X1 U808 ( .A(n296), .B(n1195), .Y(n297) );
  XNOR2X2 U809 ( .A(n298), .B(n297), .Y(PRODUCT[33]) );
  OAI22XL U810 ( .A0(n1089), .A1(n342), .B0(n1090), .B1(n300), .Y(n337) );
  XNOR2X1 U811 ( .A(n913), .B(B[23]), .Y(n340) );
  INVXL U812 ( .A(n309), .Y(n335) );
  XNOR2X1 U813 ( .A(n1118), .B(B[15]), .Y(n329) );
  OAI22XL U814 ( .A0(n1134), .A1(n329), .B0(n1132), .B1(n302), .Y(n334) );
  XNOR2X1 U815 ( .A(A[13]), .B(n630), .Y(n339) );
  OAI22XL U816 ( .A0(n1122), .A1(n339), .B0(n1123), .B1(n303), .Y(n333) );
  CMPR32X1 U817 ( .A(n307), .B(n306), .C(n305), .CO(n316), .S(n356) );
  CMPR32X1 U818 ( .A(n310), .B(n309), .C(n308), .CO(n274), .S(n355) );
  ADDFHX1 U819 ( .A(n313), .B(n312), .CI(n311), .CO(n359), .S(n354) );
  CMPR32X1 U820 ( .A(n319), .B(n318), .C(n317), .CO(n291), .S(n320) );
  NOR2XL U821 ( .A(n321), .B(n320), .Y(mult_x_1_n173) );
  NAND2XL U822 ( .A(n321), .B(n320), .Y(mult_x_1_n174) );
  NAND2XL U823 ( .A(n362), .B(n363), .Y(n325) );
  INVXL U824 ( .A(n1196), .Y(n326) );
  NAND2X1 U825 ( .A(n326), .B(n1197), .Y(n327) );
  XNOR2X4 U826 ( .A(n328), .B(n327), .Y(PRODUCT[32]) );
  OAI22XL U827 ( .A0(n1134), .A1(n346), .B0(n1132), .B1(n329), .Y(n350) );
  XNOR2X1 U828 ( .A(n920), .B(n1129), .Y(n330) );
  INVXL U829 ( .A(n330), .Y(n331) );
  CMPR32X1 U830 ( .A(n334), .B(n333), .C(n332), .CO(n311), .S(n370) );
  CMPR32X1 U831 ( .A(n337), .B(n336), .C(n335), .CO(n312), .S(n369) );
  OAI22XL U832 ( .A0(n918), .A1(n344), .B0(n916), .B1(n338), .Y(n353) );
  OAI22XL U833 ( .A0(n1094), .A1(n372), .B0(n1123), .B1(n339), .Y(n352) );
  XNOR2X1 U834 ( .A(n913), .B(B[22]), .Y(n345) );
  OAI22XL U835 ( .A0(n1041), .A1(n347), .B0(n1042), .B1(n341), .Y(n380) );
  XNOR2X1 U836 ( .A(n1043), .B(B[18]), .Y(n343) );
  OAI22XL U837 ( .A0(n1089), .A1(n343), .B0(n1090), .B1(n342), .Y(n379) );
  XNOR2X1 U838 ( .A(n1043), .B(n630), .Y(n382) );
  OAI22X1 U839 ( .A0(n1063), .A1(n382), .B0(n926), .B1(n343), .Y(n386) );
  OAI22X1 U840 ( .A0(n918), .A1(n383), .B0(n916), .B1(n344), .Y(n385) );
  INVXL U841 ( .A(n349), .Y(n384) );
  XNOR2X1 U842 ( .A(n1130), .B(B[13]), .Y(n376) );
  XNOR2X1 U843 ( .A(n480), .B(B[19]), .Y(n375) );
  ADDFHX1 U844 ( .A(n350), .B(n349), .CI(n348), .CO(n371), .S(n406) );
  CMPR32X1 U845 ( .A(n353), .B(n352), .C(n351), .CO(n392), .S(n405) );
  CMPR32X1 U846 ( .A(n356), .B(n355), .C(n354), .CO(n358), .S(n366) );
  CMPR32X1 U847 ( .A(n359), .B(n358), .C(n357), .CO(n321), .S(n360) );
  NOR2XL U848 ( .A(n361), .B(n360), .Y(mult_x_1_n184) );
  NAND2XL U849 ( .A(n361), .B(n360), .Y(mult_x_1_n185) );
  NAND2X1 U850 ( .A(n363), .B(n1199), .Y(n364) );
  XNOR2X2 U851 ( .A(n365), .B(n364), .Y(PRODUCT[31]) );
  CMPR32X1 U852 ( .A(n368), .B(n367), .C(n366), .CO(n361), .S(n394) );
  CMPR32X1 U853 ( .A(n371), .B(n370), .C(n369), .CO(n368), .S(n404) );
  XNOR2X1 U854 ( .A(A[13]), .B(B[15]), .Y(n374) );
  OAI22XL U855 ( .A0(n1094), .A1(n414), .B0(n1123), .B1(n374), .Y(n410) );
  XNOR2X1 U856 ( .A(n854), .B(n1129), .Y(n408) );
  INVXL U857 ( .A(n408), .Y(n377) );
  CMPR32X1 U858 ( .A(n380), .B(n379), .C(n378), .CO(n391), .S(n428) );
  XNOR2X1 U859 ( .A(n920), .B(B[24]), .Y(n413) );
  XNOR2X1 U860 ( .A(n1043), .B(n596), .Y(n419) );
  XNOR2X1 U861 ( .A(n894), .B(B[22]), .Y(n418) );
  OAI22XL U862 ( .A0(n918), .A1(n418), .B0(n916), .B1(n383), .Y(n424) );
  NOR2XL U863 ( .A(n394), .B(n393), .Y(mult_x_1_n191) );
  NAND2XL U864 ( .A(n394), .B(n393), .Y(mult_x_1_n192) );
  INVXL U865 ( .A(n1203), .Y(n396) );
  AOI21XL U866 ( .A0(n395), .A1(n435), .B0(n396), .Y(n397) );
  CMPR32X1 U867 ( .A(n404), .B(n403), .C(n402), .CO(n393), .S(n431) );
  CMPR32X1 U868 ( .A(n407), .B(n406), .C(n405), .CO(n390), .S(n440) );
  XNOR2X1 U869 ( .A(n1130), .B(n628), .Y(n447) );
  OAI22XL U870 ( .A0(n1134), .A1(n447), .B0(n1132), .B1(n409), .Y(n444) );
  XNOR2X1 U871 ( .A(n411), .B(n410), .Y(n452) );
  OAI22X1 U872 ( .A0(n1041), .A1(n448), .B0(n1042), .B1(n412), .Y(n459) );
  XNOR2X1 U873 ( .A(n920), .B(B[23]), .Y(n449) );
  OAI22X1 U874 ( .A0(n931), .A1(n449), .B0(n858), .B1(n413), .Y(n458) );
  CMPR32X1 U875 ( .A(n417), .B(n416), .C(n415), .CO(n429), .S(n464) );
  XNOR2X1 U876 ( .A(n894), .B(B[21]), .Y(n454) );
  OAI22X1 U877 ( .A0(n918), .A1(n454), .B0(n916), .B1(n418), .Y(n462) );
  XNOR2X1 U878 ( .A(n1043), .B(B[15]), .Y(n455) );
  OAI22XL U879 ( .A0(n1063), .A1(n455), .B0(n926), .B1(n419), .Y(n461) );
  NOR2XL U880 ( .A(n431), .B(n430), .Y(mult_x_1_n202) );
  NAND2XL U881 ( .A(n431), .B(n430), .Y(mult_x_1_n203) );
  INVXL U882 ( .A(n432), .Y(n434) );
  CMPR32X1 U883 ( .A(n440), .B(n439), .C(n438), .CO(n430), .S(n467) );
  OAI22XL U884 ( .A0(n667), .A1(n479), .B0(n1132), .B1(n447), .Y(n476) );
  XNOR2X1 U885 ( .A(n480), .B(n596), .Y(n481) );
  XNOR2X1 U886 ( .A(n920), .B(B[22]), .Y(n482) );
  OAI22X1 U887 ( .A0(n931), .A1(n482), .B0(n929), .B1(n449), .Y(n491) );
  CMPR32X1 U888 ( .A(n453), .B(n452), .C(n451), .CO(n465), .S(n497) );
  XNOR2X1 U889 ( .A(n894), .B(B[20]), .Y(n487) );
  OAI22XL U890 ( .A0(n1063), .A1(n488), .B0(n926), .B1(n455), .Y(n494) );
  CMPR32X1 U891 ( .A(n462), .B(n461), .C(n460), .CO(n475), .S(n506) );
  NOR2XL U892 ( .A(n467), .B(n466), .Y(mult_x_1_n209) );
  NAND2XL U893 ( .A(n467), .B(n466), .Y(mult_x_1_n210) );
  CMPR32X1 U894 ( .A(n475), .B(n474), .C(n473), .CO(n463), .S(n505) );
  ADDHXL U895 ( .A(n477), .B(n476), .CO(n485), .S(n518) );
  XNOR2X1 U896 ( .A(n854), .B(B[23]), .Y(n511) );
  OAI22XL U897 ( .A0(n1041), .A1(n513), .B0(n1042), .B1(n481), .Y(n524) );
  XNOR2X1 U898 ( .A(n920), .B(B[21]), .Y(n514) );
  OAI22X1 U899 ( .A0(n591), .A1(n514), .B0(n929), .B1(n482), .Y(n523) );
  XNOR2X1 U900 ( .A(n894), .B(B[19]), .Y(n519) );
  XNOR2X1 U901 ( .A(n1043), .B(B[13]), .Y(n520) );
  OAI22XL U902 ( .A0(n600), .A1(n521), .B0(n923), .B1(n489), .Y(n525) );
  CMPR32X1 U903 ( .A(n495), .B(n494), .C(n493), .CO(n508), .S(n544) );
  INVXL U904 ( .A(n1206), .Y(n501) );
  NAND2X1 U905 ( .A(n501), .B(n1207), .Y(n502) );
  CMPR32X1 U906 ( .A(n508), .B(n507), .C(n506), .CO(n496), .S(n543) );
  CMPR22X1 U907 ( .A(n510), .B(n509), .CO(n517), .S(n556) );
  OAI22X1 U908 ( .A0(n904), .A1(n549), .B0(n511), .B1(n997), .Y(n548) );
  XNOR2X1 U909 ( .A(n920), .B(B[20]), .Y(n552) );
  OAI22X1 U910 ( .A0(n591), .A1(n552), .B0(n929), .B1(n514), .Y(n561) );
  XNOR2X1 U911 ( .A(n1043), .B(B[12]), .Y(n558) );
  OAI22XL U912 ( .A0(n600), .A1(n559), .B0(n923), .B1(n521), .Y(n563) );
  ADDFHX1 U913 ( .A(n524), .B(n523), .CI(n522), .CO(n516), .S(n584) );
  CMPR32X1 U914 ( .A(n530), .B(n529), .C(n528), .CO(n504), .S(n541) );
  NOR2XL U915 ( .A(n532), .B(n531), .Y(mult_x_1_n223) );
  INVXL U916 ( .A(n533), .Y(n572) );
  NOR2XL U917 ( .A(n572), .B(n1210), .Y(n536) );
  CLKINVX3 U918 ( .A(n651), .Y(n573) );
  INVXL U919 ( .A(n534), .Y(n574) );
  OAI21XL U920 ( .A0(n574), .A1(n1210), .B0(n1211), .Y(n535) );
  NAND2X1 U921 ( .A(n538), .B(n1209), .Y(n539) );
  CMPR32X1 U922 ( .A(n543), .B(n542), .C(n541), .CO(n531), .S(n570) );
  CMPR32X1 U923 ( .A(n546), .B(n545), .C(n544), .CO(n528), .S(n582) );
  CMPR22X1 U924 ( .A(n548), .B(n547), .CO(n555), .S(n595) );
  XNOR2X1 U925 ( .A(n480), .B(B[13]), .Y(n589) );
  OAI22XL U926 ( .A0(n897), .A1(n589), .B0(n1042), .B1(n551), .Y(n603) );
  XNOR2X1 U927 ( .A(n920), .B(B[19]), .Y(n590) );
  OAI22X1 U928 ( .A0(n931), .A1(n590), .B0(n929), .B1(n552), .Y(n602) );
  ADDFHX1 U929 ( .A(n562), .B(n561), .CI(n560), .CO(n554), .S(n622) );
  NOR2XL U930 ( .A(n570), .B(n569), .Y(mult_x_1_n232) );
  NAND2XL U931 ( .A(n570), .B(n569), .Y(mult_x_1_n233) );
  NAND2XL U932 ( .A(n650), .B(n533), .Y(n576) );
  CMPR32X1 U933 ( .A(n585), .B(n584), .C(n583), .CO(n566), .S(n620) );
  XNOR2X1 U934 ( .A(n854), .B(B[20]), .Y(n626) );
  OAI22X1 U935 ( .A0(n904), .A1(n626), .B0(n587), .B1(n997), .Y(n625) );
  XNOR2X1 U936 ( .A(n480), .B(B[12]), .Y(n629) );
  OAI22XL U937 ( .A0(n1041), .A1(n629), .B0(n1042), .B1(n589), .Y(n641) );
  XNOR2X1 U938 ( .A(n920), .B(B[18]), .Y(n631) );
  OAI22X1 U939 ( .A0(n591), .A1(n631), .B0(n929), .B1(n590), .Y(n640) );
  XNOR2X1 U940 ( .A(n894), .B(n596), .Y(n636) );
  NAND2XL U941 ( .A(n611), .B(n610), .Y(mult_x_1_n242) );
  INVX1 U942 ( .A(n1214), .Y(n613) );
  NAND2XL U943 ( .A(n650), .B(n613), .Y(n615) );
  CMPR32X1 U944 ( .A(n623), .B(n622), .C(n621), .CO(n607), .S(n657) );
  CMPR22X1 U945 ( .A(n625), .B(n624), .CO(n634), .S(n674) );
  XNOR2X1 U946 ( .A(n854), .B(B[19]), .Y(n663) );
  OAI22X1 U947 ( .A0(n904), .A1(n663), .B0(n626), .B1(n997), .Y(n662) );
  OAI22X1 U948 ( .A0(n1134), .A1(n665), .B0(n1132), .B1(n627), .Y(n661) );
  XNOR2X1 U949 ( .A(n480), .B(n628), .Y(n668) );
  XNOR2X1 U950 ( .A(n894), .B(B[15]), .Y(n675) );
  OAI22XL U951 ( .A0(n918), .A1(n675), .B0(n916), .B1(n636), .Y(n685) );
  CMPR32X1 U952 ( .A(n641), .B(n640), .C(n639), .CO(n633), .S(n702) );
  NOR2XL U953 ( .A(n649), .B(n648), .Y(mult_x_1_n252) );
  NAND2XL U954 ( .A(n649), .B(n648), .Y(mult_x_1_n253) );
  INVXL U955 ( .A(n650), .Y(n652) );
  CMPR32X1 U956 ( .A(n657), .B(n656), .C(n655), .CO(n648), .S(n690) );
  CMPR22X1 U957 ( .A(n662), .B(n661), .CO(n673), .S(n713) );
  OAI22X1 U958 ( .A0(n904), .A1(n664), .B0(n663), .B1(n997), .Y(n705) );
  OAI22X1 U959 ( .A0(n667), .A1(n666), .B0(n1132), .B1(n665), .Y(n704) );
  OAI22XL U960 ( .A0(n918), .A1(n676), .B0(n916), .B1(n675), .Y(n722) );
  CMPR32X1 U961 ( .A(n685), .B(n684), .C(n683), .CO(n703), .S(n735) );
  NAND2XL U962 ( .A(n690), .B(n689), .Y(mult_x_1_n260) );
  NAND2XL U963 ( .A(n728), .B(n692), .Y(n694) );
  INVXL U964 ( .A(n1216), .Y(n695) );
  XNOR2X2 U965 ( .A(n697), .B(n696), .Y(PRODUCT[22]) );
  CMPR32X1 U966 ( .A(n700), .B(n699), .C(n698), .CO(n689), .S(n727) );
  CMPR32X1 U967 ( .A(n703), .B(n702), .C(n701), .CO(n686), .S(n734) );
  CMPR22X1 U968 ( .A(n705), .B(n704), .CO(n712), .S(n743) );
  CMPR32X1 U969 ( .A(n710), .B(n709), .C(n708), .CO(n741), .S(n745) );
  CMPR32X1 U970 ( .A(n716), .B(n715), .C(n714), .CO(n760), .S(n744) );
  CMPR32X1 U971 ( .A(n722), .B(n721), .C(n720), .CO(n737), .S(n758) );
  CMPR32X1 U972 ( .A(n725), .B(n724), .C(n723), .CO(n699), .S(n732) );
  NOR2XL U973 ( .A(n727), .B(n726), .Y(mult_x_1_n270) );
  NAND2XL U974 ( .A(n727), .B(n726), .Y(mult_x_1_n271) );
  CMPR32X1 U975 ( .A(n740), .B(n739), .C(n738), .CO(n766), .S(n762) );
  CMPR32X1 U976 ( .A(n743), .B(n742), .C(n741), .CO(n749), .S(n765) );
  CMPR32X1 U977 ( .A(n746), .B(n745), .C(n744), .CO(n764), .S(n777) );
  CMPR32X1 U978 ( .A(n749), .B(n748), .C(n747), .CO(n733), .S(n755) );
  NOR2XL U979 ( .A(n751), .B(n750), .Y(mult_x_1_n277) );
  NAND2XL U980 ( .A(n751), .B(n750), .Y(mult_x_1_n278) );
  INVXL U981 ( .A(n1220), .Y(n752) );
  NAND2X1 U982 ( .A(n752), .B(n1221), .Y(n753) );
  CMPR32X1 U983 ( .A(n757), .B(n756), .C(n755), .CO(n750), .S(n768) );
  CMPR32X1 U984 ( .A(n763), .B(n762), .C(n761), .CO(n773), .S(n775) );
  NOR2XL U985 ( .A(n768), .B(n767), .Y(mult_x_1_n288) );
  NAND2XL U986 ( .A(n768), .B(n767), .Y(mult_x_1_n289) );
  INVXL U987 ( .A(n1222), .Y(n769) );
  CMPR32X1 U988 ( .A(n774), .B(n773), .C(n772), .CO(n767), .S(n779) );
  NOR2XL U989 ( .A(n779), .B(n778), .Y(mult_x_1_n291) );
  NAND2XL U990 ( .A(n779), .B(n778), .Y(mult_x_1_n292) );
  OAI21XL U991 ( .A0(n791), .A1(n1227), .B0(n1228), .Y(n782) );
  INVXL U992 ( .A(n1225), .Y(n780) );
  XNOR2X2 U993 ( .A(n782), .B(n781), .Y(PRODUCT[18]) );
  CMPR32X1 U994 ( .A(n785), .B(n784), .C(n783), .CO(n789), .S(n793) );
  NOR2XL U995 ( .A(mult_x_1_n302), .B(mult_x_1_n299), .Y(mult_x_1_n297) );
  NAND2XL U996 ( .A(n790), .B(n789), .Y(mult_x_1_n300) );
  NAND2XL U997 ( .A(n793), .B(n792), .Y(mult_x_1_n303) );
  INVX1 U998 ( .A(n1231), .Y(n801) );
  INVXL U999 ( .A(n1232), .Y(n794) );
  AOI21X1 U1000 ( .A0(n803), .A1(n801), .B0(n794), .Y(n795) );
  NOR2XL U1001 ( .A(n798), .B(mult_x_1_n312), .Y(mult_x_1_n305) );
  INVXL U1002 ( .A(n798), .Y(n800) );
  NAND2XL U1003 ( .A(n800), .B(n799), .Y(mult_x_1_n78) );
  XNOR2X1 U1004 ( .A(n803), .B(n802), .Y(PRODUCT[15]) );
  OAI22XL U1005 ( .A0(n925), .A1(n813), .B0(n923), .B1(n914), .Y(n909) );
  XNOR2XL U1006 ( .A(n480), .B(B[0]), .Y(n804) );
  OAI22XL U1007 ( .A0(n1041), .A1(n804), .B0(n1042), .B1(n906), .Y(n908) );
  XNOR2X1 U1008 ( .A(n920), .B(n893), .Y(n808) );
  XNOR2X1 U1009 ( .A(n894), .B(B[3]), .Y(n819) );
  OAI22XL U1010 ( .A0(n895), .A1(n819), .B0(n916), .B1(n805), .Y(n821) );
  XNOR2X1 U1011 ( .A(n854), .B(B[7]), .Y(n812) );
  OAI22XL U1012 ( .A0(n904), .A1(n830), .B0(n812), .B1(n997), .Y(n827) );
  OAI22XL U1013 ( .A0(n931), .A1(n808), .B0(n929), .B1(n921), .Y(n937) );
  OAI22X1 U1014 ( .A0(n1041), .A1(n810), .B0(n1042), .B1(n809), .Y(n900) );
  OAI22X1 U1015 ( .A0(n904), .A1(n812), .B0(n811), .B1(n997), .Y(n815) );
  CMPR32X1 U1016 ( .A(n816), .B(n815), .C(n814), .CO(n935), .S(n825) );
  XNOR2XL U1017 ( .A(n913), .B(B[0]), .Y(n818) );
  OAI22X1 U1018 ( .A0(n925), .A1(n818), .B0(n923), .B1(n817), .Y(n829) );
  XNOR2XL U1019 ( .A(n894), .B(B[2]), .Y(n831) );
  OAI22X1 U1020 ( .A0(n918), .A1(n831), .B0(n916), .B1(n819), .Y(n828) );
  CMPR32X1 U1021 ( .A(n822), .B(n821), .C(n820), .CO(n945), .S(n823) );
  ADDHXL U1022 ( .A(n827), .B(n826), .CO(n820), .S(n834) );
  XNOR2XL U1023 ( .A(n894), .B(B[1]), .Y(n846) );
  NOR2XL U1024 ( .A(n987), .B(n992), .Y(n892) );
  XNOR2XL U1025 ( .A(n920), .B(B[3]), .Y(n845) );
  OAI22XL U1026 ( .A0(n904), .A1(n863), .B0(n836), .B1(n997), .Y(n849) );
  CMPR32X1 U1027 ( .A(n841), .B(n840), .C(n839), .CO(n832), .S(n842) );
  XNOR2XL U1028 ( .A(n920), .B(B[2]), .Y(n865) );
  XNOR2XL U1029 ( .A(n894), .B(B[0]), .Y(n847) );
  ADDHXL U1030 ( .A(n849), .B(n848), .CO(n843), .S(n871) );
  OR2X2 U1031 ( .A(n881), .B(n880), .Y(n1147) );
  XNOR2XL U1032 ( .A(n854), .B(B[1]), .Y(n850) );
  XNOR2XL U1033 ( .A(n854), .B(B[2]), .Y(n855) );
  OAI21XL U1034 ( .A0(n1158), .A1(n1164), .B0(n1159), .Y(n1156) );
  XNOR2XL U1035 ( .A(n854), .B(B[3]), .Y(n864) );
  OAI22X1 U1036 ( .A0(n904), .A1(n855), .B0(n864), .B1(n997), .Y(n868) );
  XNOR2XL U1037 ( .A(n920), .B(B[0]), .Y(n856) );
  XNOR2XL U1038 ( .A(n920), .B(B[1]), .Y(n866) );
  OAI22X1 U1039 ( .A0(n931), .A1(n856), .B0(n929), .B1(n866), .Y(n867) );
  CMPR22X1 U1040 ( .A(n868), .B(n867), .CO(n869), .S(n861) );
  OAI21XL U1041 ( .A0(n1153), .A1(n1150), .B0(n1151), .Y(n1168) );
  CMPR32X1 U1042 ( .A(n873), .B(n872), .C(n871), .CO(n880), .S(n878) );
  CMPR32X1 U1043 ( .A(n876), .B(n875), .C(n874), .CO(n877), .S(n870) );
  OR2X2 U1044 ( .A(n878), .B(n877), .Y(n1167) );
  NAND2XL U1045 ( .A(n881), .B(n880), .Y(n1146) );
  INVXL U1046 ( .A(n1146), .Y(n1141) );
  NAND2XL U1047 ( .A(n883), .B(n882), .Y(n1142) );
  INVXL U1048 ( .A(n1142), .Y(n884) );
  NAND2XL U1049 ( .A(n890), .B(n889), .Y(n988) );
  OAI21XL U1050 ( .A0(n987), .A1(n993), .B0(n988), .Y(n891) );
  XNOR2X1 U1051 ( .A(n894), .B(n893), .Y(n915) );
  OAI22X1 U1052 ( .A0(n897), .A1(n905), .B0(n1042), .B1(n896), .Y(n965) );
  CMPR22X1 U1053 ( .A(n899), .B(n898), .CO(n956), .S(n964) );
  CMPR22X1 U1054 ( .A(n901), .B(n900), .CO(n940), .S(n936) );
  ADDFHX1 U1055 ( .A(n912), .B(n911), .CI(n910), .CO(n960), .S(n939) );
  OAI22X2 U1056 ( .A0(n918), .A1(n917), .B0(n916), .B1(n915), .Y(n933) );
  OAI22XL U1057 ( .A0(n931), .A1(n921), .B0(n929), .B1(n930), .Y(n932) );
  OAI22XL U1058 ( .A0(n925), .A1(n924), .B0(n923), .B1(n922), .Y(n963) );
  XNOR2XL U1059 ( .A(n1043), .B(B[0]), .Y(n927) );
  OAI22XL U1060 ( .A0(n931), .A1(n930), .B0(n929), .B1(n928), .Y(n961) );
  CMPR32X1 U1061 ( .A(n937), .B(n936), .C(n935), .CO(n942), .S(n944) );
  CMPR32X1 U1062 ( .A(n946), .B(n945), .C(n944), .CO(n948), .S(n890) );
  NOR2XL U1063 ( .A(n949), .B(n948), .Y(n947) );
  NAND2XL U1064 ( .A(n42), .B(n983), .Y(n954) );
  INVXL U1065 ( .A(n982), .Y(n978) );
  NAND2XL U1066 ( .A(n951), .B(n950), .Y(n979) );
  INVXL U1067 ( .A(n979), .Y(n952) );
  OAI21XL U1068 ( .A0(n977), .A1(n954), .B0(n953), .Y(n1022) );
  CMPR32X1 U1069 ( .A(n957), .B(n956), .C(n955), .CO(n1004), .S(n1009) );
  CMPR32X1 U1070 ( .A(n963), .B(n962), .C(n961), .CO(n1003), .S(n958) );
  ADDFHX1 U1071 ( .A(n966), .B(n965), .CI(n964), .CO(n1002), .S(n972) );
  CMPR32X1 U1072 ( .A(n969), .B(n968), .C(n967), .CO(n998), .S(n1001) );
  XOR2X1 U1073 ( .A(n1027), .B(n976), .Y(n1252) );
  NAND2XL U1074 ( .A(n42), .B(n979), .Y(n980) );
  NAND2XL U1075 ( .A(n983), .B(n982), .Y(n984) );
  OAI21XL U1076 ( .A0(n996), .A1(n992), .B0(n993), .Y(n991) );
  INVXL U1077 ( .A(n987), .Y(n989) );
  CMPR32X1 U1078 ( .A(n998), .B(n999), .C(n1000), .CO(n200), .S(n1015) );
  CMPR32X1 U1079 ( .A(n1003), .B(n1002), .C(n1001), .CO(n1014), .S(n1007) );
  CMPR32X1 U1080 ( .A(n1006), .B(n1005), .C(n1004), .CO(n1011), .S(n1013) );
  CMPR32X1 U1081 ( .A(n1009), .B(n1008), .C(n1007), .CO(n1017), .S(n975) );
  NAND2XL U1082 ( .A(n1070), .B(n1026), .Y(n1025) );
  NOR2XL U1083 ( .A(n1025), .B(n1032), .Y(n1023) );
  OAI21XL U1084 ( .A0(n1024), .A1(n1032), .B0(n1033), .Y(n1021) );
  AOI21XL U1085 ( .A0(n1023), .A1(n1022), .B0(n1021), .Y(mult_x_1_n315) );
  OAI21XL U1086 ( .A0(n1027), .A1(n973), .B0(n1016), .Y(mult_x_1_n327) );
  OAI21XL U1087 ( .A0(n1179), .A1(n1029), .B0(n1028), .Y(n1031) );
  XNOR2X1 U1088 ( .A(n1118), .B(B[21]), .Y(n1061) );
  CMPR32X1 U1089 ( .A(n1048), .B(n1047), .C(n1046), .CO(n1064), .S(n1037) );
  CMPR32X1 U1090 ( .A(n1051), .B(n1050), .C(n1049), .CO(n1054), .S(n1036) );
  CMPR32X1 U1091 ( .A(n1059), .B(n1058), .C(n1057), .CO(n1102), .S(n1056) );
  XNOR2X1 U1092 ( .A(A[13]), .B(B[24]), .Y(n1082) );
  OAI22X1 U1093 ( .A0(n1063), .A1(n1062), .B0(n1090), .B1(n1087), .Y(n1097) );
  CMPR32X1 U1094 ( .A(n1066), .B(n1065), .C(n1064), .CO(n1100), .S(n1055) );
  NAND2XL U1095 ( .A(n1070), .B(n1069), .Y(mult_x_1_n81) );
  OAI21XL U1096 ( .A0(n1179), .A1(n1078), .B0(n1077), .Y(n1081) );
  XNOR2X1 U1097 ( .A(A[13]), .B(n1117), .Y(n1093) );
  CMPR32X1 U1098 ( .A(n1085), .B(n1084), .C(n1083), .CO(n1104), .S(n1101) );
  OAI22X1 U1099 ( .A0(n1094), .A1(n1093), .B0(n1123), .B1(n1120), .Y(n1128) );
  CMPR32X1 U1100 ( .A(n1097), .B(n1096), .C(n1095), .CO(n1114), .S(n1103) );
  CMPR32X1 U1101 ( .A(n1102), .B(n1101), .C(n1100), .CO(n1107), .S(n1067) );
  CMPR32X1 U1102 ( .A(n1105), .B(n1104), .C(n1103), .CO(n1099), .S(n1106) );
  OAI21XL U1103 ( .A0(n1109), .A1(n1184), .B0(n1185), .Y(n1173) );
  OAI21XL U1104 ( .A0(n1179), .A1(n1111), .B0(n1110), .Y(n1113) );
  CMPR32X1 U1105 ( .A(n1116), .B(n1115), .C(n1114), .CO(n1125), .S(n1098) );
  CMPR32X1 U1106 ( .A(n1128), .B(n1127), .C(n1126), .CO(n1137), .S(n1124) );
  XNOR2XL U1107 ( .A(n1130), .B(n1129), .Y(n1131) );
  XNOR2XL U1108 ( .A(n1169), .B(n1168), .Y(n1259) );
  AOI21XL U1109 ( .A0(n232), .A1(n1176), .B0(n1175), .Y(n1177) );
  OAI21XL U1110 ( .A0(n1179), .A1(n1178), .B0(n1177), .Y(n1180) );
endmodule


module FFT2048_DW02_mult_2_stage_J1_19 ( A, B, TC, CLK, PRODUCT );
  input [25:0] A;
  input [16:0] B;
  output [42:0] PRODUCT;
  input TC, CLK;
  wire   n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, mult_x_1_n665, mult_x_1_n650, mult_x_1_n649,
         mult_x_1_n634, mult_x_1_n633, mult_x_1_n618, mult_x_1_n617,
         mult_x_1_n602, mult_x_1_n601, mult_x_1_n586, mult_x_1_n585,
         mult_x_1_n570, mult_x_1_n569, mult_x_1_n554, mult_x_1_n553,
         mult_x_1_n538, mult_x_1_n537, mult_x_1_n522, mult_x_1_n521,
         mult_x_1_n508, mult_x_1_n507, mult_x_1_n494, mult_x_1_n321,
         mult_x_1_n316, mult_x_1_n309, mult_x_1_n305, mult_x_1_n298,
         mult_x_1_n293, mult_x_1_n292, mult_x_1_n287, mult_x_1_n286,
         mult_x_1_n282, mult_x_1_n281, mult_x_1_n195, mult_x_1_n194,
         mult_x_1_n184, mult_x_1_n183, mult_x_1_n177, mult_x_1_n176,
         mult_x_1_n170, mult_x_1_n169, mult_x_1_n161, mult_x_1_n160,
         mult_x_1_n152, mult_x_1_n151, mult_x_1_n137, mult_x_1_n136,
         mult_x_1_n130, mult_x_1_n129, mult_x_1_n121, mult_x_1_n120,
         mult_x_1_n110, mult_x_1_n109, mult_x_1_n86, mult_x_1_n85,
         mult_x_1_n84, mult_x_1_n83, mult_x_1_n58, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317;

  DFFHQXL mult_x_1_clk_r_REG12_S1 ( .D(mult_x_1_n183), .CK(CLK), .Q(n1279) );
  DFFHQXL mult_x_1_clk_r_REG16_S1 ( .D(mult_x_1_n169), .CK(CLK), .Q(n1275) );
  DFFHQXL mult_x_1_clk_r_REG18_S1 ( .D(mult_x_1_n160), .CK(CLK), .Q(n1273) );
  DFFHQXL mult_x_1_clk_r_REG20_S1 ( .D(mult_x_1_n151), .CK(CLK), .Q(n1271) );
  DFFHQX4 mult_x_1_clk_r_REG42_S1 ( .D(mult_x_1_n665), .CK(CLK), .Q(n1316) );
  DFFHQX4 mult_x_1_clk_r_REG41_S1 ( .D(mult_x_1_n650), .CK(CLK), .Q(n1315) );
  DFFHQX4 mult_x_1_clk_r_REG40_S1 ( .D(mult_x_1_n649), .CK(CLK), .Q(n1314) );
  DFFHQX4 mult_x_1_clk_r_REG39_S1 ( .D(mult_x_1_n634), .CK(CLK), .Q(n1313) );
  DFFHQX4 mult_x_1_clk_r_REG38_S1 ( .D(mult_x_1_n633), .CK(CLK), .Q(n1312) );
  DFFHQX4 mult_x_1_clk_r_REG37_S1 ( .D(mult_x_1_n618), .CK(CLK), .Q(n1311) );
  DFFHQX4 mult_x_1_clk_r_REG36_S1 ( .D(mult_x_1_n617), .CK(CLK), .Q(n1310) );
  DFFHQX4 mult_x_1_clk_r_REG35_S1 ( .D(mult_x_1_n602), .CK(CLK), .Q(n1309) );
  DFFHQX4 mult_x_1_clk_r_REG34_S1 ( .D(mult_x_1_n601), .CK(CLK), .Q(n1308) );
  DFFHQX4 mult_x_1_clk_r_REG33_S1 ( .D(mult_x_1_n586), .CK(CLK), .Q(n1307) );
  DFFHQX4 mult_x_1_clk_r_REG32_S1 ( .D(mult_x_1_n585), .CK(CLK), .Q(n1306) );
  DFFHQX4 mult_x_1_clk_r_REG31_S1 ( .D(mult_x_1_n570), .CK(CLK), .Q(n1305) );
  DFFHQX4 mult_x_1_clk_r_REG30_S1 ( .D(mult_x_1_n569), .CK(CLK), .Q(n1304) );
  DFFHQX4 mult_x_1_clk_r_REG1_S1 ( .D(mult_x_1_n554), .CK(CLK), .Q(n1303) );
  DFFHQX4 mult_x_1_clk_r_REG0_S1 ( .D(mult_x_1_n553), .CK(CLK), .Q(n1302) );
  DFFHQX4 mult_x_1_clk_r_REG3_S1 ( .D(mult_x_1_n538), .CK(CLK), .Q(n1301) );
  DFFHQX4 mult_x_1_clk_r_REG2_S1 ( .D(mult_x_1_n537), .CK(CLK), .Q(n1300) );
  DFFHQX4 mult_x_1_clk_r_REG5_S1 ( .D(mult_x_1_n522), .CK(CLK), .Q(n1299) );
  DFFHQX4 mult_x_1_clk_r_REG4_S1 ( .D(mult_x_1_n521), .CK(CLK), .Q(n1298) );
  DFFHQX4 mult_x_1_clk_r_REG7_S1 ( .D(mult_x_1_n508), .CK(CLK), .Q(n1297) );
  DFFHQX4 mult_x_1_clk_r_REG56_S1 ( .D(mult_x_1_n309), .CK(CLK), .Q(n1293) );
  DFFHQX4 mult_x_1_clk_r_REG48_S1 ( .D(mult_x_1_n292), .CK(CLK), .Q(n1287) );
  DFFHQX4 mult_x_1_clk_r_REG53_S1 ( .D(mult_x_1_n305), .CK(CLK), .Q(n1260) );
  DFFHQX4 mult_x_1_clk_r_REG54_S1 ( .D(n1317), .CK(CLK), .Q(n1259) );
  DFFHQX4 mult_x_1_clk_r_REG50_S1 ( .D(mult_x_1_n298), .CK(CLK), .Q(n1258) );
  DFFHQX4 mult_x_1_clk_r_REG51_S1 ( .D(n24), .CK(CLK), .Q(n1257) );
  DFFHQXL mult_x_1_clk_r_REG9_S1 ( .D(mult_x_1_n195), .CK(CLK), .Q(n1282) );
  DFFHQXL mult_x_1_clk_r_REG15_S1 ( .D(mult_x_1_n170), .CK(CLK), .Q(n1276) );
  DFFHQXL mult_x_1_clk_r_REG21_S1 ( .D(mult_x_1_n137), .CK(CLK), .Q(n1270) );
  DFFHQXL mult_x_1_clk_r_REG17_S1 ( .D(mult_x_1_n161), .CK(CLK), .Q(n1274) );
  DFFHQXL mult_x_1_clk_r_REG19_S1 ( .D(mult_x_1_n152), .CK(CLK), .Q(n1272) );
  DFFHQXL clk_r_REG62_S1 ( .D(n1332), .CK(CLK), .Q(PRODUCT[9]) );
  DFFHQXL mult_x_1_clk_r_REG14_S1 ( .D(mult_x_1_n176), .CK(CLK), .Q(n1277) );
  DFFHQXL mult_x_1_clk_r_REG60_S1 ( .D(mult_x_1_n321), .CK(CLK), .Q(n1261) );
  DFFHQXL mult_x_1_clk_r_REG13_S1 ( .D(mult_x_1_n177), .CK(CLK), .Q(n1278) );
  DFFHQXL mult_x_1_clk_r_REG10_S1 ( .D(mult_x_1_n194), .CK(CLK), .Q(n1281) );
  DFFHQXL clk_r_REG61_S1 ( .D(n1331), .CK(CLK), .Q(PRODUCT[10]) );
  DFFHQXL mult_x_1_clk_r_REG11_S1 ( .D(mult_x_1_n184), .CK(CLK), .Q(n1280) );
  DFFHQXL clk_r_REG68_S1 ( .D(n1338), .CK(CLK), .Q(PRODUCT[3]) );
  DFFHQXL mult_x_1_clk_r_REG28_S1 ( .D(mult_x_1_n109), .CK(CLK), .Q(n1263) );
  DFFHQXL clk_r_REG59_S1 ( .D(n1330), .CK(CLK), .Q(PRODUCT[11]) );
  DFFHQXL clk_r_REG63_S1 ( .D(n1333), .CK(CLK), .Q(PRODUCT[8]) );
  DFFHQXL clk_r_REG65_S1 ( .D(n1335), .CK(CLK), .Q(PRODUCT[6]) );
  DFFHQXL clk_r_REG67_S1 ( .D(n1337), .CK(CLK), .Q(PRODUCT[4]) );
  DFFHQXL clk_r_REG70_S1 ( .D(n1340), .CK(CLK), .Q(PRODUCT[1]) );
  DFFHQXL clk_r_REG71_S1 ( .D(n1341), .CK(CLK), .Q(PRODUCT[0]) );
  DFFHQXL clk_r_REG64_S1 ( .D(n1334), .CK(CLK), .Q(PRODUCT[7]) );
  DFFHQXL clk_r_REG66_S1 ( .D(n1336), .CK(CLK), .Q(PRODUCT[5]) );
  DFFHQXL clk_r_REG69_S1 ( .D(n1339), .CK(CLK), .Q(PRODUCT[2]) );
  DFFHQXL mult_x_1_clk_r_REG49_S1 ( .D(mult_x_1_n83), .CK(CLK), .Q(n1289) );
  DFFHQXL mult_x_1_clk_r_REG23_S1 ( .D(mult_x_1_n130), .CK(CLK), .Q(n1268) );
  DFFHQXL mult_x_1_clk_r_REG24_S1 ( .D(mult_x_1_n129), .CK(CLK), .Q(n1267) );
  DFFHQXL mult_x_1_clk_r_REG25_S1 ( .D(mult_x_1_n121), .CK(CLK), .Q(n1266) );
  DFFHQXL mult_x_1_clk_r_REG26_S1 ( .D(mult_x_1_n120), .CK(CLK), .Q(n1265) );
  DFFHQXL mult_x_1_clk_r_REG27_S1 ( .D(mult_x_1_n110), .CK(CLK), .Q(n1264) );
  DFFHQXL mult_x_1_clk_r_REG29_S1 ( .D(mult_x_1_n58), .CK(CLK), .Q(n1262) );
  DFFHQXL mult_x_1_clk_r_REG22_S1 ( .D(mult_x_1_n136), .CK(CLK), .Q(n1269) );
  DFFHQXL mult_x_1_clk_r_REG57_S1 ( .D(mult_x_1_n86), .CK(CLK), .Q(n1292) );
  DFFHQX1 mult_x_1_clk_r_REG47_S1 ( .D(mult_x_1_n293), .CK(CLK), .Q(n1288) );
  DFFHQXL mult_x_1_clk_r_REG52_S1 ( .D(mult_x_1_n84), .CK(CLK), .Q(n1290) );
  DFFHQX1 mult_x_1_clk_r_REG43_S1 ( .D(mult_x_1_n282), .CK(CLK), .Q(n1284) );
  DFFHQX1 mult_x_1_clk_r_REG46_S1 ( .D(mult_x_1_n286), .CK(CLK), .Q(n1285) );
  DFFHQX1 mult_x_1_clk_r_REG45_S1 ( .D(mult_x_1_n287), .CK(CLK), .Q(n1286) );
  DFFHQX2 mult_x_1_clk_r_REG44_S1 ( .D(mult_x_1_n281), .CK(CLK), .Q(n1283) );
  DFFHQX1 mult_x_1_clk_r_REG55_S1 ( .D(mult_x_1_n85), .CK(CLK), .Q(n1291) );
  DFFHQX1 mult_x_1_clk_r_REG58_S1 ( .D(mult_x_1_n316), .CK(CLK), .Q(n1294) );
  DFFHQX2 mult_x_1_clk_r_REG8_S1 ( .D(mult_x_1_n494), .CK(CLK), .Q(n1295) );
  DFFHQX2 mult_x_1_clk_r_REG6_S1 ( .D(mult_x_1_n507), .CK(CLK), .Q(n1296) );
  ADDFHX1 U1 ( .A(n746), .B(n745), .CI(n744), .CO(mult_x_1_n507), .S(
        mult_x_1_n508) );
  ADDFHX1 U2 ( .A(n770), .B(n769), .CI(n768), .CO(mult_x_1_n521), .S(
        mult_x_1_n522) );
  ADDFHX2 U3 ( .A(n912), .B(n911), .CI(n910), .CO(n873), .S(n913) );
  ADDFX2 U4 ( .A(n1036), .B(n1035), .CI(n1034), .CO(mult_x_1_n665), .S(n599)
         );
  ADDFHX1 U5 ( .A(n833), .B(n832), .CI(n831), .CO(n802), .S(n834) );
  ADDFHX1 U6 ( .A(n800), .B(n799), .CI(n798), .CO(n769), .S(n801) );
  ADDFHX1 U7 ( .A(n767), .B(n766), .CI(n765), .CO(n745), .S(n768) );
  ADDFHX1 U8 ( .A(n705), .B(n704), .CI(n703), .CO(n445), .S(mult_x_1_n494) );
  CMPR32X1 U9 ( .A(n909), .B(n908), .C(n907), .CO(n912), .S(n954) );
  CMPR32X1 U10 ( .A(n868), .B(n867), .C(n866), .CO(n871), .S(n910) );
  OAI21XL U11 ( .A0(n23), .A1(n22), .B0(n21), .Y(n767) );
  ADDFHX1 U12 ( .A(n1027), .B(n1026), .CI(n1025), .CO(n1032), .S(n1034) );
  ADDFHX1 U13 ( .A(n1085), .B(n1084), .CI(n1083), .CO(n659), .S(n1096) );
  ADDFHX2 U14 ( .A(n573), .B(n572), .CI(n571), .CO(n1026), .S(n604) );
  ADDFHX1 U15 ( .A(n1009), .B(n1008), .CI(n1007), .CO(n1030), .S(n1025) );
  ADDFHX1 U16 ( .A(n388), .B(n387), .CI(n386), .CO(n371), .S(n443) );
  ADDFHX2 U17 ( .A(n582), .B(n581), .CI(n580), .CO(n597), .S(n624) );
  CMPR32X1 U18 ( .A(n1091), .B(n1090), .C(n1089), .CO(n1099), .S(n1101) );
  ADDFHX1 U19 ( .A(n542), .B(n541), .CI(n540), .CO(n549), .S(n606) );
  CMPR32X1 U20 ( .A(n1071), .B(n1070), .C(n1069), .CO(n1089), .S(n1074) );
  CMPR32X1 U21 ( .A(n1065), .B(n1064), .C(n1063), .CO(n1094), .S(n1091) );
  CMPR32X1 U22 ( .A(n679), .B(n678), .C(n677), .CO(n1062), .S(n674) );
  OAI22X1 U23 ( .A0(n1161), .A1(n962), .B0(n920), .B1(n1162), .Y(n54) );
  CLKBUFX8 U24 ( .A(n397), .Y(n1162) );
  CMPR32X1 U25 ( .A(n79), .B(n78), .C(n77), .CO(n150), .S(n80) );
  CLKBUFX8 U26 ( .A(B[15]), .Y(n209) );
  BUFX8 U27 ( .A(n966), .Y(n1139) );
  BUFX3 U28 ( .A(n196), .Y(n8) );
  BUFX3 U29 ( .A(n183), .Y(n6) );
  NAND2X2 U30 ( .A(n397), .B(n14), .Y(n422) );
  BUFX4 U31 ( .A(n518), .Y(n9) );
  BUFX3 U32 ( .A(n161), .Y(n942) );
  CLKBUFX8 U33 ( .A(n212), .Y(n972) );
  BUFX4 U34 ( .A(n69), .Y(n7) );
  BUFX3 U35 ( .A(n618), .Y(n939) );
  BUFX3 U36 ( .A(n586), .Y(n937) );
  NAND2X1 U37 ( .A(n67), .B(n586), .Y(n618) );
  OAI21XL U38 ( .A0(n1250), .A1(n1048), .B0(n1049), .Y(n382) );
  XOR2X1 U39 ( .A(n1047), .B(n1046), .Y(PRODUCT[21]) );
  XOR2X1 U40 ( .A(n1250), .B(n1042), .Y(PRODUCT[29]) );
  OAI21XL U41 ( .A0(n507), .A1(n506), .B0(n238), .Y(n512) );
  XOR2X1 U42 ( .A(n241), .B(n601), .Y(PRODUCT[17]) );
  INVX2 U43 ( .A(n15), .Y(n241) );
  NAND2X1 U44 ( .A(n240), .B(n237), .Y(n242) );
  OAI21XL U45 ( .A0(n238), .A1(n508), .B0(n509), .Y(n29) );
  NOR2X1 U46 ( .A(n501), .B(n1043), .Y(n484) );
  NOR2X2 U47 ( .A(n1301), .B(n1302), .Y(n473) );
  NAND2X2 U48 ( .A(n1312), .B(n1311), .Y(n1044) );
  NOR2X1 U49 ( .A(n1297), .B(n1298), .Y(n455) );
  OAI21XL U50 ( .A0(n1281), .A1(n1040), .B0(n1282), .Y(n380) );
  NOR2X1 U51 ( .A(n1311), .B(n1312), .Y(n1043) );
  AOI21XL U52 ( .A0(n380), .A1(n252), .B0(n251), .Y(n1246) );
  XNOR2XL U53 ( .A(n312), .B(n311), .Y(PRODUCT[33]) );
  XNOR2XL U54 ( .A(B[1]), .B(n919), .Y(n73) );
  XNOR2XL U55 ( .A(n68), .B(n890), .Y(n72) );
  XNOR2XL U56 ( .A(n68), .B(n851), .Y(n651) );
  BUFX1 U57 ( .A(A[18]), .Y(n853) );
  XNOR2XL U58 ( .A(n888), .B(n887), .Y(n929) );
  BUFX1 U59 ( .A(A[12]), .Y(n883) );
  BUFX1 U60 ( .A(A[15]), .Y(n896) );
  BUFX1 U61 ( .A(A[10]), .Y(n851) );
  BUFX1 U62 ( .A(A[21]), .Y(n1119) );
  XNOR2XL U63 ( .A(n209), .B(n896), .Y(n331) );
  XNOR2XL U64 ( .A(n1220), .B(n1219), .Y(PRODUCT[39]) );
  ADDHXL U65 ( .A(n128), .B(n127), .CO(n143), .S(n151) );
  XNOR2XL U66 ( .A(n712), .B(n1119), .Y(n353) );
  XNOR2XL U67 ( .A(n362), .B(n896), .Y(n413) );
  XNOR2XL U68 ( .A(n209), .B(n1119), .Y(n230) );
  ADDFX2 U69 ( .A(n82), .B(n81), .CI(n80), .CO(n118), .S(n117) );
  BUFX8 U70 ( .A(n422), .Y(n1161) );
  ADDFX2 U71 ( .A(n673), .B(n672), .CI(n671), .CO(n1058), .S(n1069) );
  XNOR2XL U72 ( .A(n1198), .B(n1197), .Y(n1334) );
  XOR2XL U73 ( .A(n1203), .B(n1202), .Y(n1335) );
  INVX1 U74 ( .A(n712), .Y(n132) );
  BUFX3 U75 ( .A(B[9]), .Y(n712) );
  INVX1 U76 ( .A(n286), .Y(n185) );
  XOR2X1 U77 ( .A(n516), .B(n515), .Y(PRODUCT[18]) );
  NAND2X1 U78 ( .A(n39), .B(n26), .Y(n958) );
  XOR2X1 U79 ( .A(n56), .B(n1017), .Y(n1019) );
  OR2X2 U80 ( .A(n691), .B(n690), .Y(n689) );
  ADDFHX1 U81 ( .A(n874), .B(n873), .CI(n872), .CO(mult_x_1_n569), .S(
        mult_x_1_n570) );
  ADDFHX2 U82 ( .A(n871), .B(n870), .CI(n869), .CO(n835), .S(n872) );
  NAND2X1 U83 ( .A(n17), .B(n16), .Y(n344) );
  NOR2X1 U84 ( .A(n119), .B(n118), .Y(n1194) );
  ADDFHX1 U85 ( .A(n151), .B(n150), .CI(n149), .CO(n152), .S(n119) );
  NOR2X1 U86 ( .A(n1158), .B(n210), .Y(n232) );
  NOR2X1 U87 ( .A(n1158), .B(n258), .Y(n273) );
  NOR2X1 U88 ( .A(n1158), .B(n211), .Y(n222) );
  NAND2X1 U89 ( .A(n1041), .B(n1040), .Y(n1042) );
  NAND2X1 U90 ( .A(n310), .B(n1276), .Y(n311) );
  INVX1 U91 ( .A(n1279), .Y(n1051) );
  NAND2X1 U92 ( .A(n1297), .B(n1298), .Y(n456) );
  INVX1 U93 ( .A(n1265), .Y(n1211) );
  INVX1 U94 ( .A(n1271), .Y(n1172) );
  ADDFHX1 U95 ( .A(n959), .B(n958), .CI(n957), .CO(mult_x_1_n601), .S(
        mult_x_1_n602) );
  ADDFHX1 U96 ( .A(n1021), .B(n1020), .CI(n1019), .CO(mult_x_1_n633), .S(
        mult_x_1_n634) );
  NAND2X1 U97 ( .A(n1096), .B(n1095), .Y(n1097) );
  ADDFHX1 U98 ( .A(n915), .B(n914), .CI(n913), .CO(mult_x_1_n585), .S(
        mult_x_1_n586) );
  ADDFHX1 U99 ( .A(n836), .B(n835), .CI(n834), .CO(mult_x_1_n553), .S(
        mult_x_1_n554) );
  ADDFHX1 U100 ( .A(n803), .B(n802), .CI(n801), .CO(mult_x_1_n537), .S(
        mult_x_1_n538) );
  ADDFHX1 U101 ( .A(n956), .B(n955), .CI(n954), .CO(n914), .S(n957) );
  OAI2BB1XL U102 ( .A0N(n944), .A1N(n36), .B0(n35), .Y(n953) );
  ADDFHX1 U103 ( .A(n830), .B(n829), .CI(n828), .CO(n833), .S(n869) );
  ADDFHX1 U104 ( .A(n797), .B(n796), .CI(n795), .CO(n800), .S(n831) );
  NOR2X1 U105 ( .A(n117), .B(n116), .Y(n1199) );
  NOR2X1 U106 ( .A(n1158), .B(n1120), .Y(n1133) );
  NOR2X1 U107 ( .A(n1158), .B(n226), .Y(n1117) );
  OAI2BB1XL U108 ( .A0N(n845), .A1N(n972), .B0(n214), .Y(n220) );
  OAI2BB1XL U109 ( .A0N(n918), .A1N(n7), .B0(n262), .Y(n296) );
  INVXL U110 ( .A(n8), .Y(n38) );
  OAI22XL U111 ( .A0(n939), .A1(n198), .B0(n937), .B1(n652), .Y(n677) );
  NAND2X1 U112 ( .A(n62), .B(n64), .Y(n69) );
  XNOR2X1 U113 ( .A(n256), .B(n255), .Y(PRODUCT[35]) );
  NOR2X1 U114 ( .A(n1239), .B(n1177), .Y(n1209) );
  NAND2X1 U115 ( .A(n503), .B(n502), .Y(n504) );
  NAND2X1 U116 ( .A(n1045), .B(n1044), .Y(n1046) );
  INVX1 U117 ( .A(n468), .Y(n481) );
  NAND2X1 U118 ( .A(n1051), .B(n1280), .Y(n381) );
  NAND2X1 U119 ( .A(n1054), .B(n1278), .Y(n1055) );
  NAND2X1 U120 ( .A(n1299), .B(n1300), .Y(n464) );
  BUFX2 U121 ( .A(A[19]), .Y(n887) );
  BUFX2 U122 ( .A(A[23]), .Y(n1145) );
  INVXL U123 ( .A(n1293), .Y(n661) );
  INVX1 U124 ( .A(n1273), .Y(n1170) );
  BUFX2 U125 ( .A(A[17]), .Y(n894) );
  BUFX2 U126 ( .A(A[13]), .Y(n916) );
  BUFX2 U127 ( .A(A[3]), .Y(n932) );
  INVXL U128 ( .A(n1285), .Y(n600) );
  INVXL U129 ( .A(n666), .Y(n696) );
  ADDFHX1 U130 ( .A(n997), .B(n996), .CI(n995), .CO(mult_x_1_n617), .S(
        mult_x_1_n618) );
  NAND2XL U131 ( .A(n630), .B(n631), .Y(n43) );
  INVX1 U132 ( .A(n1075), .Y(n1105) );
  NAND2X1 U133 ( .A(n691), .B(n690), .Y(n1106) );
  ADDFHX1 U134 ( .A(n953), .B(n952), .CI(n951), .CO(n956), .S(n992) );
  ADDFHX2 U135 ( .A(n625), .B(n624), .CI(n623), .CO(n603), .S(n629) );
  ADDFHX1 U136 ( .A(n1074), .B(n1073), .CI(n1072), .CO(n1076), .S(n691) );
  NAND2XL U137 ( .A(n299), .B(n18), .Y(n17) );
  ADDFHX2 U138 ( .A(n373), .B(n372), .CI(n371), .CO(n375), .S(n383) );
  ADDFHX2 U139 ( .A(n425), .B(n424), .CI(n423), .CO(n441), .S(n704) );
  OR2XL U140 ( .A(n1167), .B(n1166), .Y(n1169) );
  INVXL U141 ( .A(n631), .Y(n41) );
  ADDFHX2 U142 ( .A(n176), .B(n175), .CI(n174), .CO(n177), .S(n155) );
  NAND2BXL U143 ( .AN(n300), .B(n19), .Y(n18) );
  ADDFHX1 U144 ( .A(n188), .B(n187), .CI(n186), .CO(n687), .S(n199) );
  INVXL U145 ( .A(n301), .Y(n19) );
  ADDFHX1 U146 ( .A(n401), .B(n400), .CI(n399), .CO(n392), .S(n436) );
  ADDFHX1 U147 ( .A(n843), .B(n842), .CI(n841), .CO(n827), .S(n864) );
  ADDFHX1 U148 ( .A(n882), .B(n881), .CI(n880), .CO(n865), .S(n905) );
  ADDFHX1 U149 ( .A(n809), .B(n808), .CI(n807), .CO(n794), .S(n826) );
  ADDFHX1 U150 ( .A(n776), .B(n775), .CI(n774), .CO(n764), .S(n793) );
  OR2X2 U151 ( .A(n106), .B(n105), .Y(n104) );
  ADDFHX1 U152 ( .A(n142), .B(n141), .CI(n140), .CO(n147), .S(n149) );
  ADDFHX1 U153 ( .A(n173), .B(n172), .CI(n171), .CO(n186), .S(n176) );
  ADDFHX1 U154 ( .A(n925), .B(n924), .CI(n923), .CO(n906), .S(n949) );
  INVXL U155 ( .A(n261), .Y(n262) );
  AND2XL U156 ( .A(n1224), .B(n1223), .Y(n1340) );
  INVXL U157 ( .A(n615), .Y(n47) );
  OR2XL U158 ( .A(n1222), .B(n1221), .Y(n1224) );
  OAI2BB1XL U159 ( .A0N(n937), .A1N(n939), .B0(n357), .Y(n415) );
  XNOR2X1 U160 ( .A(n1207), .B(n1206), .Y(PRODUCT[38]) );
  XNOR2X1 U161 ( .A(n1188), .B(n1187), .Y(PRODUCT[36]) );
  XNOR2X1 U162 ( .A(n1183), .B(n1182), .Y(PRODUCT[37]) );
  XNOR2X1 U163 ( .A(n495), .B(n494), .Y(PRODUCT[24]) );
  OR2XL U164 ( .A(n1239), .B(n1245), .Y(n1249) );
  XOR2X1 U165 ( .A(n507), .B(n208), .Y(PRODUCT[19]) );
  NOR2BX1 U166 ( .AN(n13), .B(n1258), .Y(n628) );
  NAND2X1 U167 ( .A(n514), .B(n1284), .Y(n515) );
  BUFX2 U168 ( .A(A[20]), .Y(n848) );
  BUFX2 U169 ( .A(A[16]), .Y(n855) );
  BUFX2 U170 ( .A(A[22]), .Y(n1135) );
  BUFX2 U171 ( .A(A[14]), .Y(n875) );
  BUFX2 U172 ( .A(A[2]), .Y(n638) );
  BUFX2 U173 ( .A(A[9]), .Y(n892) );
  BUFX2 U174 ( .A(A[7]), .Y(n921) );
  BUFX2 U175 ( .A(A[8]), .Y(n878) );
  BUFX2 U176 ( .A(A[4]), .Y(n890) );
  BUFX2 U177 ( .A(A[1]), .Y(n578) );
  BUFX2 U178 ( .A(A[11]), .Y(n926) );
  NAND2XL U179 ( .A(n1260), .B(n1257), .Y(n13) );
  XOR2X1 U180 ( .A(n60), .B(n59), .Y(PRODUCT[16]) );
  OAI21X1 U181 ( .A0(n893), .A1(n6), .B0(n37), .Y(n36) );
  BUFX4 U182 ( .A(B[11]), .Y(n286) );
  XNOR2X1 U183 ( .A(n286), .B(n892), .Y(n934) );
  OAI2BB1X1 U184 ( .A0N(n1016), .A1N(n1018), .B0(n55), .Y(n996) );
  NAND2X1 U185 ( .A(n1309), .B(n1310), .Y(n502) );
  AOI21X1 U186 ( .A0(n470), .A1(n481), .B0(n469), .Y(n471) );
  NAND4X2 U187 ( .A(n12), .B(n11), .C(n10), .D(n1288), .Y(n15) );
  NAND2BX4 U188 ( .AN(n1287), .B(n1258), .Y(n10) );
  NAND3BX4 U189 ( .AN(n1287), .B(n1257), .C(n1260), .Y(n11) );
  NAND4BX4 U190 ( .AN(n1287), .B(n1257), .C(n1293), .D(n1259), .Y(n12) );
  XOR2X2 U191 ( .A(B[14]), .B(B[15]), .Y(n14) );
  XNOR2X4 U192 ( .A(B[14]), .B(B[13]), .Y(n397) );
  OAI21X1 U193 ( .A0(n1029), .A1(n1030), .B0(n1028), .Y(n58) );
  AOI21X1 U194 ( .A0(n15), .A1(n237), .B0(n239), .Y(n507) );
  AOI21X1 U195 ( .A0(n15), .A1(n600), .B0(n513), .Y(n516) );
  NAND2XL U196 ( .A(n300), .B(n301), .Y(n16) );
  XNOR3X2 U197 ( .A(n19), .B(n300), .C(n299), .Y(n339) );
  NAND2X2 U198 ( .A(n20), .B(n518), .Y(n966) );
  XNOR2X1 U199 ( .A(B[12]), .B(B[11]), .Y(n518) );
  XOR2X1 U200 ( .A(B[12]), .B(B[13]), .Y(n20) );
  NAND2BX1 U201 ( .AN(n1285), .B(n1286), .Y(n601) );
  OAI21XL U202 ( .A0(n760), .A1(n761), .B0(n759), .Y(n21) );
  INVX1 U203 ( .A(n760), .Y(n22) );
  INVX1 U204 ( .A(n761), .Y(n23) );
  XOR3X2 U205 ( .A(n761), .B(n760), .C(n759), .Y(n799) );
  OAI21XL U206 ( .A0(n1047), .A1(n485), .B0(n496), .Y(n500) );
  NOR2X2 U207 ( .A(n468), .B(n473), .Y(n447) );
  XNOR2X2 U208 ( .A(B[15]), .B(B[16]), .Y(n328) );
  NOR2XL U209 ( .A(n1279), .B(n1277), .Y(n252) );
  OAI21XL U210 ( .A0(n1246), .A1(n1177), .B0(n1176), .Y(n1215) );
  INVXL U211 ( .A(n1243), .Y(n1176) );
  NAND2X1 U212 ( .A(n66), .B(n74), .Y(n161) );
  NAND2XL U213 ( .A(n1170), .B(n1172), .Y(n1175) );
  INVXL U214 ( .A(n1274), .Y(n1173) );
  INVXL U215 ( .A(n1269), .Y(n1186) );
  NOR2XL U216 ( .A(n460), .B(n448), .Y(n452) );
  NAND2X1 U217 ( .A(n1307), .B(n1308), .Y(n498) );
  NOR2XL U218 ( .A(n1175), .B(n1275), .Y(n1238) );
  NOR2XL U219 ( .A(n1237), .B(n1263), .Y(n1242) );
  INVXL U220 ( .A(n1237), .Y(n1214) );
  BUFX1 U221 ( .A(A[5]), .Y(n919) );
  NAND2XL U222 ( .A(n1211), .B(n1266), .Y(n1206) );
  XOR2X1 U223 ( .A(n661), .B(n1290), .Y(PRODUCT[14]) );
  XNOR2X1 U224 ( .A(n209), .B(n890), .Y(n963) );
  OAI22XL U225 ( .A0(n931), .A1(n524), .B0(n567), .B1(n1037), .Y(n570) );
  NOR2XL U226 ( .A(n1158), .B(n520), .Y(n569) );
  NAND2BXL U227 ( .AN(n1038), .B(n1156), .Y(n520) );
  NOR2XL U228 ( .A(n1158), .B(n1136), .Y(n1149) );
  INVXL U229 ( .A(n1137), .Y(n1138) );
  BUFX3 U230 ( .A(n1015), .Y(n31) );
  CMPR32X1 U231 ( .A(n982), .B(n981), .C(n980), .CO(n991), .S(n1014) );
  OAI22XL U232 ( .A0(n942), .A1(n941), .B0(n654), .B1(n940), .Y(n980) );
  OAI22XL U233 ( .A0(n939), .A1(n938), .B0(n937), .B1(n936), .Y(n981) );
  AOI21XL U234 ( .A0(n121), .A1(n1193), .B0(n120), .Y(n697) );
  NAND2XL U235 ( .A(n97), .B(n96), .Y(n1226) );
  AOI21XL U236 ( .A0(n1234), .A1(n1235), .B0(n92), .Y(n1228) );
  INVXL U237 ( .A(n1233), .Y(n92) );
  OAI22XL U238 ( .A0(n1161), .A1(n1147), .B0(n1162), .B1(n1159), .Y(n1165) );
  INVXL U239 ( .A(n1238), .Y(n1177) );
  NAND2XL U240 ( .A(n1208), .B(n1211), .Y(n1237) );
  NAND2XL U241 ( .A(n1209), .B(n1186), .Y(n1180) );
  AOI21XL U242 ( .A0(n1215), .A1(n1186), .B0(n1178), .Y(n1179) );
  INVXL U243 ( .A(n1270), .Y(n1178) );
  INVXL U244 ( .A(n1267), .Y(n1181) );
  AOI21XL U245 ( .A0(n486), .A1(n488), .B0(n487), .Y(n489) );
  INVXL U246 ( .A(n486), .Y(n496) );
  AOI21XL U247 ( .A0(n1173), .A1(n1172), .B0(n1171), .Y(n1174) );
  INVXL U248 ( .A(n1272), .Y(n1171) );
  AOI21XL U249 ( .A0(n1212), .A1(n1211), .B0(n1210), .Y(n1240) );
  INVXL U250 ( .A(n1266), .Y(n1210) );
  AOI21X2 U251 ( .A0(n239), .A1(n240), .B0(n29), .Y(n28) );
  NOR2X2 U252 ( .A(n508), .B(n506), .Y(n240) );
  INVXL U253 ( .A(n379), .Y(n1048) );
  NAND2XL U254 ( .A(n1186), .B(n1270), .Y(n1187) );
  NAND2XL U255 ( .A(n379), .B(n1051), .Y(n1053) );
  AOI21XL U256 ( .A0(n380), .A1(n1051), .B0(n1050), .Y(n1052) );
  AOI21XL U257 ( .A0(n470), .A1(n452), .B0(n451), .Y(n453) );
  AOI21XL U258 ( .A0(n470), .A1(n447), .B0(n450), .Y(n462) );
  INVXL U259 ( .A(n448), .Y(n465) );
  OAI21X1 U260 ( .A0(n491), .A1(n498), .B0(n492), .Y(n27) );
  INVXL U261 ( .A(n501), .Y(n503) );
  INVX4 U262 ( .A(n449), .Y(n1047) );
  NAND3XL U263 ( .A(n1259), .B(n1293), .C(n1257), .Y(n61) );
  XNOR2XL U264 ( .A(n837), .B(n932), .Y(n159) );
  XNOR2XL U265 ( .A(n817), .B(n919), .Y(n160) );
  XNOR2XL U266 ( .A(n837), .B(n890), .Y(n195) );
  XNOR2XL U267 ( .A(n837), .B(n919), .Y(n650) );
  XNOR2XL U268 ( .A(n817), .B(n878), .Y(n653) );
  XNOR2X1 U269 ( .A(n712), .B(n919), .Y(n616) );
  XNOR2XL U270 ( .A(n837), .B(A[6]), .Y(n649) );
  XNOR2XL U271 ( .A(n817), .B(n892), .Y(n619) );
  XNOR2XL U272 ( .A(n837), .B(n921), .Y(n635) );
  XNOR2XL U273 ( .A(n817), .B(n921), .Y(n655) );
  XNOR2XL U274 ( .A(n817), .B(A[6]), .Y(n179) );
  NAND2BXL U275 ( .AN(n1038), .B(n286), .Y(n184) );
  XNOR2X1 U276 ( .A(n209), .B(n578), .Y(n527) );
  XNOR2XL U277 ( .A(n837), .B(n878), .Y(n591) );
  XNOR2X1 U278 ( .A(n286), .B(n919), .Y(n545) );
  XNOR2XL U279 ( .A(n837), .B(n892), .Y(n547) );
  XNOR2XL U280 ( .A(n817), .B(n851), .Y(n590) );
  XNOR2XL U281 ( .A(n817), .B(n926), .Y(n574) );
  XNOR2XL U282 ( .A(n837), .B(n1145), .Y(n330) );
  NAND2BXL U283 ( .AN(n1038), .B(n817), .Y(n75) );
  CLKINVX3 U284 ( .A(B[7]), .Y(n260) );
  XNOR2XL U285 ( .A(n837), .B(n1038), .Y(n70) );
  XNOR2XL U286 ( .A(n817), .B(n638), .Y(n71) );
  XNOR2XL U287 ( .A(n837), .B(n638), .Y(n135) );
  OAI22XL U288 ( .A0(n618), .A1(n129), .B0(n937), .B1(n162), .Y(n165) );
  NAND2X1 U289 ( .A(n50), .B(n49), .Y(n48) );
  OR2X2 U290 ( .A(n579), .B(n9), .Y(n49) );
  OR2X2 U291 ( .A(n636), .B(n1139), .Y(n50) );
  NOR2BX1 U292 ( .AN(n1038), .B(n1162), .Y(n615) );
  OAI22X1 U293 ( .A0(n931), .A1(n592), .B0(n577), .B1(n1037), .Y(n614) );
  CMPR32X1 U294 ( .A(n367), .B(n366), .C(n365), .CO(n350), .S(n406) );
  INVXL U295 ( .A(n334), .Y(n365) );
  OAI22XL U296 ( .A0(n1139), .A1(n363), .B0(n9), .B1(n327), .Y(n367) );
  XNOR2XL U297 ( .A(n837), .B(n848), .Y(n420) );
  XNOR2XL U298 ( .A(n817), .B(n1119), .Y(n720) );
  OAI22XL U299 ( .A0(n7), .A1(n395), .B0(n918), .B1(n360), .Y(n399) );
  OAI22X1 U300 ( .A0(n1161), .A1(n398), .B0(n1162), .B1(n359), .Y(n400) );
  XNOR2XL U301 ( .A(n817), .B(n1145), .Y(n414) );
  OAI22XL U302 ( .A0(n422), .A1(n733), .B0(n1162), .B1(n421), .Y(n716) );
  OAI22XL U303 ( .A0(n7), .A1(n732), .B0(n918), .B1(n420), .Y(n717) );
  XNOR2XL U304 ( .A(n837), .B(n887), .Y(n732) );
  OAI22XL U305 ( .A0(n931), .A1(n889), .B0(n849), .B1(n1037), .Y(n886) );
  NOR2X1 U306 ( .A(n328), .B(n891), .Y(n42) );
  OAI22XL U307 ( .A0(n931), .A1(n929), .B0(n889), .B1(n1037), .Y(n928) );
  XNOR2X1 U308 ( .A(n286), .B(A[6]), .Y(n544) );
  XNOR2XL U309 ( .A(n817), .B(n883), .Y(n543) );
  INVXL U310 ( .A(n209), .Y(n523) );
  XNOR2XL U311 ( .A(n837), .B(n851), .Y(n546) );
  INVXL U312 ( .A(n213), .Y(n214) );
  OAI22XL U313 ( .A0(n8), .A1(n219), .B0(n6), .B1(n217), .Y(n223) );
  OAI22XL U314 ( .A0(n1161), .A1(n218), .B0(n1162), .B1(n215), .Y(n225) );
  INVXL U315 ( .A(n1247), .Y(n1248) );
  NAND2XL U316 ( .A(n1218), .B(n1264), .Y(n1219) );
  OAI22XL U317 ( .A0(n939), .A1(n355), .B0(n937), .B1(n95), .Y(n96) );
  INVXL U318 ( .A(n68), .Y(n355) );
  NAND2BXL U319 ( .AN(n1038), .B(n68), .Y(n95) );
  OAI22XL U320 ( .A0(n1161), .A1(n230), .B0(n1162), .B1(n1118), .Y(n1124) );
  OAI22XL U321 ( .A0(n1161), .A1(n1118), .B0(n1162), .B1(n1131), .Y(n1134) );
  INVXL U322 ( .A(n1150), .Y(n1132) );
  NOR2XL U323 ( .A(n328), .B(n354), .Y(n417) );
  INVXL U324 ( .A(n356), .Y(n357) );
  ADDFX2 U325 ( .A(n562), .B(n561), .CI(n560), .CO(n1009), .S(n548) );
  OAI22XL U326 ( .A0(n942), .A1(n543), .B0(n654), .B1(n564), .Y(n560) );
  OAI22X1 U327 ( .A0(n939), .A1(n538), .B0(n937), .B1(n537), .Y(n561) );
  OAI22XL U328 ( .A0(n8), .A1(n544), .B0(n6), .B1(n536), .Y(n562) );
  OAI22XL U329 ( .A0(n942), .A1(n564), .B0(n654), .B1(n941), .Y(n999) );
  OAI22XL U330 ( .A0(n972), .A1(n563), .B0(n970), .B1(n971), .Y(n1000) );
  OAI22XL U331 ( .A0(n7), .A1(n566), .B0(n64), .B1(n961), .Y(n1006) );
  OAI22XL U332 ( .A0(n7), .A1(n961), .B0(n918), .B1(n960), .Y(n1003) );
  OAI22X1 U333 ( .A0(n1161), .A1(n963), .B0(n962), .B1(n1162), .Y(n1002) );
  NOR2BXL U334 ( .AN(n1038), .B(n937), .Y(n90) );
  OAI22XL U335 ( .A0(n931), .A1(n88), .B0(n93), .B1(n1037), .Y(n91) );
  OAI22XL U336 ( .A0(n939), .A1(n101), .B0(n937), .B1(n100), .Y(n111) );
  NOR2BXL U337 ( .AN(n1038), .B(n654), .Y(n113) );
  OAI22XL U338 ( .A0(n931), .A1(n99), .B0(n98), .B1(n1037), .Y(n112) );
  OAI22XL U339 ( .A0(n939), .A1(n100), .B0(n937), .B1(n83), .Y(n110) );
  OAI22XL U340 ( .A0(n161), .A1(n85), .B0(n654), .B1(n84), .Y(n109) );
  XNOR2XL U341 ( .A(n817), .B(n1038), .Y(n85) );
  NOR2XL U342 ( .A(n1158), .B(n1157), .Y(n1164) );
  OAI2BB1XL U343 ( .A0N(n1162), .A1N(n1161), .B0(n1160), .Y(n1163) );
  INVXL U344 ( .A(n1159), .Y(n1160) );
  NOR2XL U345 ( .A(n1158), .B(n1146), .Y(n1155) );
  INVXL U346 ( .A(n1165), .Y(n1154) );
  NAND2X1 U347 ( .A(n31), .B(n1014), .Y(n32) );
  NAND2X1 U348 ( .A(n1013), .B(n34), .Y(n33) );
  OR2X2 U349 ( .A(n1015), .B(n1014), .Y(n34) );
  OAI2BB1XL U350 ( .A0N(n51), .A1N(n967), .B0(n25), .Y(n950) );
  NAND2XL U351 ( .A(n968), .B(n54), .Y(n25) );
  NAND2BXL U352 ( .AN(n968), .B(n52), .Y(n51) );
  NAND2XL U353 ( .A(n91), .B(n90), .Y(n1233) );
  INVXL U354 ( .A(n1223), .Y(n1235) );
  INVXL U355 ( .A(n1230), .Y(n107) );
  NOR2XL U356 ( .A(n115), .B(n114), .Y(n1252) );
  NAND2XL U357 ( .A(n115), .B(n114), .Y(n1253) );
  OAI22XL U358 ( .A0(n931), .A1(n1038), .B0(n88), .B1(n1037), .Y(n1222) );
  NAND2XL U359 ( .A(n89), .B(n931), .Y(n1221) );
  NAND2BXL U360 ( .AN(n1038), .B(B[1]), .Y(n89) );
  NAND2XL U361 ( .A(n1222), .B(n1221), .Y(n1223) );
  NAND2XL U362 ( .A(n106), .B(n105), .Y(n1230) );
  INVXL U363 ( .A(n1193), .Y(n1202) );
  NOR2XL U364 ( .A(n1269), .B(n1267), .Y(n1208) );
  INVXL U365 ( .A(n1209), .Y(n1185) );
  INVXL U366 ( .A(n1215), .Y(n1184) );
  OAI21X1 U367 ( .A0(n1286), .A1(n1283), .B0(n1284), .Y(n239) );
  NAND2XL U368 ( .A(n1209), .B(n1208), .Y(n1205) );
  NAND2XL U369 ( .A(n1181), .B(n1268), .Y(n1182) );
  INVXL U370 ( .A(n1275), .Y(n310) );
  INVXL U371 ( .A(n480), .Y(n469) );
  NAND2XL U372 ( .A(n1301), .B(n1302), .Y(n474) );
  INVXL U373 ( .A(n473), .Y(n475) );
  INVXL U374 ( .A(n491), .Y(n493) );
  XNOR2X1 U375 ( .A(n500), .B(n499), .Y(PRODUCT[23]) );
  INVXL U376 ( .A(n484), .Y(n485) );
  INVXL U377 ( .A(n1286), .Y(n513) );
  XNOR2XL U378 ( .A(n286), .B(n1038), .Y(n197) );
  XNOR2XL U379 ( .A(n286), .B(n578), .Y(n648) );
  XNOR2XL U380 ( .A(n888), .B(n926), .Y(n646) );
  OAI22XL U381 ( .A0(n169), .A1(n168), .B0(n181), .B1(n1037), .Y(n190) );
  OAI22X1 U382 ( .A0(n972), .A1(n170), .B0(n970), .B1(n180), .Y(n189) );
  XNOR2XL U383 ( .A(n1156), .B(n916), .Y(n329) );
  XNOR2XL U384 ( .A(n888), .B(A[25]), .Y(n714) );
  XNOR2XL U385 ( .A(n888), .B(A[24]), .Y(n727) );
  XNOR2XL U386 ( .A(n286), .B(n875), .Y(n750) );
  XNOR2XL U387 ( .A(n68), .B(n1135), .Y(n751) );
  XNOR2XL U388 ( .A(n817), .B(n848), .Y(n752) );
  XNOR2XL U389 ( .A(n286), .B(n916), .Y(n783) );
  XNOR2XL U390 ( .A(n68), .B(n1119), .Y(n784) );
  XNOR2XL U391 ( .A(n817), .B(n887), .Y(n785) );
  XNOR2XL U392 ( .A(n286), .B(n883), .Y(n815) );
  XNOR2XL U393 ( .A(n68), .B(n848), .Y(n816) );
  XNOR2XL U394 ( .A(n817), .B(n853), .Y(n818) );
  NAND2BXL U395 ( .AN(n1038), .B(n209), .Y(n522) );
  XNOR2XL U396 ( .A(n888), .B(n894), .Y(n567) );
  XNOR2XL U397 ( .A(n1156), .B(n855), .Y(n259) );
  XNOR2XL U398 ( .A(n1156), .B(n896), .Y(n290) );
  XNOR2XL U399 ( .A(n1156), .B(n875), .Y(n313) );
  XNOR2XL U400 ( .A(n68), .B(A[6]), .Y(n129) );
  AOI21XL U401 ( .A0(n1243), .A1(n1242), .B0(n1241), .Y(n1244) );
  NAND2XL U402 ( .A(n1238), .B(n1242), .Y(n1245) );
  NAND2XL U403 ( .A(n1209), .B(n1214), .Y(n1217) );
  INVXL U404 ( .A(n1240), .Y(n1213) );
  INVXL U405 ( .A(n1263), .Y(n1218) );
  NAND2XL U406 ( .A(n1170), .B(n1274), .Y(n284) );
  NAND2XL U407 ( .A(n1172), .B(n1272), .Y(n255) );
  OAI21XL U408 ( .A0(n1250), .A1(n254), .B0(n253), .Y(n256) );
  INVXL U409 ( .A(n1039), .Y(n1041) );
  XNOR2X1 U410 ( .A(n459), .B(n458), .Y(PRODUCT[28]) );
  NAND2XL U411 ( .A(n457), .B(n456), .Y(n458) );
  OAI21XL U412 ( .A0(n454), .A1(n1047), .B0(n453), .Y(n459) );
  XNOR2X1 U413 ( .A(n467), .B(n466), .Y(PRODUCT[27]) );
  NAND2XL U414 ( .A(n465), .B(n464), .Y(n466) );
  XNOR2X1 U415 ( .A(n477), .B(n476), .Y(PRODUCT[26]) );
  NAND2XL U416 ( .A(n475), .B(n474), .Y(n476) );
  OAI21XL U417 ( .A0(n1047), .A1(n472), .B0(n471), .Y(n477) );
  NAND2XL U418 ( .A(n481), .B(n480), .Y(n482) );
  OAI21XL U419 ( .A0(n1047), .A1(n1043), .B0(n1044), .Y(n505) );
  NOR2BXL U420 ( .AN(n1288), .B(n1287), .Y(n59) );
  NAND2XL U421 ( .A(n628), .B(n61), .Y(n60) );
  OAI22XL U422 ( .A0(n939), .A1(n162), .B0(n586), .B1(n198), .Y(n192) );
  OAI22XL U423 ( .A0(n161), .A1(n160), .B0(n654), .B1(n179), .Y(n193) );
  OAI22XL U424 ( .A0(n7), .A1(n159), .B0(n918), .B1(n195), .Y(n194) );
  OAI22XL U425 ( .A0(n161), .A1(n125), .B0(n654), .B1(n160), .Y(n171) );
  OAI22X1 U426 ( .A0(n7), .A1(n135), .B0(n918), .B1(n159), .Y(n173) );
  OAI22XL U427 ( .A0(n942), .A1(n655), .B0(n654), .B1(n653), .Y(n683) );
  OAI22XL U428 ( .A0(n939), .A1(n652), .B0(n937), .B1(n651), .Y(n684) );
  OAI22XL U429 ( .A0(n7), .A1(n650), .B0(n918), .B1(n649), .Y(n685) );
  NAND2BXL U430 ( .AN(n1038), .B(n1121), .Y(n593) );
  OAI22XL U431 ( .A0(n942), .A1(n653), .B0(n654), .B1(n619), .Y(n1066) );
  OAI22XL U432 ( .A0(n972), .A1(n667), .B0(n970), .B1(n616), .Y(n1068) );
  XNOR2XL U433 ( .A(n1156), .B(n1135), .Y(n1136) );
  XNOR2XL U434 ( .A(n1156), .B(n1119), .Y(n1120) );
  OAI22XL U435 ( .A0(n939), .A1(n617), .B0(n586), .B1(n585), .Y(n620) );
  OAI22XL U436 ( .A0(n972), .A1(n616), .B0(n970), .B1(n583), .Y(n622) );
  OAI22XL U437 ( .A0(n8), .A1(n647), .B0(n6), .B1(n639), .Y(n1063) );
  ADDFX2 U438 ( .A(n642), .B(n641), .CI(n640), .CO(n632), .S(n1093) );
  OAI22X1 U439 ( .A0(n7), .A1(n635), .B0(n918), .B1(n591), .Y(n641) );
  OAI22XL U440 ( .A0(n942), .A1(n619), .B0(n654), .B1(n590), .Y(n642) );
  OAI22XL U441 ( .A0(n942), .A1(n179), .B0(n654), .B1(n655), .Y(n682) );
  OAI22XL U442 ( .A0(n972), .A1(n180), .B0(n970), .B1(n668), .Y(n681) );
  XNOR2XL U443 ( .A(B[16]), .B(n883), .Y(n354) );
  OAI22XL U444 ( .A0(n1139), .A1(n413), .B0(n9), .B1(n363), .Y(n403) );
  OAI22XL U445 ( .A0(n972), .A1(n418), .B0(n845), .B1(n361), .Y(n404) );
  INVXL U446 ( .A(n714), .Y(n428) );
  XNOR2XL U447 ( .A(n286), .B(n896), .Y(n718) );
  XNOR2XL U448 ( .A(n68), .B(n1145), .Y(n719) );
  XNOR2XL U449 ( .A(n837), .B(n853), .Y(n771) );
  OAI22XL U450 ( .A0(n931), .A1(n813), .B0(n781), .B1(n780), .Y(n812) );
  OAI22XL U451 ( .A0(n972), .A1(n777), .B0(n845), .B1(n724), .Y(n758) );
  ADDFX2 U452 ( .A(n755), .B(n754), .CI(n753), .CO(n761), .S(n796) );
  OAI22XL U453 ( .A0(n942), .A1(n752), .B0(n654), .B1(n720), .Y(n753) );
  OAI22X1 U454 ( .A0(n939), .A1(n751), .B0(n937), .B1(n719), .Y(n754) );
  OAI22XL U455 ( .A0(n8), .A1(n750), .B0(n6), .B1(n718), .Y(n755) );
  XNOR2XL U456 ( .A(n837), .B(n894), .Y(n804) );
  XNOR2XL U457 ( .A(n712), .B(n875), .Y(n844) );
  ADDFX2 U458 ( .A(n788), .B(n787), .CI(n786), .CO(n797), .S(n829) );
  OAI22XL U459 ( .A0(n942), .A1(n785), .B0(n654), .B1(n752), .Y(n786) );
  OAI22X1 U460 ( .A0(n939), .A1(n784), .B0(n937), .B1(n751), .Y(n787) );
  OAI22XL U461 ( .A0(n8), .A1(n783), .B0(n6), .B1(n750), .Y(n788) );
  XNOR2XL U462 ( .A(n837), .B(n855), .Y(n838) );
  CMPR32X1 U463 ( .A(n821), .B(n820), .C(n819), .CO(n830), .S(n867) );
  OAI22XL U464 ( .A0(n942), .A1(n818), .B0(n654), .B1(n785), .Y(n819) );
  OAI22XL U465 ( .A0(n939), .A1(n816), .B0(n937), .B1(n784), .Y(n820) );
  OAI22XL U466 ( .A0(n8), .A1(n815), .B0(n6), .B1(n783), .Y(n821) );
  CMPR32X1 U467 ( .A(n859), .B(n858), .C(n857), .CO(n868), .S(n908) );
  OAI22XL U468 ( .A0(n942), .A1(n856), .B0(n654), .B1(n818), .Y(n857) );
  OAI22XL U469 ( .A0(n939), .A1(n854), .B0(n937), .B1(n816), .Y(n858) );
  OAI22XL U470 ( .A0(n8), .A1(n852), .B0(n6), .B1(n815), .Y(n859) );
  XNOR2XL U471 ( .A(n837), .B(n896), .Y(n876) );
  XNOR2XL U472 ( .A(n286), .B(n926), .Y(n852) );
  XNOR2XL U473 ( .A(n68), .B(n887), .Y(n854) );
  XNOR2XL U474 ( .A(n817), .B(n894), .Y(n856) );
  XNOR2XL U475 ( .A(n817), .B(n855), .Y(n897) );
  XNOR2XL U476 ( .A(n286), .B(n851), .Y(n893) );
  XNOR2XL U477 ( .A(n68), .B(n853), .Y(n895) );
  XNOR2XL U478 ( .A(n837), .B(n875), .Y(n917) );
  XNOR2X1 U479 ( .A(n209), .B(A[6]), .Y(n920) );
  XNOR2XL U480 ( .A(n1121), .B(n878), .Y(n922) );
  OAI22XL U481 ( .A0(n931), .A1(n930), .B0(n929), .B1(n1037), .Y(n974) );
  XNOR2XL U482 ( .A(n817), .B(n896), .Y(n940) );
  XNOR2XL U483 ( .A(n68), .B(n894), .Y(n936) );
  XNOR2XL U484 ( .A(n68), .B(n875), .Y(n538) );
  XNOR2XL U485 ( .A(n712), .B(n851), .Y(n971) );
  XNOR2XL U486 ( .A(n817), .B(n875), .Y(n941) );
  XNOR2XL U487 ( .A(n817), .B(n916), .Y(n564) );
  XNOR2XL U488 ( .A(n837), .B(n916), .Y(n960) );
  XNOR2XL U489 ( .A(n837), .B(n883), .Y(n961) );
  XNOR2X1 U490 ( .A(n1121), .B(A[6]), .Y(n965) );
  ADDFX2 U491 ( .A(n589), .B(n588), .CI(n587), .CO(n580), .S(n633) );
  OAI22X1 U492 ( .A0(n1161), .A1(n528), .B0(n1162), .B1(n527), .Y(n588) );
  OAI22XL U493 ( .A0(n972), .A1(n583), .B0(n970), .B1(n533), .Y(n589) );
  NOR2BXL U494 ( .AN(n1038), .B(n328), .Y(n531) );
  OAI22XL U495 ( .A0(n931), .A1(n525), .B0(n524), .B1(n1037), .Y(n530) );
  OAI22X1 U496 ( .A0(n1161), .A1(n527), .B0(n1162), .B1(n526), .Y(n529) );
  XNOR2XL U497 ( .A(B[16]), .B(n578), .Y(n517) );
  XNOR2XL U498 ( .A(n1121), .B(n890), .Y(n534) );
  XNOR2XL U499 ( .A(n1121), .B(n919), .Y(n565) );
  OAI22XL U500 ( .A0(n7), .A1(n591), .B0(n64), .B1(n547), .Y(n608) );
  OAI22XL U501 ( .A0(n939), .A1(n585), .B0(n937), .B1(n539), .Y(n610) );
  OAI22XL U502 ( .A0(n7), .A1(n547), .B0(n64), .B1(n546), .Y(n551) );
  OAI22XL U503 ( .A0(n942), .A1(n574), .B0(n654), .B1(n543), .Y(n553) );
  OAI22XL U504 ( .A0(n942), .A1(n590), .B0(n654), .B1(n574), .Y(n613) );
  OAI21XL U505 ( .A0(n47), .A1(n46), .B0(n45), .Y(n611) );
  XNOR2XL U506 ( .A(n286), .B(n1119), .Y(n292) );
  INVXL U507 ( .A(n221), .Y(n269) );
  OAI22XL U508 ( .A0(n1139), .A1(n288), .B0(n9), .B1(n268), .Y(n293) );
  OAI22XL U509 ( .A0(n972), .A1(n289), .B0(n845), .B1(n266), .Y(n295) );
  ADDFX2 U510 ( .A(n318), .B(n317), .CI(n316), .CO(n299), .S(n348) );
  OAI22XL U511 ( .A0(n8), .A1(n325), .B0(n6), .B1(n292), .Y(n316) );
  OAI22X1 U512 ( .A0(n1161), .A1(n323), .B0(n1162), .B1(n291), .Y(n317) );
  NOR2XL U513 ( .A(n1158), .B(n290), .Y(n318) );
  ADDFX2 U514 ( .A(n321), .B(n320), .CI(n319), .CO(n300), .S(n347) );
  INVXL U515 ( .A(n297), .Y(n319) );
  OAI22X1 U516 ( .A0(n972), .A1(n324), .B0(n845), .B1(n289), .Y(n320) );
  OAI22X1 U517 ( .A0(n1139), .A1(n326), .B0(n9), .B1(n288), .Y(n321) );
  CMPR32X1 U518 ( .A(n335), .B(n334), .C(n333), .CO(n349), .S(n387) );
  OAI2BB1XL U519 ( .A0N(n74), .A1N(n942), .B0(n315), .Y(n333) );
  NOR2XL U520 ( .A(n1158), .B(n313), .Y(n335) );
  INVXL U521 ( .A(n314), .Y(n315) );
  OAI22XL U522 ( .A0(n972), .A1(n353), .B0(n845), .B1(n324), .Y(n336) );
  OAI22XL U523 ( .A0(n7), .A1(n330), .B0(n918), .B1(n322), .Y(n338) );
  OAI22XL U524 ( .A0(n1161), .A1(n331), .B0(n1162), .B1(n323), .Y(n337) );
  OAI22XL U525 ( .A0(n8), .A1(n364), .B0(n6), .B1(n332), .Y(n368) );
  OAI22XL U526 ( .A0(n7), .A1(n360), .B0(n918), .B1(n330), .Y(n370) );
  OAI22XL U527 ( .A0(n8), .A1(n332), .B0(n6), .B1(n325), .Y(n352) );
  XNOR2XL U528 ( .A(n888), .B(n932), .Y(n99) );
  XNOR2XL U529 ( .A(n68), .B(n638), .Y(n100) );
  XNOR2XL U530 ( .A(n68), .B(n932), .Y(n83) );
  INVXL U531 ( .A(n817), .Y(n76) );
  NAND2BXL U532 ( .AN(n1038), .B(n837), .Y(n63) );
  OAI22XL U533 ( .A0(n161), .A1(n71), .B0(n654), .B1(n126), .Y(n140) );
  OAI22X1 U534 ( .A0(n7), .A1(n70), .B0(n918), .B1(n136), .Y(n141) );
  CMPR32X1 U535 ( .A(n145), .B(n144), .C(n143), .CO(n175), .S(n146) );
  OAI22XL U536 ( .A0(n618), .A1(n124), .B0(n937), .B1(n129), .Y(n145) );
  OAI22XL U537 ( .A0(n942), .A1(n126), .B0(n654), .B1(n125), .Y(n144) );
  OAI22XL U538 ( .A0(n7), .A1(n136), .B0(n918), .B1(n135), .Y(n137) );
  NOR2BXL U539 ( .AN(n1038), .B(n970), .Y(n139) );
  OAI2BB1XL U540 ( .A0N(n6), .A1N(n8), .B0(n228), .Y(n1115) );
  INVXL U541 ( .A(n227), .Y(n228) );
  OAI21XL U542 ( .A0(n697), .A1(n158), .B0(n157), .Y(n666) );
  NAND2X1 U543 ( .A(n700), .B(n1190), .Y(n158) );
  AOI21XL U544 ( .A0(n700), .A1(n698), .B0(n156), .Y(n157) );
  OAI22XL U545 ( .A0(n972), .A1(n361), .B0(n845), .B1(n353), .Y(n394) );
  CMPR32X1 U546 ( .A(n711), .B(n710), .C(n709), .CO(n437), .S(n730) );
  NOR2XL U547 ( .A(n328), .B(n396), .Y(n710) );
  OAI22XL U548 ( .A0(n7), .A1(n420), .B0(n918), .B1(n395), .Y(n711) );
  OAI22XL U549 ( .A0(n942), .A1(n720), .B0(n654), .B1(n706), .Y(n737) );
  ADDFX2 U550 ( .A(n437), .B(n436), .CI(n435), .CO(n424), .S(n742) );
  INVXL U551 ( .A(n416), .Y(n429) );
  OAI22XL U552 ( .A0(n942), .A1(n706), .B0(n654), .B1(n414), .Y(n430) );
  OAI22XL U553 ( .A0(n972), .A1(n713), .B0(n845), .B1(n418), .Y(n434) );
  OAI22XL U554 ( .A0(n8), .A1(n426), .B0(n6), .B1(n419), .Y(n433) );
  OR2XL U555 ( .A(n717), .B(n716), .Y(n432) );
  ADDFX2 U556 ( .A(n723), .B(n722), .CI(n721), .CO(n749), .S(n760) );
  OAI2BB1XL U557 ( .A0N(n1037), .A1N(n931), .B0(n428), .Y(n721) );
  OAI22XL U558 ( .A0(n939), .A1(n719), .B0(n937), .B1(n427), .Y(n722) );
  OAI22XL U559 ( .A0(n8), .A1(n718), .B0(n6), .B1(n426), .Y(n723) );
  AND2XL U560 ( .A(n928), .B(n42), .Y(n901) );
  CMPR32X1 U561 ( .A(n900), .B(n899), .C(n898), .CO(n909), .S(n952) );
  OAI22XL U562 ( .A0(n942), .A1(n897), .B0(n654), .B1(n856), .Y(n898) );
  OAI22XL U563 ( .A0(n939), .A1(n895), .B0(n937), .B1(n854), .Y(n899) );
  OAI22XL U564 ( .A0(n8), .A1(n893), .B0(n6), .B1(n852), .Y(n900) );
  NAND2BXL U565 ( .AN(n934), .B(n38), .Y(n37) );
  OAI22XL U566 ( .A0(n939), .A1(n537), .B0(n937), .B1(n938), .Y(n977) );
  OAI22XL U567 ( .A0(n8), .A1(n536), .B0(n6), .B1(n935), .Y(n979) );
  OAI22XL U568 ( .A0(n7), .A1(n546), .B0(n918), .B1(n566), .Y(n559) );
  INVXL U569 ( .A(n1116), .Y(n231) );
  OAI22XL U570 ( .A0(n1161), .A1(n215), .B0(n1162), .B1(n230), .Y(n233) );
  OAI22XL U571 ( .A0(n1139), .A1(n216), .B0(n9), .B1(n229), .Y(n236) );
  OAI22XL U572 ( .A0(n1139), .A1(n268), .B0(n9), .B1(n257), .Y(n274) );
  XNOR2XL U573 ( .A(n1156), .B(n894), .Y(n258) );
  OAI22XL U574 ( .A0(n8), .A1(n292), .B0(n6), .B1(n287), .Y(n301) );
  OAI22XL U575 ( .A0(n1161), .A1(n1131), .B0(n1162), .B1(n1147), .Y(n1144) );
  XOR2X1 U576 ( .A(n40), .B(n629), .Y(n660) );
  XNOR2X1 U577 ( .A(n630), .B(n41), .Y(n40) );
  NAND2XL U578 ( .A(n1110), .B(n1109), .Y(n1111) );
  CMPR32X1 U579 ( .A(n743), .B(n742), .C(n741), .CO(n703), .S(n744) );
  ADDFX2 U580 ( .A(n749), .B(n748), .CI(n747), .CO(n743), .S(n770) );
  NAND2X1 U581 ( .A(n44), .B(n43), .Y(n626) );
  OAI21XL U582 ( .A0(n630), .A1(n631), .B0(n629), .Y(n44) );
  NOR2XL U583 ( .A(n1152), .B(n1151), .Y(mult_x_1_n109) );
  NAND2XL U584 ( .A(n1227), .B(n1226), .Y(n1229) );
  INVXL U585 ( .A(n1225), .Y(n1227) );
  NAND2XL U586 ( .A(n409), .B(n408), .Y(mult_x_1_n184) );
  NOR2XL U587 ( .A(n1108), .B(n1107), .Y(mult_x_1_n136) );
  INVXL U588 ( .A(n1111), .Y(mult_x_1_n305) );
  NAND2XL U589 ( .A(n1169), .B(n1168), .Y(mult_x_1_n58) );
  NAND2XL U590 ( .A(n1167), .B(n1166), .Y(n1168) );
  NAND2XL U591 ( .A(n1152), .B(n1151), .Y(mult_x_1_n110) );
  NOR2XL U592 ( .A(n1141), .B(n1140), .Y(mult_x_1_n120) );
  NAND2XL U593 ( .A(n1141), .B(n1140), .Y(mult_x_1_n121) );
  NOR2XL U594 ( .A(n1127), .B(n1126), .Y(mult_x_1_n129) );
  NAND2XL U595 ( .A(n1127), .B(n1126), .Y(mult_x_1_n130) );
  NAND2XL U596 ( .A(n1317), .B(n1111), .Y(mult_x_1_n84) );
  NAND2X1 U597 ( .A(n993), .B(n994), .Y(n39) );
  OAI21XL U598 ( .A0(n993), .A1(n994), .B0(n992), .Y(n26) );
  NAND2X1 U599 ( .A(n58), .B(n57), .Y(n1020) );
  NAND2X1 U600 ( .A(n1029), .B(n1030), .Y(n57) );
  NAND2XL U601 ( .A(n1234), .B(n1233), .Y(n1236) );
  NAND2XL U602 ( .A(n1254), .B(n1253), .Y(n1256) );
  INVXL U603 ( .A(n1252), .Y(n1254) );
  NAND2XL U604 ( .A(n1196), .B(n1195), .Y(n1197) );
  NOR2BXL U605 ( .AN(n1038), .B(n1037), .Y(n1341) );
  NAND2XL U606 ( .A(n104), .B(n1230), .Y(n1232) );
  NAND2XL U607 ( .A(n1201), .B(n1200), .Y(n1203) );
  INVXL U608 ( .A(n1199), .Y(n1201) );
  NAND2XL U609 ( .A(n1190), .B(n1189), .Y(n1191) );
  XNOR2X1 U610 ( .A(B[6]), .B(B[5]), .Y(n64) );
  CLKINVX3 U611 ( .A(B[13]), .Y(n594) );
  NOR2X2 U612 ( .A(n1307), .B(n1308), .Y(n497) );
  BUFX3 U613 ( .A(B[3]), .Y(n68) );
  NOR2X1 U614 ( .A(n1299), .B(n1300), .Y(n448) );
  NAND2X1 U615 ( .A(n243), .B(n484), .Y(n446) );
  OAI21XL U616 ( .A0(n473), .A1(n480), .B0(n474), .Y(n450) );
  OR2X2 U617 ( .A(n1096), .B(n1095), .Y(n24) );
  OAI22X1 U618 ( .A0(n7), .A1(n260), .B0(n918), .B1(n63), .Y(n127) );
  CMPR22X1 U619 ( .A(n779), .B(n778), .CO(n756), .S(n790) );
  CMPR22X1 U620 ( .A(n847), .B(n846), .CO(n822), .S(n861) );
  CMPR22X1 U621 ( .A(n976), .B(n975), .CO(n983), .S(n1005) );
  OAI22X1 U622 ( .A0(n169), .A1(n133), .B0(n168), .B1(n1037), .Y(n167) );
  NAND2X1 U623 ( .A(B[1]), .B(n780), .Y(n169) );
  CMPR22X1 U624 ( .A(n726), .B(n725), .CO(n739), .S(n757) );
  CMPR22X1 U625 ( .A(n87), .B(n86), .CO(n81), .S(n108) );
  CMPR22X1 U626 ( .A(n644), .B(n643), .CO(n640), .S(n1059) );
  OAI22X1 U627 ( .A0(n1139), .A1(n594), .B0(n9), .B1(n593), .Y(n643) );
  OAI22X1 U628 ( .A0(n212), .A1(n266), .B0(n845), .B1(n213), .Y(n221) );
  CMPR22X1 U629 ( .A(n103), .B(n102), .CO(n105), .S(n97) );
  OAI22X1 U630 ( .A0(n618), .A1(n94), .B0(n937), .B1(n101), .Y(n102) );
  CMPR22X1 U631 ( .A(n670), .B(n669), .CO(n1070), .S(n680) );
  OAI22X1 U632 ( .A0(n7), .A1(n960), .B0(n918), .B1(n917), .Y(n968) );
  NAND2X1 U633 ( .A(n510), .B(n509), .Y(n511) );
  XNOR2X2 U634 ( .A(n505), .B(n504), .Y(PRODUCT[22]) );
  ADDFX2 U635 ( .A(n191), .B(n190), .CI(n189), .CO(n676), .S(n187) );
  XOR3X2 U636 ( .A(n944), .B(n36), .C(n943), .Y(n990) );
  OAI21XL U637 ( .A0(n614), .A1(n615), .B0(n48), .Y(n45) );
  XOR2X1 U638 ( .A(n42), .B(n928), .Y(n946) );
  INVX8 U639 ( .A(n260), .Y(n837) );
  XOR2X1 U640 ( .A(B[9]), .B(B[8]), .Y(n122) );
  AOI21X2 U641 ( .A0(n486), .A1(n243), .B0(n27), .Y(n479) );
  NOR2X2 U642 ( .A(n497), .B(n491), .Y(n243) );
  NOR2X2 U643 ( .A(n1305), .B(n1306), .Y(n491) );
  OAI21X2 U644 ( .A0(n501), .A1(n1044), .B0(n502), .Y(n486) );
  NOR2X4 U645 ( .A(n1309), .B(n1310), .Y(n501) );
  OAI21X4 U646 ( .A0(n241), .A1(n242), .B0(n28), .Y(n449) );
  XOR2X1 U647 ( .A(n1289), .B(n30), .Y(PRODUCT[15]) );
  AOI21X1 U648 ( .A0(n1259), .A1(n1293), .B0(n1260), .Y(n30) );
  NAND2X1 U649 ( .A(n33), .B(n32), .Y(n1018) );
  XOR3X2 U650 ( .A(n1014), .B(n31), .C(n1013), .Y(n1028) );
  OAI21XL U651 ( .A0(n944), .A1(n36), .B0(n943), .Y(n35) );
  XOR3X2 U652 ( .A(n992), .B(n994), .C(n993), .Y(n995) );
  INVXL U653 ( .A(n614), .Y(n46) );
  XOR3X2 U654 ( .A(n614), .B(n615), .C(n48), .Y(n1088) );
  INVXL U655 ( .A(n54), .Y(n52) );
  XOR2X1 U656 ( .A(n967), .B(n53), .Y(n987) );
  XOR2X1 U657 ( .A(n968), .B(n54), .Y(n53) );
  OAI21XL U658 ( .A0(n1018), .A1(n1016), .B0(n1017), .Y(n55) );
  XOR2X1 U659 ( .A(n1016), .B(n1018), .Y(n56) );
  XOR3X2 U660 ( .A(n1030), .B(n1028), .C(n1029), .Y(n1031) );
  NOR2X1 U661 ( .A(n203), .B(n202), .Y(n663) );
  CMPR22X1 U662 ( .A(n167), .B(n166), .CO(n188), .S(n164) );
  NOR2X1 U663 ( .A(n178), .B(n177), .Y(n692) );
  BUFX3 U664 ( .A(n130), .Y(n845) );
  AOI21XL U665 ( .A0(n666), .A1(n665), .B0(n664), .Y(n1082) );
  CMPR22X1 U666 ( .A(n576), .B(n575), .CO(n582), .S(n612) );
  NOR2X2 U667 ( .A(n1313), .B(n1314), .Y(n508) );
  NOR2X2 U668 ( .A(n1315), .B(n1316), .Y(n506) );
  NAND2X2 U669 ( .A(n1303), .B(n1304), .Y(n480) );
  NAND2X1 U670 ( .A(n379), .B(n252), .Y(n1239) );
  OAI22X1 U671 ( .A0(n8), .A1(n185), .B0(n6), .B1(n184), .Y(n669) );
  XNOR2X1 U672 ( .A(B[4]), .B(B[3]), .Y(n74) );
  XNOR2XL U673 ( .A(n817), .B(n932), .Y(n126) );
  XNOR2XL U674 ( .A(n888), .B(n1119), .Y(n849) );
  XNOR2XL U675 ( .A(n888), .B(n853), .Y(n930) );
  XNOR2XL U676 ( .A(n1156), .B(n853), .Y(n211) );
  XNOR2XL U677 ( .A(n817), .B(n578), .Y(n84) );
  BUFX3 U678 ( .A(B[16]), .Y(n1156) );
  XNOR2XL U679 ( .A(n1156), .B(n848), .Y(n226) );
  XNOR2XL U680 ( .A(n817), .B(n1135), .Y(n706) );
  XNOR2XL U681 ( .A(n1156), .B(n887), .Y(n210) );
  XNOR2XL U682 ( .A(n1156), .B(n1145), .Y(n1146) );
  OAI22X1 U683 ( .A0(n1161), .A1(n920), .B0(n1162), .B1(n877), .Y(n924) );
  OAI22X1 U684 ( .A0(n1161), .A1(n526), .B0(n1162), .B1(n521), .Y(n556) );
  ADDFX2 U685 ( .A(n991), .B(n990), .CI(n989), .CO(n994), .S(n1016) );
  INVX1 U686 ( .A(B[0]), .Y(n780) );
  INVX1 U687 ( .A(B[1]), .Y(n519) );
  XNOR2X1 U688 ( .A(B[1]), .B(A[6]), .Y(n65) );
  XNOR2X1 U689 ( .A(n888), .B(n921), .Y(n134) );
  BUFX3 U690 ( .A(n780), .Y(n1037) );
  OAI22X1 U691 ( .A0(n169), .A1(n65), .B0(n134), .B1(n1037), .Y(n128) );
  XOR2X1 U692 ( .A(B[6]), .B(B[7]), .Y(n62) );
  BUFX3 U693 ( .A(n64), .Y(n918) );
  BUFX3 U694 ( .A(A[0]), .Y(n1038) );
  NOR2BX1 U695 ( .AN(n1038), .B(n918), .Y(n79) );
  BUFX3 U696 ( .A(n169), .Y(n931) );
  OAI22X2 U697 ( .A0(n931), .A1(n73), .B0(n65), .B1(n1037), .Y(n78) );
  XOR2X1 U698 ( .A(B[4]), .B(B[5]), .Y(n66) );
  BUFX4 U699 ( .A(B[5]), .Y(n817) );
  BUFX3 U700 ( .A(n74), .Y(n654) );
  OAI22X1 U701 ( .A0(n942), .A1(n84), .B0(n654), .B1(n71), .Y(n77) );
  XOR2XL U702 ( .A(B[2]), .B(B[3]), .Y(n67) );
  XNOR2X1 U703 ( .A(B[2]), .B(B[1]), .Y(n586) );
  XNOR2X1 U704 ( .A(n68), .B(n919), .Y(n124) );
  OAI22X1 U705 ( .A0(n939), .A1(n72), .B0(n937), .B1(n124), .Y(n142) );
  XNOR2X1 U706 ( .A(n837), .B(n578), .Y(n136) );
  OAI22X1 U707 ( .A0(n939), .A1(n83), .B0(n586), .B1(n72), .Y(n82) );
  XNOR2X1 U708 ( .A(n888), .B(n890), .Y(n98) );
  OAI22X1 U709 ( .A0(n931), .A1(n98), .B0(n73), .B1(n1037), .Y(n87) );
  OAI22X1 U710 ( .A0(n942), .A1(n76), .B0(n654), .B1(n75), .Y(n86) );
  NOR2XL U711 ( .A(n1194), .B(n1199), .Y(n121) );
  XNOR2X1 U712 ( .A(B[1]), .B(n578), .Y(n88) );
  XNOR2X1 U713 ( .A(B[1]), .B(n638), .Y(n93) );
  OR2X2 U714 ( .A(n91), .B(n90), .Y(n1234) );
  OAI22X1 U715 ( .A0(n931), .A1(n93), .B0(n99), .B1(n1037), .Y(n103) );
  XNOR2X1 U716 ( .A(n68), .B(n1038), .Y(n94) );
  XNOR2XL U717 ( .A(n68), .B(n578), .Y(n101) );
  NOR2XL U718 ( .A(n97), .B(n96), .Y(n1225) );
  OAI21XL U719 ( .A0(n1228), .A1(n1225), .B0(n1226), .Y(n1231) );
  AOI21XL U720 ( .A0(n1231), .A1(n104), .B0(n107), .Y(n1255) );
  CMPR32X1 U721 ( .A(n110), .B(n109), .C(n108), .CO(n116), .S(n115) );
  CMPR32X1 U722 ( .A(n113), .B(n112), .C(n111), .CO(n114), .S(n106) );
  OAI21XL U723 ( .A0(n1255), .A1(n1252), .B0(n1253), .Y(n1193) );
  NAND2X1 U724 ( .A(n117), .B(n116), .Y(n1200) );
  NAND2XL U725 ( .A(n119), .B(n118), .Y(n1195) );
  OAI21XL U726 ( .A0(n1194), .A1(n1200), .B0(n1195), .Y(n120) );
  XNOR2X1 U727 ( .A(B[8]), .B(B[7]), .Y(n130) );
  NAND2X1 U728 ( .A(n122), .B(n130), .Y(n212) );
  XNOR2X1 U729 ( .A(n712), .B(n1038), .Y(n123) );
  BUFX3 U730 ( .A(n130), .Y(n970) );
  XNOR2X1 U731 ( .A(n712), .B(n578), .Y(n170) );
  OAI22X1 U732 ( .A0(n972), .A1(n123), .B0(n970), .B1(n170), .Y(n172) );
  XNOR2X1 U733 ( .A(n817), .B(n890), .Y(n125) );
  XNOR2X1 U734 ( .A(n68), .B(n921), .Y(n162) );
  XNOR2XL U735 ( .A(n888), .B(n878), .Y(n133) );
  XNOR2XL U736 ( .A(B[1]), .B(n892), .Y(n168) );
  NAND2BX1 U737 ( .AN(n1038), .B(n712), .Y(n131) );
  OAI22X2 U738 ( .A0(n212), .A1(n132), .B0(n845), .B1(n131), .Y(n166) );
  OAI22X1 U739 ( .A0(n169), .A1(n134), .B0(n133), .B1(n1037), .Y(n138) );
  ADDFHX1 U740 ( .A(n139), .B(n138), .CI(n137), .CO(n163), .S(n148) );
  OR2X2 U741 ( .A(n155), .B(n154), .Y(n700) );
  CMPR32X1 U742 ( .A(n148), .B(n147), .C(n146), .CO(n154), .S(n153) );
  OR2X2 U743 ( .A(n153), .B(n152), .Y(n1190) );
  NAND2XL U744 ( .A(n153), .B(n152), .Y(n1189) );
  INVXL U745 ( .A(n1189), .Y(n698) );
  NAND2XL U746 ( .A(n155), .B(n154), .Y(n699) );
  INVXL U747 ( .A(n699), .Y(n156) );
  XNOR2X1 U748 ( .A(n68), .B(n878), .Y(n198) );
  CMPR32X1 U749 ( .A(n165), .B(n164), .C(n163), .CO(n200), .S(n174) );
  XNOR2X1 U750 ( .A(B[10]), .B(B[9]), .Y(n183) );
  NOR2BX1 U751 ( .AN(n1038), .B(n6), .Y(n191) );
  XNOR2XL U752 ( .A(B[1]), .B(n851), .Y(n181) );
  XNOR2X1 U753 ( .A(n712), .B(n638), .Y(n180) );
  NAND2XL U754 ( .A(n178), .B(n177), .Y(n693) );
  OAI21XL U755 ( .A0(n696), .A1(n692), .B0(n693), .Y(n206) );
  XNOR2X1 U756 ( .A(n712), .B(n932), .Y(n668) );
  OAI22X1 U757 ( .A0(n931), .A1(n181), .B0(n646), .B1(n1037), .Y(n670) );
  XOR2X1 U758 ( .A(B[10]), .B(B[11]), .Y(n182) );
  NAND2XL U759 ( .A(n182), .B(n183), .Y(n196) );
  CMPR32X1 U760 ( .A(n194), .B(n193), .C(n192), .CO(n675), .S(n201) );
  OAI22X1 U761 ( .A0(n7), .A1(n195), .B0(n918), .B1(n650), .Y(n679) );
  OAI22X1 U762 ( .A0(n8), .A1(n197), .B0(n6), .B1(n648), .Y(n678) );
  XNOR2X1 U763 ( .A(n68), .B(n892), .Y(n652) );
  CMPR32X1 U764 ( .A(n201), .B(n200), .C(n199), .CO(n202), .S(n178) );
  INVXL U765 ( .A(n663), .Y(n204) );
  NAND2XL U766 ( .A(n203), .B(n202), .Y(n662) );
  NAND2XL U767 ( .A(n204), .B(n662), .Y(n205) );
  XNOR2X1 U768 ( .A(n206), .B(n205), .Y(n1330) );
  NOR2X1 U769 ( .A(n1283), .B(n1285), .Y(n237) );
  INVXL U770 ( .A(n506), .Y(n207) );
  NAND2X1 U771 ( .A(n1315), .B(n1316), .Y(n238) );
  NAND2XL U772 ( .A(n207), .B(n238), .Y(n208) );
  XNOR2X1 U773 ( .A(n209), .B(n848), .Y(n215) );
  BUFX3 U774 ( .A(n328), .Y(n1158) );
  XNOR2XL U775 ( .A(n286), .B(A[24]), .Y(n217) );
  XNOR2XL U776 ( .A(B[11]), .B(A[25]), .Y(n227) );
  OAI22X1 U777 ( .A0(n8), .A1(n217), .B0(n6), .B1(n227), .Y(n1116) );
  CLKINVX3 U778 ( .A(n594), .Y(n362) );
  XNOR2XL U779 ( .A(n362), .B(n1135), .Y(n216) );
  XNOR2X1 U780 ( .A(n362), .B(n1145), .Y(n229) );
  XNOR2XL U781 ( .A(n712), .B(A[24]), .Y(n266) );
  XNOR2X1 U782 ( .A(n712), .B(A[25]), .Y(n213) );
  XNOR2X1 U783 ( .A(n209), .B(n887), .Y(n218) );
  XNOR2X1 U784 ( .A(n362), .B(n1119), .Y(n257) );
  OAI22XL U785 ( .A0(n1139), .A1(n257), .B0(n9), .B1(n216), .Y(n224) );
  XNOR2XL U786 ( .A(n286), .B(n1145), .Y(n219) );
  XNOR2X1 U787 ( .A(n209), .B(n853), .Y(n267) );
  OAI22XL U788 ( .A0(n1161), .A1(n267), .B0(n1162), .B1(n218), .Y(n271) );
  XNOR2X1 U789 ( .A(B[11]), .B(n1135), .Y(n287) );
  OAI22XL U790 ( .A0(n8), .A1(n287), .B0(n6), .B1(n219), .Y(n270) );
  CMPR32X1 U791 ( .A(n222), .B(n221), .C(n220), .CO(n235), .S(n264) );
  CMPR32X1 U792 ( .A(n225), .B(n224), .C(n223), .CO(n234), .S(n263) );
  XNOR2XL U793 ( .A(n362), .B(A[24]), .Y(n1122) );
  OAI22XL U794 ( .A0(n1139), .A1(n229), .B0(n9), .B1(n1122), .Y(n1125) );
  XNOR2X1 U795 ( .A(n209), .B(n1135), .Y(n1118) );
  CMPR32X1 U796 ( .A(n233), .B(n232), .C(n231), .CO(n1123), .S(n277) );
  CMPR32X1 U797 ( .A(n236), .B(n235), .C(n234), .CO(n1112), .S(n276) );
  NAND2XL U798 ( .A(n1108), .B(n1107), .Y(mult_x_1_n137) );
  NOR2X1 U799 ( .A(n1303), .B(n1304), .Y(n468) );
  NOR2X1 U800 ( .A(n448), .B(n455), .Y(n245) );
  NAND2X1 U801 ( .A(n447), .B(n245), .Y(n247) );
  NOR2XL U802 ( .A(n446), .B(n247), .Y(n249) );
  NAND2X1 U803 ( .A(n1313), .B(n1314), .Y(n509) );
  NAND2X1 U804 ( .A(n1305), .B(n1306), .Y(n492) );
  OAI21XL U805 ( .A0(n455), .A1(n464), .B0(n456), .Y(n244) );
  AOI21XL U806 ( .A0(n245), .A1(n450), .B0(n244), .Y(n246) );
  OAI21X1 U807 ( .A0(n479), .A1(n247), .B0(n246), .Y(n248) );
  AOI21X2 U808 ( .A0(n249), .A1(n449), .B0(n248), .Y(n250) );
  BUFX8 U809 ( .A(n250), .Y(n1250) );
  NOR2X1 U810 ( .A(n1296), .B(n1295), .Y(n1039) );
  NOR2XL U811 ( .A(n1039), .B(n1281), .Y(n379) );
  NOR2XL U812 ( .A(n1239), .B(n1275), .Y(n280) );
  NAND2XL U813 ( .A(n280), .B(n1170), .Y(n254) );
  NAND2X1 U814 ( .A(n1296), .B(n1295), .Y(n1040) );
  OAI21XL U815 ( .A0(n1277), .A1(n1280), .B0(n1278), .Y(n251) );
  OAI21XL U816 ( .A0(n1246), .A1(n1275), .B0(n1276), .Y(n281) );
  AOI21XL U817 ( .A0(n281), .A1(n1170), .B0(n1173), .Y(n253) );
  XNOR2X1 U818 ( .A(n362), .B(n848), .Y(n268) );
  NOR2X1 U819 ( .A(n1158), .B(n259), .Y(n298) );
  XNOR2XL U820 ( .A(n837), .B(A[24]), .Y(n322) );
  XNOR2XL U821 ( .A(n837), .B(A[25]), .Y(n261) );
  OAI22X1 U822 ( .A0(n7), .A1(n322), .B0(n918), .B1(n261), .Y(n297) );
  CMPR32X1 U823 ( .A(n265), .B(n264), .C(n263), .CO(n275), .S(n306) );
  XNOR2X1 U824 ( .A(n712), .B(n1145), .Y(n289) );
  XNOR2X1 U825 ( .A(n209), .B(n894), .Y(n291) );
  OAI22XL U826 ( .A0(n1161), .A1(n291), .B0(n1162), .B1(n267), .Y(n294) );
  XNOR2X1 U827 ( .A(n362), .B(n887), .Y(n288) );
  CMPR32X1 U828 ( .A(n271), .B(n270), .C(n269), .CO(n265), .S(n303) );
  CMPR32X1 U829 ( .A(n274), .B(n273), .C(n272), .CO(n307), .S(n302) );
  CMPR32X1 U830 ( .A(n277), .B(n276), .C(n275), .CO(n1108), .S(n278) );
  NOR2XL U831 ( .A(n279), .B(n278), .Y(mult_x_1_n151) );
  NAND2XL U832 ( .A(n279), .B(n278), .Y(mult_x_1_n152) );
  INVXL U833 ( .A(n280), .Y(n283) );
  INVXL U834 ( .A(n281), .Y(n282) );
  OAI21XL U835 ( .A0(n1250), .A1(n283), .B0(n282), .Y(n285) );
  XNOR2X1 U836 ( .A(n285), .B(n284), .Y(PRODUCT[34]) );
  XNOR2X1 U837 ( .A(n362), .B(n853), .Y(n326) );
  XNOR2X1 U838 ( .A(n712), .B(n1135), .Y(n324) );
  XNOR2X1 U839 ( .A(n209), .B(n855), .Y(n323) );
  XNOR2X1 U840 ( .A(n286), .B(n848), .Y(n325) );
  CMPR32X1 U841 ( .A(n295), .B(n294), .C(n293), .CO(n304), .S(n341) );
  CMPR32X1 U842 ( .A(n298), .B(n297), .C(n296), .CO(n272), .S(n340) );
  CMPR32X1 U843 ( .A(n304), .B(n303), .C(n302), .CO(n305), .S(n342) );
  CMPR32X1 U844 ( .A(n307), .B(n306), .C(n305), .CO(n279), .S(n308) );
  NOR2XL U845 ( .A(n309), .B(n308), .Y(mult_x_1_n160) );
  NAND2XL U846 ( .A(n309), .B(n308), .Y(mult_x_1_n161) );
  OAI21X1 U847 ( .A0(n1250), .A1(n1239), .B0(n1246), .Y(n312) );
  XNOR2XL U848 ( .A(n817), .B(A[24]), .Y(n358) );
  XNOR2XL U849 ( .A(n817), .B(A[25]), .Y(n314) );
  OAI22X1 U850 ( .A0(n942), .A1(n358), .B0(n654), .B1(n314), .Y(n334) );
  XNOR2X1 U851 ( .A(B[11]), .B(n887), .Y(n332) );
  XNOR2X1 U852 ( .A(n362), .B(n894), .Y(n327) );
  OAI22XL U853 ( .A0(n1139), .A1(n327), .B0(n9), .B1(n326), .Y(n351) );
  XNOR2X1 U854 ( .A(n362), .B(n855), .Y(n363) );
  NOR2XL U855 ( .A(n328), .B(n329), .Y(n366) );
  XNOR2X1 U856 ( .A(n837), .B(n1135), .Y(n360) );
  XNOR2X1 U857 ( .A(n209), .B(n875), .Y(n359) );
  OAI22X1 U858 ( .A0(n1161), .A1(n359), .B0(n1162), .B1(n331), .Y(n369) );
  XNOR2XL U859 ( .A(n286), .B(n853), .Y(n364) );
  CMPR32X1 U860 ( .A(n338), .B(n337), .C(n336), .CO(n373), .S(n386) );
  CMPR32X1 U861 ( .A(n341), .B(n340), .C(n339), .CO(n343), .S(n374) );
  CMPR32X1 U862 ( .A(n344), .B(n343), .C(n342), .CO(n309), .S(n345) );
  NOR2XL U863 ( .A(n346), .B(n345), .Y(mult_x_1_n169) );
  NAND2XL U864 ( .A(n346), .B(n345), .Y(mult_x_1_n170) );
  CMPR32X1 U865 ( .A(n349), .B(n348), .C(n347), .CO(n376), .S(n385) );
  CMPR32X1 U866 ( .A(n352), .B(n351), .C(n350), .CO(n372), .S(n391) );
  XNOR2X1 U867 ( .A(n712), .B(n848), .Y(n361) );
  XNOR2XL U868 ( .A(n68), .B(A[24]), .Y(n427) );
  XNOR2X1 U869 ( .A(n68), .B(A[25]), .Y(n356) );
  OAI22X2 U870 ( .A0(n939), .A1(n427), .B0(n937), .B1(n356), .Y(n416) );
  OAI22X1 U871 ( .A0(n942), .A1(n414), .B0(n654), .B1(n358), .Y(n401) );
  XNOR2X1 U872 ( .A(n209), .B(n916), .Y(n398) );
  XNOR2X1 U873 ( .A(n837), .B(n1119), .Y(n395) );
  XNOR2X1 U874 ( .A(n712), .B(n887), .Y(n418) );
  XNOR2X1 U875 ( .A(n286), .B(n894), .Y(n419) );
  OAI22XL U876 ( .A0(n8), .A1(n419), .B0(n6), .B1(n364), .Y(n402) );
  CMPR32X1 U877 ( .A(n370), .B(n369), .C(n368), .CO(n388), .S(n405) );
  CMPR32X1 U878 ( .A(n376), .B(n375), .C(n374), .CO(n346), .S(n377) );
  NOR2XL U879 ( .A(n378), .B(n377), .Y(mult_x_1_n176) );
  NAND2XL U880 ( .A(n378), .B(n377), .Y(mult_x_1_n177) );
  INVXL U881 ( .A(n380), .Y(n1049) );
  XNOR2X2 U882 ( .A(n382), .B(n381), .Y(PRODUCT[31]) );
  ADDFHX1 U883 ( .A(n385), .B(n384), .CI(n383), .CO(n378), .S(n409) );
  CMPR32X1 U884 ( .A(n391), .B(n390), .C(n389), .CO(n384), .S(n442) );
  CMPR32X1 U885 ( .A(n394), .B(n393), .C(n392), .CO(n390), .S(n425) );
  XNOR2X1 U886 ( .A(B[16]), .B(n926), .Y(n396) );
  XNOR2X1 U887 ( .A(n209), .B(n883), .Y(n421) );
  OAI22XL U888 ( .A0(n422), .A1(n421), .B0(n1162), .B1(n398), .Y(n709) );
  CMPR32X1 U889 ( .A(n404), .B(n403), .C(n402), .CO(n407), .S(n435) );
  CMPR32X1 U890 ( .A(n407), .B(n406), .C(n405), .CO(n389), .S(n423) );
  NOR2XL U891 ( .A(n409), .B(n408), .Y(mult_x_1_n183) );
  OAI21X2 U892 ( .A0(n1250), .A1(n1039), .B0(n1040), .Y(n412) );
  INVXL U893 ( .A(n1281), .Y(n410) );
  NAND2X1 U894 ( .A(n410), .B(n1282), .Y(n411) );
  XNOR2X2 U895 ( .A(n412), .B(n411), .Y(PRODUCT[30]) );
  CLKINVX3 U896 ( .A(n594), .Y(n1121) );
  XNOR2X1 U897 ( .A(n1121), .B(n875), .Y(n708) );
  OAI22XL U898 ( .A0(n1139), .A1(n708), .B0(n9), .B1(n413), .Y(n431) );
  ADDFHX1 U899 ( .A(n417), .B(n416), .CI(n415), .CO(n393), .S(n439) );
  XNOR2XL U900 ( .A(n712), .B(n853), .Y(n713) );
  XNOR2X1 U901 ( .A(n286), .B(n855), .Y(n426) );
  XNOR2X1 U902 ( .A(n209), .B(n926), .Y(n733) );
  CMPR32X1 U903 ( .A(n431), .B(n430), .C(n429), .CO(n440), .S(n748) );
  CMPR32X1 U904 ( .A(n434), .B(n433), .C(n432), .CO(n438), .S(n747) );
  CMPR32X1 U905 ( .A(n440), .B(n439), .C(n438), .CO(n705), .S(n741) );
  ADDFHX1 U906 ( .A(n443), .B(n442), .CI(n441), .CO(n408), .S(n444) );
  NOR2XL U907 ( .A(n445), .B(n444), .Y(mult_x_1_n194) );
  NAND2XL U908 ( .A(n445), .B(n444), .Y(mult_x_1_n195) );
  INVXL U909 ( .A(n446), .Y(n478) );
  INVXL U910 ( .A(n447), .Y(n460) );
  NAND2XL U911 ( .A(n478), .B(n452), .Y(n454) );
  INVX1 U912 ( .A(n479), .Y(n470) );
  INVXL U913 ( .A(n450), .Y(n461) );
  OAI21XL U914 ( .A0(n461), .A1(n448), .B0(n464), .Y(n451) );
  INVXL U915 ( .A(n455), .Y(n457) );
  NAND2XL U916 ( .A(n478), .B(n447), .Y(n463) );
  OAI21XL U917 ( .A0(n1047), .A1(n463), .B0(n462), .Y(n467) );
  NAND2XL U918 ( .A(n478), .B(n481), .Y(n472) );
  OAI21XL U919 ( .A0(n1047), .A1(n446), .B0(n479), .Y(n483) );
  XNOR2X1 U920 ( .A(n483), .B(n482), .Y(PRODUCT[25]) );
  INVXL U921 ( .A(n497), .Y(n488) );
  NAND2XL U922 ( .A(n484), .B(n488), .Y(n490) );
  INVXL U923 ( .A(n498), .Y(n487) );
  OAI21XL U924 ( .A0(n1047), .A1(n490), .B0(n489), .Y(n495) );
  NAND2XL U925 ( .A(n493), .B(n492), .Y(n494) );
  NAND2XL U926 ( .A(n488), .B(n498), .Y(n499) );
  INVXL U927 ( .A(n508), .Y(n510) );
  XNOR2X2 U928 ( .A(n512), .B(n511), .Y(PRODUCT[20]) );
  INVXL U929 ( .A(n1283), .Y(n514) );
  XNOR2X1 U930 ( .A(n209), .B(n638), .Y(n526) );
  XNOR2X1 U931 ( .A(n209), .B(n932), .Y(n521) );
  NOR2XL U932 ( .A(n328), .B(n517), .Y(n555) );
  OAI22XL U933 ( .A0(n1139), .A1(n534), .B0(n9), .B1(n565), .Y(n554) );
  XNOR2X1 U934 ( .A(n837), .B(n926), .Y(n566) );
  XNOR2X1 U935 ( .A(n712), .B(n878), .Y(n532) );
  XNOR2X1 U936 ( .A(n712), .B(n892), .Y(n563) );
  OAI22XL U937 ( .A0(n972), .A1(n532), .B0(n970), .B1(n563), .Y(n558) );
  CLKINVX3 U938 ( .A(n519), .Y(n888) );
  XNOR2X1 U939 ( .A(n888), .B(n855), .Y(n524) );
  XNOR2X1 U940 ( .A(n286), .B(n921), .Y(n536) );
  XNOR2X1 U941 ( .A(n286), .B(n878), .Y(n935) );
  OAI22X1 U942 ( .A0(n1161), .A1(n521), .B0(n1162), .B1(n963), .Y(n978) );
  XNOR2X1 U943 ( .A(n68), .B(n896), .Y(n537) );
  XNOR2X1 U944 ( .A(n68), .B(n855), .Y(n938) );
  XNOR2X1 U945 ( .A(n888), .B(n875), .Y(n577) );
  XNOR2X1 U946 ( .A(n888), .B(n896), .Y(n525) );
  OAI22X1 U947 ( .A0(n931), .A1(n577), .B0(n525), .B1(n1037), .Y(n576) );
  OAI22X2 U948 ( .A0(n1161), .A1(n523), .B0(n1162), .B1(n522), .Y(n575) );
  XNOR2X1 U949 ( .A(n712), .B(A[6]), .Y(n583) );
  XNOR2X1 U950 ( .A(n712), .B(n921), .Y(n533) );
  XNOR2X1 U951 ( .A(n209), .B(n1038), .Y(n528) );
  XNOR2X1 U952 ( .A(n1121), .B(n638), .Y(n579) );
  XNOR2X1 U953 ( .A(n1121), .B(n932), .Y(n535) );
  OAI22XL U954 ( .A0(n1139), .A1(n579), .B0(n9), .B1(n535), .Y(n587) );
  CMPR32X1 U955 ( .A(n531), .B(n530), .C(n529), .CO(n550), .S(n581) );
  OAI22X1 U956 ( .A0(n972), .A1(n533), .B0(n970), .B1(n532), .Y(n542) );
  XNOR2X1 U957 ( .A(n68), .B(n916), .Y(n539) );
  OAI22X2 U958 ( .A0(n939), .A1(n539), .B0(n937), .B1(n538), .Y(n541) );
  OAI22XL U959 ( .A0(n1139), .A1(n535), .B0(n9), .B1(n534), .Y(n540) );
  XNOR2X1 U960 ( .A(n68), .B(n883), .Y(n585) );
  XNOR2X1 U961 ( .A(n286), .B(n890), .Y(n584) );
  OAI22X1 U962 ( .A0(n8), .A1(n584), .B0(n6), .B1(n545), .Y(n609) );
  OAI22X1 U963 ( .A0(n8), .A1(n545), .B0(n6), .B1(n544), .Y(n552) );
  ADDFHX1 U964 ( .A(n550), .B(n549), .CI(n548), .CO(n1027), .S(n596) );
  CMPR32X1 U965 ( .A(n553), .B(n552), .C(n551), .CO(n573), .S(n605) );
  CMPR32X1 U966 ( .A(n556), .B(n555), .C(n554), .CO(n1024), .S(n572) );
  CMPR32X1 U967 ( .A(n559), .B(n558), .C(n557), .CO(n1023), .S(n571) );
  OAI22XL U968 ( .A0(n1139), .A1(n565), .B0(n9), .B1(n965), .Y(n998) );
  OAI22X1 U969 ( .A0(n931), .A1(n567), .B0(n930), .B1(n780), .Y(n976) );
  XNOR2XL U970 ( .A(B[16]), .B(n638), .Y(n568) );
  NOR2XL U971 ( .A(n328), .B(n568), .Y(n975) );
  ADDHXL U972 ( .A(n570), .B(n569), .CO(n1004), .S(n557) );
  XNOR2X1 U973 ( .A(B[1]), .B(n916), .Y(n592) );
  XNOR2X1 U974 ( .A(n1121), .B(n578), .Y(n636) );
  XNOR2X1 U975 ( .A(n286), .B(n932), .Y(n639) );
  OAI22X1 U976 ( .A0(n8), .A1(n639), .B0(n6), .B1(n584), .Y(n621) );
  XNOR2XL U977 ( .A(n68), .B(n926), .Y(n617) );
  XNOR2X1 U978 ( .A(n888), .B(n883), .Y(n645) );
  OAI22X1 U979 ( .A0(n931), .A1(n645), .B0(n592), .B1(n1037), .Y(n644) );
  ADDFHX1 U980 ( .A(n597), .B(n596), .CI(n595), .CO(n1035), .S(n602) );
  NOR2XL U981 ( .A(n599), .B(n598), .Y(mult_x_1_n281) );
  NAND2XL U982 ( .A(n599), .B(n598), .Y(mult_x_1_n282) );
  CMPR32X1 U983 ( .A(n604), .B(n603), .C(n602), .CO(n598), .S(n627) );
  CMPR32X1 U984 ( .A(n607), .B(n606), .C(n605), .CO(n595), .S(n631) );
  CMPR32X1 U985 ( .A(n610), .B(n609), .C(n608), .CO(n607), .S(n658) );
  CMPR32X1 U986 ( .A(n613), .B(n612), .C(n611), .CO(n625), .S(n657) );
  XNOR2X1 U987 ( .A(n712), .B(n890), .Y(n667) );
  OAI22XL U988 ( .A0(n618), .A1(n651), .B0(n937), .B1(n617), .Y(n1067) );
  CMPR32X1 U989 ( .A(n622), .B(n621), .C(n620), .CO(n634), .S(n1086) );
  NOR2XL U990 ( .A(n627), .B(n626), .Y(mult_x_1_n286) );
  NAND2XL U991 ( .A(n627), .B(n626), .Y(mult_x_1_n287) );
  ADDFHX1 U992 ( .A(n634), .B(n633), .CI(n632), .CO(n623), .S(n1085) );
  OAI22X1 U993 ( .A0(n7), .A1(n649), .B0(n918), .B1(n635), .Y(n1065) );
  XNOR2XL U994 ( .A(n1121), .B(n1038), .Y(n637) );
  OAI22X1 U995 ( .A0(n1139), .A1(n637), .B0(n9), .B1(n636), .Y(n1064) );
  XNOR2X1 U996 ( .A(n286), .B(n638), .Y(n647) );
  NOR2BX1 U997 ( .AN(n1038), .B(n9), .Y(n673) );
  OAI22X1 U998 ( .A0(n931), .A1(n646), .B0(n645), .B1(n1037), .Y(n672) );
  OAI22X1 U999 ( .A0(n8), .A1(n648), .B0(n6), .B1(n647), .Y(n671) );
  CMPR32X1 U1000 ( .A(n658), .B(n657), .C(n656), .CO(n630), .S(n1083) );
  NOR2XL U1001 ( .A(n660), .B(n659), .Y(mult_x_1_n292) );
  NAND2XL U1002 ( .A(n660), .B(n659), .Y(mult_x_1_n293) );
  XOR2X1 U1003 ( .A(n1294), .B(n1291), .Y(PRODUCT[13]) );
  XNOR2X1 U1004 ( .A(n1261), .B(n1292), .Y(PRODUCT[12]) );
  NOR2XL U1005 ( .A(n663), .B(n692), .Y(n665) );
  OAI21XL U1006 ( .A0(n663), .A1(n693), .B0(n662), .Y(n664) );
  INVXL U1007 ( .A(n1082), .Y(mult_x_1_n321) );
  OAI22XL U1008 ( .A0(n972), .A1(n668), .B0(n970), .B1(n667), .Y(n1071) );
  ADDFHX1 U1009 ( .A(n676), .B(n675), .CI(n674), .CO(n1073), .S(n686) );
  CMPR32X1 U1010 ( .A(n682), .B(n681), .C(n680), .CO(n1061), .S(n688) );
  CMPR32X1 U1011 ( .A(n685), .B(n684), .C(n683), .CO(n1057), .S(n1060) );
  CMPR32X1 U1012 ( .A(n688), .B(n687), .C(n686), .CO(n690), .S(n203) );
  INVXL U1013 ( .A(n1106), .Y(n1079) );
  AOI21XL U1014 ( .A0(mult_x_1_n321), .A1(n689), .B0(n1079), .Y(mult_x_1_n316)
         );
  INVXL U1015 ( .A(n692), .Y(n694) );
  NAND2XL U1016 ( .A(n694), .B(n693), .Y(n695) );
  XOR2X1 U1017 ( .A(n696), .B(n695), .Y(n1331) );
  INVXL U1018 ( .A(n697), .Y(n1192) );
  AOI21XL U1019 ( .A0(n1192), .A1(n1190), .B0(n698), .Y(n702) );
  NAND2XL U1020 ( .A(n700), .B(n699), .Y(n701) );
  XOR2X1 U1021 ( .A(n702), .B(n701), .Y(n1332) );
  XNOR2X1 U1022 ( .A(B[16]), .B(n851), .Y(n707) );
  NOR2XL U1023 ( .A(n328), .B(n707), .Y(n736) );
  XNOR2X1 U1024 ( .A(n1121), .B(n916), .Y(n734) );
  OAI22XL U1025 ( .A0(n1139), .A1(n734), .B0(n9), .B1(n708), .Y(n735) );
  XNOR2X1 U1026 ( .A(n712), .B(n894), .Y(n724) );
  OAI22XL U1027 ( .A0(n972), .A1(n724), .B0(n845), .B1(n713), .Y(n740) );
  OAI22X1 U1028 ( .A0(n931), .A1(n727), .B0(n714), .B1(n1037), .Y(n726) );
  XNOR2X1 U1029 ( .A(B[16]), .B(n892), .Y(n715) );
  NOR2XL U1030 ( .A(n328), .B(n715), .Y(n725) );
  XNOR2X1 U1031 ( .A(n717), .B(n716), .Y(n738) );
  XNOR2XL U1032 ( .A(n712), .B(n855), .Y(n777) );
  XNOR2X1 U1033 ( .A(n888), .B(n1145), .Y(n781) );
  OAI22X1 U1034 ( .A0(n931), .A1(n781), .B0(n727), .B1(n780), .Y(n779) );
  XNOR2XL U1035 ( .A(B[16]), .B(n878), .Y(n728) );
  NOR2XL U1036 ( .A(n328), .B(n728), .Y(n778) );
  CMPR32X1 U1037 ( .A(n731), .B(n730), .C(n729), .CO(n746), .S(n766) );
  OAI22X1 U1038 ( .A0(n7), .A1(n771), .B0(n918), .B1(n732), .Y(n776) );
  XNOR2X1 U1039 ( .A(n209), .B(n851), .Y(n772) );
  OAI22X1 U1040 ( .A0(n1161), .A1(n772), .B0(n1162), .B1(n733), .Y(n775) );
  XNOR2X1 U1041 ( .A(n1121), .B(n883), .Y(n773) );
  OAI22XL U1042 ( .A0(n1139), .A1(n773), .B0(n9), .B1(n734), .Y(n774) );
  CMPR32X1 U1043 ( .A(n737), .B(n736), .C(n735), .CO(n731), .S(n763) );
  CMPR32X1 U1044 ( .A(n740), .B(n739), .C(n738), .CO(n729), .S(n762) );
  CMPR32X1 U1045 ( .A(n758), .B(n757), .C(n756), .CO(n759), .S(n795) );
  CMPR32X1 U1046 ( .A(n764), .B(n763), .C(n762), .CO(n765), .S(n798) );
  OAI22X1 U1047 ( .A0(n7), .A1(n804), .B0(n918), .B1(n771), .Y(n809) );
  XNOR2X1 U1048 ( .A(n209), .B(n892), .Y(n805) );
  OAI22X1 U1049 ( .A0(n1161), .A1(n805), .B0(n1162), .B1(n772), .Y(n808) );
  XNOR2X1 U1050 ( .A(n1121), .B(n926), .Y(n806) );
  OAI22XL U1051 ( .A0(n1139), .A1(n806), .B0(n9), .B1(n773), .Y(n807) );
  XNOR2XL U1052 ( .A(n712), .B(n896), .Y(n810) );
  OAI22XL U1053 ( .A0(n972), .A1(n810), .B0(n845), .B1(n777), .Y(n791) );
  XNOR2X1 U1054 ( .A(n888), .B(n1135), .Y(n813) );
  XNOR2XL U1055 ( .A(B[16]), .B(n921), .Y(n782) );
  NOR2XL U1056 ( .A(n1158), .B(n782), .Y(n811) );
  CMPR32X1 U1057 ( .A(n791), .B(n790), .C(n789), .CO(n792), .S(n828) );
  CMPR32X1 U1058 ( .A(n794), .B(n793), .C(n792), .CO(n803), .S(n832) );
  OAI22X1 U1059 ( .A0(n7), .A1(n838), .B0(n918), .B1(n804), .Y(n843) );
  XNOR2X1 U1060 ( .A(n209), .B(n878), .Y(n839) );
  OAI22X1 U1061 ( .A0(n1161), .A1(n839), .B0(n1162), .B1(n805), .Y(n842) );
  XNOR2X1 U1062 ( .A(n1121), .B(n851), .Y(n840) );
  OAI22XL U1063 ( .A0(n966), .A1(n840), .B0(n9), .B1(n806), .Y(n841) );
  OAI22XL U1064 ( .A0(n972), .A1(n844), .B0(n845), .B1(n810), .Y(n824) );
  ADDHXL U1065 ( .A(n812), .B(n811), .CO(n789), .S(n823) );
  OAI22X1 U1066 ( .A0(n931), .A1(n849), .B0(n813), .B1(n1037), .Y(n847) );
  XNOR2XL U1067 ( .A(B[16]), .B(A[6]), .Y(n814) );
  NOR2XL U1068 ( .A(n328), .B(n814), .Y(n846) );
  CMPR32X1 U1069 ( .A(n824), .B(n822), .C(n823), .CO(n825), .S(n866) );
  CMPR32X1 U1070 ( .A(n827), .B(n826), .C(n825), .CO(n836), .S(n870) );
  OAI22X1 U1071 ( .A0(n7), .A1(n876), .B0(n918), .B1(n838), .Y(n882) );
  XNOR2X1 U1072 ( .A(n209), .B(n921), .Y(n877) );
  OAI22X1 U1073 ( .A0(n1161), .A1(n877), .B0(n1162), .B1(n839), .Y(n881) );
  XNOR2X1 U1074 ( .A(n1121), .B(n892), .Y(n879) );
  OAI22XL U1075 ( .A0(n1139), .A1(n879), .B0(n9), .B1(n840), .Y(n880) );
  XNOR2XL U1076 ( .A(n712), .B(n916), .Y(n884) );
  OAI22XL U1077 ( .A0(n972), .A1(n884), .B0(n845), .B1(n844), .Y(n862) );
  XNOR2X1 U1078 ( .A(n888), .B(n848), .Y(n889) );
  XNOR2XL U1079 ( .A(B[16]), .B(n919), .Y(n850) );
  NOR2XL U1080 ( .A(n1158), .B(n850), .Y(n885) );
  CMPR32X1 U1081 ( .A(n862), .B(n861), .C(n860), .CO(n863), .S(n907) );
  CMPR32X1 U1082 ( .A(n865), .B(n864), .C(n863), .CO(n874), .S(n911) );
  OAI22X1 U1083 ( .A0(n7), .A1(n917), .B0(n918), .B1(n876), .Y(n925) );
  OAI22XL U1084 ( .A0(n966), .A1(n922), .B0(n9), .B1(n879), .Y(n923) );
  XNOR2XL U1085 ( .A(n712), .B(n883), .Y(n927) );
  OAI22XL U1086 ( .A0(n972), .A1(n927), .B0(n970), .B1(n884), .Y(n903) );
  ADDHXL U1087 ( .A(n886), .B(n885), .CO(n860), .S(n902) );
  XNOR2XL U1088 ( .A(B[16]), .B(n890), .Y(n891) );
  OAI22X1 U1089 ( .A0(n939), .A1(n936), .B0(n937), .B1(n895), .Y(n944) );
  OAI22X1 U1090 ( .A0(n942), .A1(n940), .B0(n654), .B1(n897), .Y(n943) );
  CMPR32X1 U1091 ( .A(n903), .B(n901), .C(n902), .CO(n904), .S(n951) );
  CMPR32X1 U1092 ( .A(n906), .B(n905), .C(n904), .CO(n915), .S(n955) );
  XNOR2X1 U1093 ( .A(n209), .B(n919), .Y(n962) );
  XNOR2XL U1094 ( .A(n1121), .B(n921), .Y(n964) );
  OAI22XL U1095 ( .A0(n966), .A1(n964), .B0(n9), .B1(n922), .Y(n967) );
  XNOR2XL U1096 ( .A(n712), .B(n926), .Y(n969) );
  OAI22XL U1097 ( .A0(n972), .A1(n969), .B0(n970), .B1(n927), .Y(n947) );
  XNOR2XL U1098 ( .A(B[16]), .B(n932), .Y(n933) );
  NOR2XL U1099 ( .A(n1158), .B(n933), .Y(n973) );
  OAI22X1 U1100 ( .A0(n8), .A1(n935), .B0(n6), .B1(n934), .Y(n982) );
  CMPR32X1 U1101 ( .A(n947), .B(n946), .C(n945), .CO(n948), .S(n989) );
  CMPR32X1 U1102 ( .A(n950), .B(n949), .C(n948), .CO(n959), .S(n993) );
  OAI22XL U1103 ( .A0(n966), .A1(n965), .B0(n9), .B1(n964), .Y(n1001) );
  OAI22XL U1104 ( .A0(n972), .A1(n971), .B0(n970), .B1(n969), .Y(n985) );
  ADDHXL U1105 ( .A(n974), .B(n973), .CO(n945), .S(n984) );
  CMPR32X1 U1106 ( .A(n979), .B(n978), .C(n977), .CO(n1015), .S(n1022) );
  CMPR32X1 U1107 ( .A(n985), .B(n983), .C(n984), .CO(n986), .S(n1013) );
  CMPR32X1 U1108 ( .A(n988), .B(n987), .C(n986), .CO(n997), .S(n1017) );
  CMPR32X1 U1109 ( .A(n1000), .B(n999), .C(n998), .CO(n1012), .S(n1008) );
  CMPR32X1 U1110 ( .A(n1003), .B(n1002), .C(n1001), .CO(n988), .S(n1011) );
  CMPR32X1 U1111 ( .A(n1006), .B(n1005), .C(n1004), .CO(n1010), .S(n1007) );
  CMPR32X1 U1112 ( .A(n1012), .B(n1011), .C(n1010), .CO(n1021), .S(n1029) );
  CMPR32X1 U1113 ( .A(n1024), .B(n1023), .C(n1022), .CO(n1033), .S(n1036) );
  CMPR32X1 U1114 ( .A(n1033), .B(n1032), .C(n1031), .CO(mult_x_1_n649), .S(
        mult_x_1_n650) );
  INVXL U1115 ( .A(n1043), .Y(n1045) );
  INVXL U1116 ( .A(n1280), .Y(n1050) );
  OAI21XL U1117 ( .A0(n1250), .A1(n1053), .B0(n1052), .Y(n1056) );
  INVXL U1118 ( .A(n1277), .Y(n1054) );
  XNOR2X2 U1119 ( .A(n1056), .B(n1055), .Y(PRODUCT[32]) );
  CMPR32X1 U1120 ( .A(n1059), .B(n1058), .C(n1057), .CO(n1092), .S(n1103) );
  ADDFHX1 U1121 ( .A(n1062), .B(n1061), .CI(n1060), .CO(n1102), .S(n1072) );
  CMPR32X1 U1122 ( .A(n1068), .B(n1067), .C(n1066), .CO(n1087), .S(n1090) );
  NOR2X1 U1123 ( .A(n1077), .B(n1076), .Y(n1075) );
  NAND2XL U1124 ( .A(n1105), .B(n689), .Y(n1081) );
  NAND2XL U1125 ( .A(n1077), .B(n1076), .Y(n1104) );
  INVXL U1126 ( .A(n1104), .Y(n1078) );
  AOI21XL U1127 ( .A0(n1105), .A1(n1079), .B0(n1078), .Y(n1080) );
  OAI21XL U1128 ( .A0(n1082), .A1(n1081), .B0(n1080), .Y(mult_x_1_n309) );
  ADDFHX1 U1129 ( .A(n1088), .B(n1087), .CI(n1086), .CO(n656), .S(n1100) );
  CMPR32X1 U1130 ( .A(n1094), .B(n1093), .C(n1092), .CO(n1084), .S(n1098) );
  INVXL U1131 ( .A(n1097), .Y(mult_x_1_n298) );
  NAND2XL U1132 ( .A(n24), .B(n1097), .Y(mult_x_1_n83) );
  CMPR32X1 U1133 ( .A(n1100), .B(n1099), .C(n1098), .CO(n1095), .S(n1110) );
  ADDFHX1 U1134 ( .A(n1103), .B(n1102), .CI(n1101), .CO(n1109), .S(n1077) );
  OR2X2 U1135 ( .A(n1110), .B(n1109), .Y(n1317) );
  NAND2XL U1136 ( .A(n1105), .B(n1104), .Y(mult_x_1_n85) );
  NAND2XL U1137 ( .A(n689), .B(n1106), .Y(mult_x_1_n86) );
  CMPR32X1 U1138 ( .A(n1114), .B(n1113), .C(n1112), .CO(n1127), .S(n1107) );
  CMPR32X1 U1139 ( .A(n1117), .B(n1116), .C(n1115), .CO(n1130), .S(n1114) );
  XNOR2X1 U1140 ( .A(n209), .B(n1145), .Y(n1131) );
  XNOR2XL U1141 ( .A(n1121), .B(A[25]), .Y(n1137) );
  OAI22X1 U1142 ( .A0(n1139), .A1(n1122), .B0(n9), .B1(n1137), .Y(n1150) );
  CMPR32X1 U1143 ( .A(n1125), .B(n1124), .C(n1123), .CO(n1128), .S(n1113) );
  CMPR32X1 U1144 ( .A(n1130), .B(n1129), .C(n1128), .CO(n1141), .S(n1126) );
  XNOR2XL U1145 ( .A(n209), .B(A[24]), .Y(n1147) );
  CMPR32X1 U1146 ( .A(n1134), .B(n1133), .C(n1132), .CO(n1143), .S(n1129) );
  OAI2BB1X1 U1147 ( .A0N(n9), .A1N(n1139), .B0(n1138), .Y(n1148) );
  CMPR32X1 U1148 ( .A(n1144), .B(n1143), .C(n1142), .CO(n1152), .S(n1140) );
  XNOR2XL U1149 ( .A(n209), .B(A[25]), .Y(n1159) );
  CMPR32X1 U1150 ( .A(n1150), .B(n1149), .C(n1148), .CO(n1153), .S(n1142) );
  CMPR32X1 U1151 ( .A(n1155), .B(n1154), .C(n1153), .CO(n1167), .S(n1151) );
  XNOR2XL U1152 ( .A(n1156), .B(A[24]), .Y(n1157) );
  XOR3X2 U1153 ( .A(n1165), .B(n1164), .C(n1163), .Y(n1166) );
  OAI21XL U1154 ( .A0(n1175), .A1(n1276), .B0(n1174), .Y(n1243) );
  OAI21XL U1155 ( .A0(n1250), .A1(n1180), .B0(n1179), .Y(n1183) );
  OAI21XL U1156 ( .A0(n1250), .A1(n1185), .B0(n1184), .Y(n1188) );
  XNOR2X1 U1157 ( .A(n1192), .B(n1191), .Y(n1333) );
  OAI21XL U1158 ( .A0(n1202), .A1(n1199), .B0(n1200), .Y(n1198) );
  INVXL U1159 ( .A(n1194), .Y(n1196) );
  OAI21XL U1160 ( .A0(n1267), .A1(n1270), .B0(n1268), .Y(n1212) );
  AOI21XL U1161 ( .A0(n1215), .A1(n1208), .B0(n1212), .Y(n1204) );
  OAI21XL U1162 ( .A0(n1250), .A1(n1205), .B0(n1204), .Y(n1207) );
  AOI21XL U1163 ( .A0(n1215), .A1(n1214), .B0(n1213), .Y(n1216) );
  OAI21XL U1164 ( .A0(n1250), .A1(n1217), .B0(n1216), .Y(n1220) );
  XOR2XL U1165 ( .A(n1229), .B(n1228), .Y(n1338) );
  XNOR2XL U1166 ( .A(n1232), .B(n1231), .Y(n1337) );
  XNOR2XL U1167 ( .A(n1236), .B(n1235), .Y(n1339) );
  OAI21XL U1168 ( .A0(n1240), .A1(n1263), .B0(n1264), .Y(n1241) );
  OAI21XL U1169 ( .A0(n1246), .A1(n1245), .B0(n1244), .Y(n1247) );
  OAI21XL U1170 ( .A0(n1250), .A1(n1249), .B0(n1248), .Y(n1251) );
  XNOR2XL U1171 ( .A(n1251), .B(n1262), .Y(PRODUCT[40]) );
  XOR2XL U1172 ( .A(n1256), .B(n1255), .Y(n1336) );
endmodule


module FFT2048_DW02_mult_2_stage_J1_18 ( A, B, TC, CLK, PRODUCT );
  input [15:0] A;
  input [26:0] B;
  output [42:0] PRODUCT;
  input TC, CLK;
  wire   n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, mult_x_1_n679, mult_x_1_n666, mult_x_1_n665, mult_x_1_n652,
         mult_x_1_n651, mult_x_1_n638, mult_x_1_n637, mult_x_1_n625,
         mult_x_1_n624, mult_x_1_n623, mult_x_1_n614, mult_x_1_n612,
         mult_x_1_n611, mult_x_1_n600, mult_x_1_n598, mult_x_1_n597,
         mult_x_1_n586, mult_x_1_n584, mult_x_1_n583, mult_x_1_n572,
         mult_x_1_n570, mult_x_1_n569, mult_x_1_n558, mult_x_1_n556,
         mult_x_1_n555, mult_x_1_n544, mult_x_1_n542, mult_x_1_n541,
         mult_x_1_n530, mult_x_1_n528, mult_x_1_n527, mult_x_1_n516,
         mult_x_1_n514, mult_x_1_n513, mult_x_1_n502, mult_x_1_n500,
         mult_x_1_n499, mult_x_1_n488, mult_x_1_n487, mult_x_1_n486,
         mult_x_1_n485, mult_x_1_n474, mult_x_1_n473, mult_x_1_n464,
         mult_x_1_n463, mult_x_1_n462, mult_x_1_n461, mult_x_1_n453,
         mult_x_1_n452, mult_x_1_n451, mult_x_1_n443, mult_x_1_n442,
         mult_x_1_n441, mult_x_1_n434, mult_x_1_n433, mult_x_1_n428,
         mult_x_1_n427, mult_x_1_n426, mult_x_1_n425, mult_x_1_n421,
         mult_x_1_n420, mult_x_1_n419, mult_x_1_n414, mult_x_1_n408,
         mult_x_1_n407, mult_x_1_n404, mult_x_1_n388, mult_x_1_n387,
         mult_x_1_n361, mult_x_1_n317, mult_x_1_n312, mult_x_1_n310,
         mult_x_1_n305, mult_x_1_n297, mult_x_1_n296, mult_x_1_n100,
         mult_x_1_n81, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198;

  DFFHQX1 mult_x_1_clk_r_REG9_S1 ( .D(mult_x_1_n611), .CK(CLK), .Q(n1186) );
  DFFHQXL mult_x_1_clk_r_REG1_S1 ( .D(mult_x_1_n666), .CK(CLK), .Q(n1197) );
  DFFHQXL mult_x_1_clk_r_REG66_S1 ( .D(mult_x_1_n679), .CK(CLK), .Q(n1198) );
  DFFHQXL mult_x_1_clk_r_REG3_S1 ( .D(mult_x_1_n652), .CK(CLK), .Q(n1195) );
  DFFHQXL mult_x_1_clk_r_REG5_S1 ( .D(mult_x_1_n638), .CK(CLK), .Q(n1193) );
  DFFHQXL mult_x_1_clk_r_REG4_S1 ( .D(mult_x_1_n637), .CK(CLK), .Q(n1192) );
  DFFHQXL mult_x_1_clk_r_REG7_S1 ( .D(mult_x_1_n624), .CK(CLK), .Q(n1190) );
  DFFHQXL mult_x_1_clk_r_REG6_S1 ( .D(mult_x_1_n623), .CK(CLK), .Q(n1189) );
  DFFHQX4 mult_x_1_clk_r_REG11_S1 ( .D(mult_x_1_n614), .CK(CLK), .Q(n1188) );
  DFFHQXL mult_x_1_clk_r_REG67_S1 ( .D(mult_x_1_n297), .CK(CLK), .Q(n1127) );
  DFFHQXL mult_x_1_clk_r_REG22_S1 ( .D(mult_x_1_n500), .CK(CLK), .Q(n1163) );
  DFFHQXL mult_x_1_clk_r_REG19_S1 ( .D(mult_x_1_n514), .CK(CLK), .Q(n1166) );
  DFFHQXL mult_x_1_clk_r_REG25_S1 ( .D(mult_x_1_n486), .CK(CLK), .Q(n1159) );
  DFFHQXL mult_x_1_clk_r_REG37_S1 ( .D(mult_x_1_n584), .CK(CLK), .Q(n1181) );
  DFFHQX1 mult_x_1_clk_r_REG70_S1 ( .D(mult_x_1_n387), .CK(CLK), .Q(n1122) );
  DFFHQXL mult_x_1_clk_r_REG53_S1 ( .D(mult_x_1_n451), .CK(CLK), .Q(n1149) );
  DFFHQXL mult_x_1_clk_r_REG16_S1 ( .D(mult_x_1_n528), .CK(CLK), .Q(n1169) );
  DFFHQXL mult_x_1_clk_r_REG28_S1 ( .D(mult_x_1_n542), .CK(CLK), .Q(n1172) );
  DFFHQX4 mult_x_1_clk_r_REG15_S1 ( .D(mult_x_1_n527), .CK(CLK), .Q(n1168) );
  DFFHQXL mult_x_1_clk_r_REG24_S1 ( .D(mult_x_1_n485), .CK(CLK), .Q(n1158) );
  DFFHQXL mult_x_1_clk_r_REG41_S1 ( .D(mult_x_1_n474), .CK(CLK), .Q(n1157) );
  DFFHQXL mult_x_1_clk_r_REG43_S1 ( .D(mult_x_1_n462), .CK(CLK), .Q(n1153) );
  DFFHQXL mult_x_1_clk_r_REG74_S1 ( .D(mult_x_1_n312), .CK(CLK), .Q(n1131) );
  DFFHQXL mult_x_1_clk_r_REG63_S1 ( .D(mult_x_1_n407), .CK(CLK), .Q(n1134) );
  DFFHQXL mult_x_1_clk_r_REG46_S1 ( .D(mult_x_1_n433), .CK(CLK), .Q(n1144) );
  DFFHQXL mult_x_1_clk_r_REG64_S1 ( .D(mult_x_1_n408), .CK(CLK), .Q(n1135) );
  DFFHQXL mult_x_1_clk_r_REG77_S1 ( .D(mult_x_1_n317), .CK(CLK), .Q(n1132) );
  DFFHQXL mult_x_1_clk_r_REG56_S1 ( .D(mult_x_1_n441), .CK(CLK), .Q(n1146) );
  DFFHQXL mult_x_1_clk_r_REG49_S1 ( .D(mult_x_1_n426), .CK(CLK), .Q(n1141) );
  DFFHQXL clk_r_REG78_S1 ( .D(n1211), .CK(CLK), .Q(PRODUCT[9]) );
  DFFHQXL mult_x_1_clk_r_REG13_S1 ( .D(mult_x_1_n598), .CK(CLK), .Q(n1184) );
  DFFHQXL mult_x_1_clk_r_REG54_S1 ( .D(mult_x_1_n452), .CK(CLK), .Q(n1150) );
  DFFHQXL mult_x_1_clk_r_REG68_S1 ( .D(mult_x_1_n296), .CK(CLK), .Q(n1126) );
  DFFHQXL mult_x_1_clk_r_REG0_S1 ( .D(mult_x_1_n665), .CK(CLK), .Q(n1196) );
  DFFHQXL clk_r_REG80_S1 ( .D(n1213), .CK(CLK), .Q(PRODUCT[7]) );
  DFFHQXL mult_x_1_clk_r_REG2_S1 ( .D(mult_x_1_n651), .CK(CLK), .Q(n1194) );
  DFFHQXL mult_x_1_clk_r_REG75_S1 ( .D(mult_x_1_n421), .CK(CLK), .Q(n1139) );
  DFFHQXL mult_x_1_clk_r_REG38_S1 ( .D(mult_x_1_n487), .CK(CLK), .Q(n1160) );
  DFFHQXL mult_x_1_clk_r_REG30_S1 ( .D(mult_x_1_n570), .CK(CLK), .Q(n1178) );
  DFFHQXL clk_r_REG76_S1 ( .D(n1210), .CK(CLK), .Q(PRODUCT[10]) );
  DFFHQXL clk_r_REG79_S1 ( .D(n1212), .CK(CLK), .Q(PRODUCT[8]) );
  DFFHQXL clk_r_REG81_S1 ( .D(n1214), .CK(CLK), .Q(PRODUCT[6]) );
  DFFHQXL clk_r_REG82_S1 ( .D(n1215), .CK(CLK), .Q(PRODUCT[5]) );
  DFFHQXL clk_r_REG83_S1 ( .D(n1216), .CK(CLK), .Q(PRODUCT[4]) );
  DFFHQXL clk_r_REG84_S1 ( .D(n1217), .CK(CLK), .Q(PRODUCT[3]) );
  DFFHQXL clk_r_REG85_S1 ( .D(n1218), .CK(CLK), .Q(PRODUCT[2]) );
  DFFHQXL clk_r_REG86_S1 ( .D(n1219), .CK(CLK), .Q(PRODUCT[1]) );
  DFFHQXL clk_r_REG87_S1 ( .D(n1220), .CK(CLK), .Q(PRODUCT[0]) );
  DFFHQX1 mult_x_1_clk_r_REG35_S1 ( .D(mult_x_1_n600), .CK(CLK), .Q(n1185) );
  DFFHQX1 mult_x_1_clk_r_REG33_S1 ( .D(mult_x_1_n586), .CK(CLK), .Q(n1182) );
  DFFHQX1 mult_x_1_clk_r_REG36_S1 ( .D(mult_x_1_n583), .CK(CLK), .Q(n1180) );
  DFFHQX1 mult_x_1_clk_r_REG34_S1 ( .D(mult_x_1_n572), .CK(CLK), .Q(n1179) );
  DFFHQX1 mult_x_1_clk_r_REG29_S1 ( .D(mult_x_1_n569), .CK(CLK), .Q(n1177) );
  DFFHQX1 mult_x_1_clk_r_REG26_S1 ( .D(mult_x_1_n558), .CK(CLK), .Q(n1176) );
  DFFHQX1 mult_x_1_clk_r_REG14_S1 ( .D(mult_x_1_n544), .CK(CLK), .Q(n1173) );
  DFFHQX1 mult_x_1_clk_r_REG17_S1 ( .D(mult_x_1_n530), .CK(CLK), .Q(n1170) );
  DFFHQX1 mult_x_1_clk_r_REG20_S1 ( .D(mult_x_1_n516), .CK(CLK), .Q(n1167) );
  DFFHQXL mult_x_1_clk_r_REG39_S1 ( .D(mult_x_1_n488), .CK(CLK), .Q(n1161) );
  DFFHQXL mult_x_1_clk_r_REG42_S1 ( .D(mult_x_1_n461), .CK(CLK), .Q(n1152) );
  DFFHQXL mult_x_1_clk_r_REG55_S1 ( .D(mult_x_1_n443), .CK(CLK), .Q(n1148) );
  DFFHQXL mult_x_1_clk_r_REG57_S1 ( .D(mult_x_1_n442), .CK(CLK), .Q(n1147) );
  DFFHQXL mult_x_1_clk_r_REG47_S1 ( .D(mult_x_1_n434), .CK(CLK), .Q(n1145) );
  DFFHQXL mult_x_1_clk_r_REG51_S1 ( .D(mult_x_1_n428), .CK(CLK), .Q(n1143) );
  DFFHQXL mult_x_1_clk_r_REG50_S1 ( .D(mult_x_1_n427), .CK(CLK), .Q(n1142) );
  DFFHQXL mult_x_1_clk_r_REG48_S1 ( .D(mult_x_1_n425), .CK(CLK), .Q(n1140) );
  DFFHQXL mult_x_1_clk_r_REG59_S1 ( .D(mult_x_1_n420), .CK(CLK), .Q(n1138) );
  DFFHQXL mult_x_1_clk_r_REG58_S1 ( .D(mult_x_1_n419), .CK(CLK), .Q(n1137) );
  DFFHQXL mult_x_1_clk_r_REG62_S1 ( .D(mult_x_1_n414), .CK(CLK), .Q(n1136) );
  DFFHQXL mult_x_1_clk_r_REG65_S1 ( .D(mult_x_1_n404), .CK(CLK), .Q(n1133) );
  DFFHQXL mult_x_1_clk_r_REG73_S1 ( .D(mult_x_1_n81), .CK(CLK), .Q(n1130) );
  DFFHQX2 mult_x_1_clk_r_REG71_S1 ( .D(mult_x_1_n310), .CK(CLK), .Q(n1129) );
  DFFHQXL mult_x_1_clk_r_REG60_S1 ( .D(mult_x_1_n100), .CK(CLK), .Q(n1125) );
  DFFHQXL mult_x_1_clk_r_REG61_S1 ( .D(mult_x_1_n361), .CK(CLK), .Q(n1124) );
  DFFHQX1 mult_x_1_clk_r_REG69_S1 ( .D(mult_x_1_n305), .CK(CLK), .Q(n1128) );
  DFFHQXL mult_x_1_clk_r_REG44_S1 ( .D(mult_x_1_n463), .CK(CLK), .Q(n1154) );
  DFFHQXL mult_x_1_clk_r_REG45_S1 ( .D(mult_x_1_n464), .CK(CLK), .Q(n1155) );
  DFFHQXL mult_x_1_clk_r_REG52_S1 ( .D(mult_x_1_n453), .CK(CLK), .Q(n1151) );
  DFFHQX1 mult_x_1_clk_r_REG10_S1 ( .D(mult_x_1_n612), .CK(CLK), .Q(n1187) );
  DFFHQXL mult_x_1_clk_r_REG32_S1 ( .D(mult_x_1_n556), .CK(CLK), .Q(n1175) );
  DFFHQXL mult_x_1_clk_r_REG21_S1 ( .D(mult_x_1_n499), .CK(CLK), .Q(n1162) );
  DFFHQX4 mult_x_1_clk_r_REG31_S1 ( .D(mult_x_1_n555), .CK(CLK), .Q(n1174) );
  DFFHQXL mult_x_1_clk_r_REG40_S1 ( .D(mult_x_1_n473), .CK(CLK), .Q(n1156) );
  DFFHQX1 mult_x_1_clk_r_REG27_S1 ( .D(mult_x_1_n541), .CK(CLK), .Q(n1171) );
  DFFHQX1 mult_x_1_clk_r_REG23_S1 ( .D(mult_x_1_n502), .CK(CLK), .Q(n1164) );
  DFFHQX2 mult_x_1_clk_r_REG8_S1 ( .D(mult_x_1_n625), .CK(CLK), .Q(n1191) );
  DFFHQX1 mult_x_1_clk_r_REG72_S1 ( .D(mult_x_1_n388), .CK(CLK), .Q(n1123) );
  DFFHQX1 mult_x_1_clk_r_REG12_S1 ( .D(mult_x_1_n597), .CK(CLK), .Q(n1183) );
  DFFHQX2 mult_x_1_clk_r_REG18_S1 ( .D(mult_x_1_n513), .CK(CLK), .Q(n1165) );
  ADDFHX1 U1 ( .A(n950), .B(n949), .CI(n948), .CO(mult_x_1_n637), .S(
        mult_x_1_n638) );
  ADDFHX1 U2 ( .A(n684), .B(n683), .CI(n682), .CO(mult_x_1_n513), .S(
        mult_x_1_n514) );
  ADDFHX1 U3 ( .A(n552), .B(n551), .CI(n550), .CO(mult_x_1_n451), .S(
        mult_x_1_n452) );
  ADDFHX1 U4 ( .A(n971), .B(n970), .CI(n969), .CO(mult_x_1_n651), .S(
        mult_x_1_n652) );
  ADDFHX2 U5 ( .A(n947), .B(n946), .CI(n945), .CO(n919), .S(n948) );
  NAND2XL U6 ( .A(n29), .B(n575), .Y(n30) );
  ADDFHX1 U7 ( .A(n968), .B(n967), .CI(n966), .CO(n949), .S(n969) );
  ADDFHX1 U8 ( .A(n687), .B(n686), .CI(n685), .CO(n656), .S(mult_x_1_n516) );
  ADDFHX1 U9 ( .A(n875), .B(n874), .CI(n873), .CO(n867), .S(n920) );
  ADDFHX1 U10 ( .A(n715), .B(n714), .CI(n713), .CO(n682), .S(mult_x_1_n530) );
  ADDFHX2 U11 ( .A(n681), .B(n680), .CI(n679), .CO(n686), .S(n713) );
  CMPR32X1 U12 ( .A(n962), .B(n961), .C(n960), .CO(n968), .S(n978) );
  ADDFHX1 U13 ( .A(n926), .B(n925), .CI(n924), .CO(n921), .S(n950) );
  ADDFHX1 U14 ( .A(n944), .B(n943), .CI(n942), .CO(n947), .S(n966) );
  ADDFHX1 U15 ( .A(n697), .B(n696), .CI(n695), .CO(n714), .S(n707) );
  ADDFHX1 U16 ( .A(n974), .B(n48), .CI(n972), .CO(n967), .S(n982) );
  INVX1 U17 ( .A(n29), .Y(n28) );
  ADDFHX2 U18 ( .A(n914), .B(n913), .CI(n912), .CO(n925), .S(n951) );
  ADDFHX1 U19 ( .A(n917), .B(n916), .CI(n915), .CO(n874), .S(n924) );
  OAI22X2 U20 ( .A0(n590), .A1(n257), .B0(n614), .B1(n258), .Y(n611) );
  ADDFHX1 U21 ( .A(n900), .B(n901), .CI(n899), .CO(n917), .S(n913) );
  ADDFHX1 U22 ( .A(n42), .B(n861), .CI(n860), .CO(n866), .S(n916) );
  ADDFHX1 U23 ( .A(n363), .B(n362), .CI(n361), .CO(n456), .S(n455) );
  ADDFHX1 U24 ( .A(n929), .B(n928), .CI(n927), .CO(n962), .S(n955) );
  ADDFHX1 U25 ( .A(n878), .B(n877), .CI(n876), .CO(n941), .S(n928) );
  CMPR22X1 U26 ( .A(n290), .B(n289), .CO(n877), .S(n286) );
  ADDFX2 U27 ( .A(n417), .B(n416), .CI(n415), .CO(n422), .S(n421) );
  ADDFHX1 U28 ( .A(n367), .B(n366), .CI(n365), .CO(n373), .S(n383) );
  CLKBUFX3 U29 ( .A(n288), .Y(n529) );
  BUFX3 U30 ( .A(n572), .Y(n102) );
  INVX1 U31 ( .A(A[13]), .Y(n264) );
  CLKBUFX3 U32 ( .A(n497), .Y(n499) );
  INVX4 U33 ( .A(n498), .Y(n8) );
  INVX4 U34 ( .A(n275), .Y(n7) );
  XNOR2X2 U35 ( .A(A[4]), .B(A[3]), .Y(n528) );
  OAI21XL U36 ( .A0(n1038), .A1(n1037), .B0(n1036), .Y(n1104) );
  XNOR2X2 U37 ( .A(n167), .B(n166), .Y(PRODUCT[31]) );
  INVX1 U38 ( .A(n34), .Y(n1029) );
  XNOR2X1 U39 ( .A(n230), .B(n229), .Y(PRODUCT[21]) );
  XNOR2X1 U40 ( .A(n93), .B(n92), .Y(PRODUCT[20]) );
  AOI21X2 U41 ( .A0(n213), .A1(n123), .B0(n20), .Y(n69) );
  NOR2X2 U42 ( .A(n208), .B(n215), .Y(n123) );
  OAI21X2 U43 ( .A0(n222), .A1(n227), .B0(n223), .Y(n213) );
  NOR2X2 U44 ( .A(n118), .B(n117), .Y(n222) );
  CMPR32X1 U45 ( .A(n1151), .B(n1147), .C(n1149), .CO(n146), .S(n140) );
  NAND2X1 U46 ( .A(n116), .B(n115), .Y(n227) );
  NOR2X1 U47 ( .A(n116), .B(n115), .Y(n220) );
  NAND2X1 U48 ( .A(n35), .B(n236), .Y(n108) );
  ADDFHX1 U49 ( .A(n1185), .B(n1186), .CI(n1184), .CO(n115), .S(n90) );
  ADDFHX1 U50 ( .A(n1176), .B(n1177), .CI(n1175), .CO(n121), .S(n120) );
  ADDFHX1 U51 ( .A(n1173), .B(n1174), .CI(n1172), .CO(n124), .S(n122) );
  XNOR2X2 U52 ( .A(B[7]), .B(n856), .Y(n765) );
  OAI22X1 U53 ( .A0(n742), .A1(n529), .B0(n790), .B1(n102), .Y(n793) );
  CMPR22X1 U54 ( .A(n793), .B(n792), .CO(n767), .S(n827) );
  INVXL U55 ( .A(n357), .Y(n5) );
  INVXL U56 ( .A(n5), .Y(n6) );
  AOI21XL U57 ( .A0(n159), .A1(n143), .B0(n142), .Y(n23) );
  NOR2X2 U58 ( .A(n220), .B(n222), .Y(n214) );
  XNOR2XL U59 ( .A(B[4]), .B(n858), .Y(n886) );
  XNOR2XL U60 ( .A(B[6]), .B(n9), .Y(n327) );
  XNOR2XL U61 ( .A(B[15]), .B(A[11]), .Y(n49) );
  XNOR2XL U62 ( .A(B[6]), .B(n858), .Y(n859) );
  XNOR2XL U63 ( .A(B[6]), .B(n895), .Y(n282) );
  INVX4 U64 ( .A(n264), .Y(n856) );
  XNOR2XL U65 ( .A(B[13]), .B(n856), .Y(n639) );
  XNOR2XL U66 ( .A(B[14]), .B(A[7]), .Y(n773) );
  XNOR2XL U67 ( .A(B[26]), .B(A[7]), .Y(n500) );
  XNOR2XL U68 ( .A(B[19]), .B(A[5]), .Y(n717) );
  XNOR2XL U69 ( .A(B[9]), .B(n858), .Y(n794) );
  XNOR2XL U70 ( .A(B[9]), .B(n895), .Y(n931) );
  XNOR2XL U71 ( .A(B[25]), .B(A[11]), .Y(n489) );
  BUFX3 U72 ( .A(n665), .Y(n258) );
  XOR2X2 U73 ( .A(n576), .B(n575), .Y(n13) );
  NOR2XL U74 ( .A(n1028), .B(n1027), .Y(n996) );
  NAND2X1 U75 ( .A(n457), .B(n456), .Y(n1025) );
  ADDFHX1 U76 ( .A(n630), .B(n629), .CI(n628), .CO(n635), .S(n659) );
  INVX1 U77 ( .A(n547), .Y(n583) );
  ADDFHX1 U78 ( .A(n778), .B(n777), .CI(n776), .CO(n770), .S(n811) );
  OAI2BB1X1 U79 ( .A0N(n832), .A1N(n665), .B0(n96), .Y(n472) );
  OAI2BB1X1 U80 ( .A0N(n497), .A1N(n8), .B0(n496), .Y(n508) );
  NAND2XL U81 ( .A(n839), .B(n840), .Y(n72) );
  OR2X2 U82 ( .A(n423), .B(n422), .Y(n403) );
  NAND2BX1 U83 ( .AN(n1006), .B(n34), .Y(n26) );
  XOR2X2 U84 ( .A(n226), .B(n225), .Y(PRODUCT[22]) );
  NAND3X2 U85 ( .A(n25), .B(n24), .C(n23), .Y(n34) );
  XNOR2X1 U86 ( .A(n248), .B(n247), .Y(PRODUCT[16]) );
  INVXL U87 ( .A(n1104), .Y(n1039) );
  INVX1 U88 ( .A(n239), .Y(n248) );
  NAND2X1 U89 ( .A(n91), .B(n109), .Y(n92) );
  NAND2X1 U90 ( .A(n1017), .B(n1016), .Y(n1018) );
  XNOR2X1 U91 ( .A(n9), .B(A[6]), .Y(n497) );
  NAND2X4 U92 ( .A(n617), .B(n256), .Y(n329) );
  NAND2X1 U93 ( .A(n1030), .B(n1035), .Y(n1038) );
  INVX1 U94 ( .A(n1011), .Y(n1013) );
  AND2X2 U95 ( .A(n1035), .B(n1032), .Y(n1009) );
  AND2X2 U96 ( .A(n1103), .B(n1056), .Y(n1042) );
  NAND2X1 U97 ( .A(n135), .B(n134), .Y(n180) );
  NAND2X1 U98 ( .A(n139), .B(n138), .Y(n164) );
  NAND2X1 U99 ( .A(n125), .B(n124), .Y(n1012) );
  NOR2X1 U100 ( .A(n125), .B(n124), .Y(n1011) );
  CLKINVX3 U101 ( .A(n518), .Y(n895) );
  XOR2X1 U102 ( .A(A[3]), .B(A[2]), .Y(n256) );
  NAND2X1 U103 ( .A(n28), .B(n27), .Y(n31) );
  INVX1 U104 ( .A(n575), .Y(n27) );
  ADDFHX1 U105 ( .A(n661), .B(n659), .CI(n660), .CO(n622), .S(mult_x_1_n502)
         );
  BUFX3 U106 ( .A(n576), .Y(n29) );
  ADDFHX1 U107 ( .A(n812), .B(n811), .CI(n810), .CO(n782), .S(mult_x_1_n586)
         );
  NAND2BXL U108 ( .AN(n578), .B(n17), .Y(n15) );
  INVXL U109 ( .A(n578), .Y(n16) );
  OAI22XL U110 ( .A0(n766), .A1(n884), .B0(n765), .B1(n882), .Y(n800) );
  ADDFHX1 U111 ( .A(n384), .B(n383), .CI(n382), .CO(n376), .S(n386) );
  XOR2X1 U112 ( .A(n1075), .B(n1074), .Y(PRODUCT[38]) );
  NAND2X1 U113 ( .A(n26), .B(n1005), .Y(n1010) );
  OAI21XL U114 ( .A0(n1029), .A1(n1106), .B0(n1105), .Y(n1110) );
  OAI2BB1X1 U115 ( .A0N(n1101), .A1N(n34), .B0(n1039), .Y(n1043) );
  NAND3BX1 U116 ( .AN(n144), .B(n11), .C(n1014), .Y(n25) );
  AOI21X1 U117 ( .A0(n230), .A1(n214), .B0(n213), .Y(n219) );
  OAI22XL U118 ( .A0(n304), .A1(n486), .B0(n485), .B1(n501), .Y(n339) );
  NAND2BX1 U119 ( .AN(n144), .B(n170), .Y(n24) );
  NAND2BXL U120 ( .AN(n986), .B(n856), .Y(n263) );
  NAND2X1 U121 ( .A(n228), .B(n227), .Y(n229) );
  NAND2X1 U122 ( .A(n198), .B(n197), .Y(n199) );
  NAND2X1 U123 ( .A(n217), .B(n216), .Y(n218) );
  NAND2X1 U124 ( .A(n12), .B(n1037), .Y(n147) );
  NAND2X1 U125 ( .A(n175), .B(n174), .Y(n176) );
  NAND2X1 U126 ( .A(n181), .B(n180), .Y(n182) );
  INVX1 U127 ( .A(n227), .Y(n221) );
  INVX1 U128 ( .A(n168), .Y(n181) );
  BUFX3 U129 ( .A(n617), .Y(n328) );
  NAND2X1 U130 ( .A(n129), .B(n128), .Y(n197) );
  NAND2X4 U131 ( .A(n267), .B(n268), .Y(n485) );
  BUFX3 U132 ( .A(n267), .Y(n486) );
  NOR2X1 U133 ( .A(n129), .B(n128), .Y(n184) );
  NOR2X1 U134 ( .A(n135), .B(n134), .Y(n168) );
  BUFX3 U135 ( .A(n832), .Y(n257) );
  NAND2X1 U136 ( .A(n832), .B(n95), .Y(n665) );
  XNOR2X1 U137 ( .A(A[1]), .B(A[2]), .Y(n617) );
  NAND2X1 U138 ( .A(n146), .B(n145), .Y(n1037) );
  NAND2X1 U139 ( .A(n288), .B(n94), .Y(n572) );
  NOR2X1 U140 ( .A(n145), .B(n146), .Y(n1031) );
  INVXL U141 ( .A(A[3]), .Y(n19) );
  CLKINVX3 U142 ( .A(A[0]), .Y(n934) );
  INVX4 U143 ( .A(n74), .Y(n9) );
  INVX1 U144 ( .A(A[1]), .Y(n10) );
  OAI2BB1X1 U145 ( .A0N(n31), .A1N(n574), .B0(n30), .Y(mult_x_1_n461) );
  NAND2XL U146 ( .A(n316), .B(n315), .Y(mult_x_1_n297) );
  ADDFHX2 U147 ( .A(n920), .B(n919), .CI(n918), .CO(mult_x_1_n623), .S(
        mult_x_1_n624) );
  ADDFHX2 U148 ( .A(n658), .B(n657), .CI(n656), .CO(mult_x_1_n499), .S(
        mult_x_1_n500) );
  ADDFHX1 U149 ( .A(n784), .B(n783), .CI(n782), .CO(mult_x_1_n569), .S(
        mult_x_1_n570) );
  OAI21XL U150 ( .A0(n16), .A1(n17), .B0(n14), .Y(n586) );
  ADDFHX1 U151 ( .A(n709), .B(n708), .CI(n707), .CO(n710), .S(mult_x_1_n544)
         );
  ADDFHX1 U152 ( .A(n809), .B(n808), .CI(n807), .CO(mult_x_1_n583), .S(
        mult_x_1_n584) );
  ADDFHX1 U153 ( .A(n923), .B(n922), .CI(n921), .CO(mult_x_1_n625), .S(n918)
         );
  ADDFHX1 U154 ( .A(n633), .B(n46), .CI(n631), .CO(n595), .S(n634) );
  ADDFHX1 U155 ( .A(n647), .B(n646), .CI(n645), .CO(n642), .S(n687) );
  ADDFHX1 U156 ( .A(n762), .B(n761), .CI(n760), .CO(n734), .S(mult_x_1_n558)
         );
  NAND2XL U157 ( .A(n15), .B(n577), .Y(n14) );
  NOR2X1 U158 ( .A(n457), .B(n456), .Y(n1024) );
  ADDFHX1 U159 ( .A(n906), .B(n44), .CI(n904), .CO(n923), .S(n946) );
  INVXL U160 ( .A(n37), .Y(n38) );
  ADDFHX1 U161 ( .A(n787), .B(n786), .CI(n785), .CO(n757), .S(mult_x_1_n572)
         );
  NAND2X1 U162 ( .A(n455), .B(n454), .Y(n1020) );
  ADDFHX1 U163 ( .A(n800), .B(n799), .CI(n798), .CO(n795), .S(n846) );
  ADDFHX1 U164 ( .A(n546), .B(n547), .CI(n545), .CO(n535), .S(n554) );
  ADDFHX1 U165 ( .A(n673), .B(n672), .CI(n671), .CO(n668), .S(n715) );
  INVXL U166 ( .A(n632), .Y(n45) );
  INVXL U167 ( .A(n58), .Y(n54) );
  XNOR3X2 U168 ( .A(n957), .B(n955), .C(n956), .Y(n58) );
  INVX1 U169 ( .A(n61), .Y(n605) );
  XNOR2X1 U170 ( .A(B[8]), .B(n895), .Y(n930) );
  OR2X2 U171 ( .A(n413), .B(n412), .Y(n411) );
  XOR2X1 U172 ( .A(n1110), .B(n1109), .Y(PRODUCT[37]) );
  AND2XL U173 ( .A(n1097), .B(n1096), .Y(n1219) );
  ADDFHX1 U174 ( .A(n280), .B(n279), .CI(n278), .CO(n272), .S(n294) );
  OR2XL U175 ( .A(n1095), .B(n1094), .Y(n1097) );
  NAND2X1 U176 ( .A(n33), .B(n1037), .Y(n32) );
  XOR2X1 U177 ( .A(n1043), .B(n1042), .Y(PRODUCT[36]) );
  XNOR2X1 U178 ( .A(n254), .B(n253), .Y(PRODUCT[15]) );
  NAND2XL U179 ( .A(n329), .B(n617), .Y(n18) );
  NOR2BXL U180 ( .AN(n986), .B(n528), .Y(n417) );
  NAND2BXL U181 ( .AN(n986), .B(A[1]), .Y(n405) );
  NOR2BXL U182 ( .AN(n986), .B(n497), .Y(n429) );
  XOR2X1 U183 ( .A(n1118), .B(n1117), .Y(PRODUCT[14]) );
  BUFX3 U184 ( .A(B[0]), .Y(n986) );
  BUFX3 U185 ( .A(n882), .Y(n99) );
  AND2X2 U186 ( .A(n528), .B(n255), .Y(n275) );
  AND2X2 U187 ( .A(n497), .B(n262), .Y(n498) );
  BUFX3 U188 ( .A(n573), .Y(n369) );
  NAND2X1 U189 ( .A(n1013), .B(n1012), .Y(n201) );
  NOR2X1 U190 ( .A(n1038), .B(n1031), .Y(n1101) );
  INVX1 U191 ( .A(n179), .Y(n11) );
  NAND2X1 U192 ( .A(A[1]), .B(n934), .Y(n573) );
  INVX1 U193 ( .A(n232), .Y(n21) );
  AND2XL U194 ( .A(n1073), .B(n1072), .Y(n1074) );
  AND2XL U195 ( .A(n1108), .B(n1107), .Y(n1109) );
  INVXL U196 ( .A(n1012), .Y(n68) );
  INVX1 U197 ( .A(n220), .Y(n228) );
  NAND2X1 U198 ( .A(n122), .B(n121), .Y(n209) );
  NOR2X1 U199 ( .A(n141), .B(n140), .Y(n154) );
  INVX1 U200 ( .A(n1031), .Y(n12) );
  INVX1 U201 ( .A(n231), .Y(n236) );
  INVX1 U202 ( .A(n1189), .Y(n22) );
  ADDFHX2 U203 ( .A(n1188), .B(n1191), .CI(n1187), .CO(n89), .S(n87) );
  ADDFHX1 U204 ( .A(n1154), .B(n1152), .CI(n1150), .CO(n141), .S(n139) );
  AND2XL U205 ( .A(n1124), .B(n1125), .Y(n1063) );
  INVX1 U206 ( .A(A[11]), .Y(n488) );
  INVX1 U207 ( .A(A[7]), .Y(n518) );
  XNOR2X1 U208 ( .A(B[21]), .B(A[7]), .Y(n619) );
  XNOR2X1 U209 ( .A(B[1]), .B(A[9]), .Y(n306) );
  ADDHXL U210 ( .A(n339), .B(n338), .CO(n325), .S(n357) );
  OAI22X1 U211 ( .A0(n519), .A1(n499), .B0(n539), .B1(n8), .Y(n541) );
  XOR2X1 U212 ( .A(B[13]), .B(n518), .Y(n801) );
  OAI22X1 U213 ( .A0(n619), .A1(n8), .B0(n587), .B1(n499), .Y(n609) );
  XNOR2X1 U214 ( .A(B[11]), .B(n9), .Y(n932) );
  XNOR2X1 U215 ( .A(B[22]), .B(A[9]), .Y(n544) );
  XOR2X1 U216 ( .A(n574), .B(n13), .Y(mult_x_1_n462) );
  XNOR3X2 U217 ( .A(n577), .B(n17), .C(n578), .Y(n592) );
  AND2X2 U218 ( .A(n561), .B(n18), .Y(n17) );
  XOR2X1 U219 ( .A(n1023), .B(n1022), .Y(n1210) );
  XOR2X1 U220 ( .A(n599), .B(n600), .Y(n77) );
  XOR2X1 U221 ( .A(B[22]), .B(n19), .Y(n698) );
  XOR2X1 U222 ( .A(B[22]), .B(n10), .Y(n730) );
  OAI22X4 U223 ( .A0(n528), .A1(n567), .B0(n570), .B1(n7), .Y(n580) );
  XNOR2X4 U224 ( .A(B[24]), .B(n9), .Y(n570) );
  XOR2X4 U225 ( .A(B[25]), .B(n74), .Y(n567) );
  XOR2X2 U226 ( .A(n202), .B(n201), .Y(PRODUCT[25]) );
  OAI21X2 U227 ( .A0(n208), .A1(n216), .B0(n209), .Y(n20) );
  NAND2X1 U228 ( .A(n120), .B(n119), .Y(n216) );
  NOR2X2 U229 ( .A(n122), .B(n121), .Y(n208) );
  XNOR2X1 U230 ( .A(B[26]), .B(n10), .Y(n61) );
  XNOR2X1 U231 ( .A(B[1]), .B(n856), .Y(n291) );
  XNOR2X4 U232 ( .A(B[16]), .B(A[11]), .Y(n614) );
  XNOR2X4 U233 ( .A(B[17]), .B(A[11]), .Y(n590) );
  XOR2X1 U234 ( .A(n58), .B(n57), .Y(n56) );
  XNOR2X1 U235 ( .A(B[11]), .B(A[9]), .Y(n802) );
  OAI21X4 U236 ( .A0(n111), .A1(n110), .B0(n109), .Y(n112) );
  NOR2X2 U237 ( .A(n90), .B(n89), .Y(n110) );
  AOI21X2 U238 ( .A0(n35), .A1(n88), .B0(n21), .Y(n111) );
  NAND2X1 U239 ( .A(n87), .B(n1189), .Y(n232) );
  NAND2BX4 U240 ( .AN(n87), .B(n22), .Y(n35) );
  NOR2X1 U241 ( .A(n139), .B(n138), .Y(n163) );
  XOR2X2 U242 ( .A(n32), .B(n1002), .Y(PRODUCT[34]) );
  NAND2X1 U243 ( .A(n34), .B(n12), .Y(n33) );
  OAI21X4 U244 ( .A0(n70), .A1(n204), .B0(n69), .Y(n1014) );
  NOR2X2 U245 ( .A(n120), .B(n119), .Y(n215) );
  XNOR2X1 U246 ( .A(B[3]), .B(n858), .Y(n287) );
  OAI22X2 U247 ( .A0(n291), .A1(n884), .B0(n265), .B1(n882), .Y(n289) );
  XNOR2X1 U248 ( .A(n986), .B(n856), .Y(n265) );
  OAI21X1 U249 ( .A0(n1015), .A1(n1012), .B0(n1016), .Y(n194) );
  XOR2X1 U250 ( .A(n1010), .B(n1009), .Y(PRODUCT[35]) );
  INVX1 U251 ( .A(n856), .Y(n73) );
  OAI22X1 U252 ( .A0(n306), .A1(n486), .B0(n305), .B1(n485), .Y(n338) );
  INVXL U253 ( .A(A[9]), .Y(n501) );
  CMPR22X1 U254 ( .A(n274), .B(n273), .CO(n279), .S(n311) );
  OAI22X1 U255 ( .A0(n259), .A1(n257), .B0(n258), .B1(n488), .Y(n274) );
  OAI22X1 U256 ( .A0(n261), .A1(n257), .B0(n260), .B1(n258), .Y(n273) );
  NAND2BXL U257 ( .AN(n986), .B(A[11]), .Y(n259) );
  NAND2BXL U258 ( .AN(n986), .B(A[7]), .Y(n350) );
  NAND2X1 U259 ( .A(n35), .B(n232), .Y(n233) );
  OAI21XL U260 ( .A0(n202), .A1(n196), .B0(n195), .Y(n200) );
  INVXL U261 ( .A(n194), .Y(n195) );
  XNOR2X2 U262 ( .A(n177), .B(n176), .Y(PRODUCT[30]) );
  OAI21XL U263 ( .A0(n202), .A1(n172), .B0(n171), .Y(n177) );
  INVXL U264 ( .A(n1131), .Y(n1084) );
  INVXL U265 ( .A(n1126), .Y(n1116) );
  OAI22X1 U266 ( .A0(n818), .A1(n529), .B0(n817), .B1(n102), .Y(n854) );
  XNOR2XL U267 ( .A(B[7]), .B(A[9]), .Y(n902) );
  XNOR2XL U268 ( .A(B[7]), .B(n858), .Y(n833) );
  XNOR2XL U269 ( .A(B[8]), .B(A[9]), .Y(n903) );
  OAI22X1 U270 ( .A0(n391), .A1(n528), .B0(n390), .B1(n7), .Y(n397) );
  INVXL U271 ( .A(n1071), .Y(n1073) );
  NAND2XL U272 ( .A(n1101), .B(n1103), .Y(n1106) );
  XNOR2X1 U273 ( .A(B[26]), .B(A[11]), .Y(n97) );
  XNOR2XL U274 ( .A(B[25]), .B(A[9]), .Y(n502) );
  XNOR2X1 U275 ( .A(B[25]), .B(A[7]), .Y(n519) );
  XNOR2XL U276 ( .A(B[18]), .B(A[15]), .Y(n510) );
  OAI22X1 U277 ( .A0(n529), .A1(n563), .B0(n571), .B1(n102), .Y(n577) );
  XOR2X1 U278 ( .A(B[11]), .B(n73), .Y(n675) );
  OAI22X1 U279 ( .A0(n791), .A1(n884), .B0(n829), .B1(n882), .Y(n819) );
  XNOR2XL U280 ( .A(B[9]), .B(n9), .Y(n297) );
  XNOR2XL U281 ( .A(B[26]), .B(A[9]), .Y(n487) );
  INVX1 U282 ( .A(n385), .Y(n464) );
  XNOR2XL U283 ( .A(B[24]), .B(A[11]), .Y(n495) );
  XNOR2XL U284 ( .A(B[23]), .B(A[11]), .Y(n503) );
  AOI21XL U285 ( .A0(n170), .A1(n160), .B0(n159), .Y(n161) );
  INVX1 U286 ( .A(n114), .Y(n238) );
  OAI22XL U287 ( .A0(n353), .A1(n499), .B0(n352), .B1(n8), .Y(n365) );
  NAND2X1 U288 ( .A(n71), .B(n186), .Y(n192) );
  OAI21XL U289 ( .A0(n202), .A1(n179), .B0(n178), .Y(n183) );
  NAND2XL U290 ( .A(n1103), .B(n1108), .Y(n1065) );
  INVXL U291 ( .A(n1032), .Y(n1033) );
  NOR2XL U292 ( .A(n1134), .B(n1133), .Y(n1071) );
  XNOR2XL U293 ( .A(n1132), .B(n1130), .Y(PRODUCT[11]) );
  OAI22XL U294 ( .A0(n340), .A1(n499), .B0(n353), .B1(n8), .Y(n356) );
  XNOR2XL U295 ( .A(B[8]), .B(A[3]), .Y(n342) );
  OAI22XL U296 ( .A0(n276), .A1(n486), .B0(n307), .B1(n485), .Y(n310) );
  NAND2BXL U297 ( .AN(n986), .B(A[3]), .Y(n399) );
  OAI22XL U298 ( .A0(n392), .A1(n528), .B0(n391), .B1(n7), .Y(n427) );
  XNOR2XL U299 ( .A(B[10]), .B(A[1]), .Y(n349) );
  NOR2XL U300 ( .A(n1065), .B(n1071), .Y(n1060) );
  XOR2XL U301 ( .A(n1082), .B(n1081), .Y(PRODUCT[13]) );
  NAND2XL U302 ( .A(n1122), .B(n1128), .Y(n1081) );
  XNOR2XL U303 ( .A(n1084), .B(n1083), .Y(PRODUCT[12]) );
  NAND2XL U304 ( .A(n1123), .B(n1129), .Y(n1083) );
  INVXL U305 ( .A(n100), .Y(n101) );
  XNOR2XL U306 ( .A(B[23]), .B(A[7]), .Y(n568) );
  XNOR2XL U307 ( .A(B[22]), .B(A[7]), .Y(n587) );
  XNOR2XL U308 ( .A(B[24]), .B(A[3]), .Y(n616) );
  OAI22X1 U309 ( .A0(n615), .A1(n102), .B0(n613), .B1(n529), .Y(n621) );
  XNOR2X1 U310 ( .A(B[25]), .B(A[1]), .Y(n648) );
  XOR2X1 U311 ( .A(B[14]), .B(n59), .Y(n664) );
  INVXL U312 ( .A(n858), .Y(n59) );
  OAI22X1 U313 ( .A0(n674), .A1(n529), .B0(n694), .B1(n102), .Y(n692) );
  OAI22X1 U314 ( .A0(n747), .A1(n258), .B0(n702), .B1(n257), .Y(n737) );
  XNOR2XL U315 ( .A(B[10]), .B(n856), .Y(n719) );
  XNOR2X1 U316 ( .A(B[15]), .B(A[7]), .Y(n740) );
  XNOR2XL U317 ( .A(B[13]), .B(A[9]), .Y(n748) );
  CMPR22X1 U318 ( .A(n767), .B(n768), .CO(n777), .S(n799) );
  OAI22X1 U319 ( .A0(n741), .A1(n529), .B0(n742), .B1(n102), .Y(n768) );
  XNOR2XL U320 ( .A(B[8]), .B(n858), .Y(n821) );
  XNOR2XL U321 ( .A(B[15]), .B(A[3]), .Y(n890) );
  INVX1 U322 ( .A(n41), .Y(n42) );
  CMPR22X1 U323 ( .A(n831), .B(n830), .CO(n840), .S(n861) );
  OAI22X1 U324 ( .A0(n814), .A1(n529), .B0(n818), .B1(n102), .Y(n831) );
  XNOR2XL U325 ( .A(B[9]), .B(A[9]), .Y(n863) );
  XNOR2XL U326 ( .A(B[10]), .B(n895), .Y(n911) );
  OAI22XL U327 ( .A0(n903), .A1(n486), .B0(n902), .B1(n485), .Y(n912) );
  XNOR2XL U328 ( .A(B[8]), .B(n9), .Y(n296) );
  OAI22XL U329 ( .A0(n277), .A1(n486), .B0(n276), .B1(n485), .Y(n295) );
  OAI22X1 U330 ( .A0(n930), .A1(n499), .B0(n283), .B1(n8), .Y(n956) );
  OAI22X1 U331 ( .A0(n821), .A1(n257), .B0(n833), .B1(n258), .Y(n838) );
  XNOR2XL U332 ( .A(B[18]), .B(A[1]), .Y(n853) );
  XNOR2XL U333 ( .A(B[1]), .B(A[1]), .Y(n404) );
  OAI22XL U334 ( .A0(n418), .A1(n892), .B0(n408), .B1(n369), .Y(n413) );
  OAI22XL U335 ( .A0(n419), .A1(n892), .B0(n418), .B1(n369), .Y(n420) );
  OAI22XL U336 ( .A0(n402), .A1(n328), .B0(n401), .B1(n329), .Y(n415) );
  CMPR32X1 U337 ( .A(n376), .B(n375), .C(n374), .CO(n454), .S(n450) );
  OAI22XL U338 ( .A0(n370), .A1(n892), .B0(n381), .B1(n369), .Y(n375) );
  OAI21XL U339 ( .A0(n453), .A1(n461), .B0(n452), .Y(n460) );
  NAND2XL U340 ( .A(n464), .B(n1053), .Y(n453) );
  AOI21XL U341 ( .A0(n464), .A1(n462), .B0(n451), .Y(n452) );
  AOI2BB1X2 U342 ( .A0N(n566), .A1N(n884), .B0(n66), .Y(n65) );
  INVXL U343 ( .A(n97), .Y(n96) );
  XNOR2XL U344 ( .A(B[23]), .B(A[13]), .Y(n482) );
  OAI22XL U345 ( .A0(n525), .A1(n258), .B0(n503), .B1(n257), .Y(n512) );
  OAI22XL U346 ( .A0(n510), .A1(n102), .B0(n1045), .B1(n529), .Y(n514) );
  XNOR2XL U347 ( .A(B[23]), .B(A[9]), .Y(n543) );
  OAI22XL U348 ( .A0(n565), .A1(n884), .B0(n589), .B1(n882), .Y(n627) );
  OR2XL U349 ( .A(n603), .B(n602), .Y(n631) );
  INVX1 U350 ( .A(n45), .Y(n46) );
  OAI22XL U351 ( .A0(n604), .A1(n99), .B0(n589), .B1(n884), .Y(n612) );
  CMPR32X1 U352 ( .A(n746), .B(n745), .C(n744), .CO(n736), .S(n758) );
  OAI22XL U353 ( .A0(n739), .A1(n7), .B0(n717), .B1(n528), .Y(n745) );
  OAI22XL U354 ( .A0(n822), .A1(n369), .B0(n788), .B1(n934), .Y(n825) );
  OAI22XL U355 ( .A0(n297), .A1(n7), .B0(n933), .B1(n528), .Y(n965) );
  OAI22XL U356 ( .A0(n404), .A1(n892), .B0(n986), .B1(n369), .Y(n1095) );
  NAND2XL U357 ( .A(n369), .B(n405), .Y(n1094) );
  NOR2XL U358 ( .A(n407), .B(n406), .Y(n1090) );
  NAND2XL U359 ( .A(n407), .B(n406), .Y(n1091) );
  NAND2XL U360 ( .A(n1095), .B(n1094), .Y(n1096) );
  NAND2XL U361 ( .A(n413), .B(n412), .Y(n1098) );
  NAND2XL U362 ( .A(n421), .B(n420), .Y(n1112) );
  AOI21XL U363 ( .A0(n1099), .A1(n411), .B0(n414), .Y(n1114) );
  INVXL U364 ( .A(n1098), .Y(n414) );
  NAND2XL U365 ( .A(n436), .B(n435), .Y(n1086) );
  INVXL U366 ( .A(n460), .Y(n1023) );
  OAI2BB1XL U367 ( .A0N(n486), .A1N(n485), .B0(n484), .Y(n494) );
  OAI22XL U368 ( .A0(n489), .A1(n257), .B0(n495), .B1(n258), .Y(n493) );
  INVXL U369 ( .A(n487), .Y(n484) );
  ADDFX2 U370 ( .A(n478), .B(n477), .CI(n476), .CO(mult_x_1_n407), .S(
        mult_x_1_n408) );
  OAI22XL U371 ( .A0(n474), .A1(n102), .B0(n470), .B1(n529), .Y(n478) );
  AOI21XL U372 ( .A0(n1122), .A1(n1080), .B0(n78), .Y(n79) );
  NAND2BXL U373 ( .AN(n986), .B(A[9]), .Y(n304) );
  NAND2X1 U374 ( .A(n90), .B(n89), .Y(n109) );
  OAI21XL U375 ( .A0(n205), .A1(n215), .B0(n216), .Y(n206) );
  AOI21XL U376 ( .A0(n170), .A1(n181), .B0(n169), .Y(n171) );
  NAND2XL U377 ( .A(n137), .B(n136), .Y(n174) );
  NAND2XL U378 ( .A(n1001), .B(n1000), .Y(n1003) );
  NOR2XL U379 ( .A(n1015), .B(n1011), .Y(n193) );
  NOR2X1 U380 ( .A(n137), .B(n136), .Y(n173) );
  NAND2XL U381 ( .A(n1008), .B(n1007), .Y(n1032) );
  INVXL U382 ( .A(n1003), .Y(n1034) );
  INVXL U383 ( .A(n1065), .Y(n1068) );
  INVXL U384 ( .A(n1056), .Y(n1102) );
  XNOR2XL U385 ( .A(B[2]), .B(n895), .Y(n353) );
  XNOR2XL U386 ( .A(B[3]), .B(n895), .Y(n340) );
  XNOR2XL U387 ( .A(B[1]), .B(A[15]), .Y(n817) );
  CMPR22X1 U388 ( .A(n881), .B(n880), .CO(n855), .S(n898) );
  OAI22X1 U389 ( .A0(n815), .A1(n529), .B0(n102), .B1(n51), .Y(n881) );
  OAI22X1 U390 ( .A0(n817), .A1(n529), .B0(n816), .B1(n102), .Y(n880) );
  NAND2BXL U391 ( .AN(n986), .B(A[15]), .Y(n815) );
  NAND2BXL U392 ( .AN(n986), .B(n9), .Y(n389) );
  XNOR2XL U393 ( .A(B[4]), .B(n9), .Y(n364) );
  XNOR2XL U394 ( .A(B[3]), .B(n9), .Y(n379) );
  NAND2XL U395 ( .A(n1041), .B(n1040), .Y(n1056) );
  INVXL U396 ( .A(n163), .Y(n165) );
  OAI21XL U397 ( .A0(n153), .A1(n202), .B0(n152), .Y(n158) );
  INVXL U398 ( .A(n154), .Y(n156) );
  NAND2XL U399 ( .A(n133), .B(n193), .Y(n179) );
  OAI21XL U400 ( .A0(n188), .A1(n197), .B0(n189), .Y(n132) );
  AOI21XL U401 ( .A0(n1102), .A1(n1108), .B0(n1058), .Y(n1066) );
  INVXL U402 ( .A(n1107), .Y(n1058) );
  AOI21XL U403 ( .A0(n1104), .A1(n1068), .B0(n1067), .Y(n1069) );
  INVXL U404 ( .A(n1066), .Y(n1067) );
  NAND2XL U405 ( .A(n1101), .B(n1068), .Y(n1070) );
  NAND2XL U406 ( .A(n1134), .B(n1133), .Y(n1072) );
  NAND2XL U407 ( .A(n1057), .B(n1135), .Y(n1107) );
  AOI21XL U408 ( .A0(n1104), .A1(n1103), .B0(n1102), .Y(n1105) );
  INVX1 U409 ( .A(n1129), .Y(n1080) );
  NOR2BXL U410 ( .AN(n986), .B(n832), .Y(n326) );
  XNOR2XL U411 ( .A(B[12]), .B(A[15]), .Y(n613) );
  XNOR2XL U412 ( .A(B[11]), .B(A[15]), .Y(n615) );
  XNOR2XL U413 ( .A(B[10]), .B(A[15]), .Y(n651) );
  XNOR2XL U414 ( .A(B[9]), .B(A[15]), .Y(n674) );
  XNOR2XL U415 ( .A(B[8]), .B(A[15]), .Y(n694) );
  XOR2XL U416 ( .A(B[5]), .B(n73), .Y(n829) );
  XOR2XL U417 ( .A(B[4]), .B(n51), .Y(n790) );
  XNOR2XL U418 ( .A(B[3]), .B(A[9]), .Y(n276) );
  NOR2BXL U419 ( .AN(n986), .B(n884), .Y(n280) );
  OAI22XL U420 ( .A0(n266), .A1(n257), .B0(n261), .B1(n258), .Y(n278) );
  XNOR2XL U421 ( .A(B[2]), .B(A[1]), .Y(n408) );
  XNOR2XL U422 ( .A(B[3]), .B(A[1]), .Y(n418) );
  XNOR2XL U423 ( .A(B[9]), .B(A[1]), .Y(n370) );
  OAI22XL U424 ( .A0(n354), .A1(n328), .B0(n368), .B1(n329), .Y(n372) );
  CMPR32X1 U425 ( .A(n337), .B(n336), .C(n335), .CO(n332), .S(n995) );
  OAI22XL U426 ( .A0(n308), .A1(n528), .B0(n327), .B1(n7), .Y(n336) );
  OAI22XL U427 ( .A0(n349), .A1(n369), .B0(n331), .B1(n934), .Y(n346) );
  OAI22XL U428 ( .A0(n330), .A1(n328), .B0(n342), .B1(n329), .Y(n347) );
  XNOR2XL U429 ( .A(B[21]), .B(A[9]), .Y(n559) );
  XNOR2XL U430 ( .A(B[24]), .B(A[7]), .Y(n539) );
  XNOR2XL U431 ( .A(B[26]), .B(A[3]), .Y(n564) );
  OAI22XL U432 ( .A0(n601), .A1(n7), .B0(n570), .B1(n528), .Y(n632) );
  NAND2X1 U433 ( .A(n61), .B(n60), .Y(n602) );
  NAND2XL U434 ( .A(n573), .B(n892), .Y(n60) );
  XNOR2XL U435 ( .A(B[18]), .B(A[11]), .Y(n569) );
  XOR2XL U436 ( .A(B[14]), .B(n73), .Y(n604) );
  XNOR2XL U437 ( .A(B[20]), .B(A[7]), .Y(n638) );
  XNOR2XL U438 ( .A(B[16]), .B(A[9]), .Y(n652) );
  XNOR2XL U439 ( .A(B[24]), .B(A[1]), .Y(n678) );
  CMPR22X1 U440 ( .A(n677), .B(n676), .CO(n679), .S(n696) );
  OAI22X1 U441 ( .A0(n674), .A1(n102), .B0(n651), .B1(n529), .Y(n677) );
  OAI22X1 U442 ( .A0(n652), .A1(n486), .B0(n700), .B1(n485), .Y(n676) );
  XNOR2XL U443 ( .A(B[20]), .B(A[3]), .Y(n729) );
  XNOR2XL U444 ( .A(B[8]), .B(n856), .Y(n766) );
  XNOR2XL U445 ( .A(n264), .B(A[12]), .Y(n52) );
  OAI22XL U446 ( .A0(n894), .A1(n329), .B0(n890), .B1(n328), .Y(n905) );
  XNOR2XL U447 ( .A(B[12]), .B(n9), .Y(n889) );
  CMPR32X1 U448 ( .A(n322), .B(n321), .C(n320), .CO(n312), .S(n992) );
  XNOR2XL U449 ( .A(B[11]), .B(A[3]), .Y(n269) );
  XNOR2XL U450 ( .A(B[10]), .B(n9), .Y(n933) );
  XNOR2XL U451 ( .A(B[15]), .B(A[1]), .Y(n935) );
  OAI22XL U452 ( .A0(n902), .A1(n267), .B0(n879), .B1(n485), .Y(n940) );
  OAI22XL U453 ( .A0(n863), .A1(n486), .B0(n903), .B1(n485), .Y(n915) );
  OAI22XL U454 ( .A0(n408), .A1(n892), .B0(n404), .B1(n369), .Y(n407) );
  NOR2BXL U455 ( .AN(n986), .B(n617), .Y(n406) );
  CMPR22X1 U456 ( .A(n410), .B(n409), .CO(n416), .S(n412) );
  OAI22XL U457 ( .A0(n431), .A1(n892), .B0(n430), .B1(n369), .Y(n440) );
  OAI22XL U458 ( .A0(n426), .A1(n328), .B0(n425), .B1(n329), .Y(n442) );
  XOR2XL U459 ( .A(n1064), .B(n1063), .Y(PRODUCT[39]) );
  OAI22XL U460 ( .A0(n717), .A1(n7), .B0(n699), .B1(n528), .Y(n722) );
  OAI22XL U461 ( .A0(n104), .A1(n288), .B0(n103), .B1(n102), .Y(n105) );
  OAI2BB1XL U462 ( .A0N(n884), .A1N(n99), .B0(n101), .Y(n107) );
  ADDFX2 U463 ( .A(n523), .B(n522), .CI(n521), .CO(n516), .S(n533) );
  OAI22XL U464 ( .A0(n531), .A1(n102), .B0(n510), .B1(n529), .Y(n522) );
  CMPR32X1 U465 ( .A(n670), .B(n669), .C(n668), .CO(n658), .S(n683) );
  OAI22XL U466 ( .A0(n641), .A1(n8), .B0(n638), .B1(n499), .Y(n669) );
  OAI22XL U467 ( .A0(n663), .A1(n7), .B0(n637), .B1(n528), .Y(n670) );
  OAI22XL U468 ( .A0(n662), .A1(n329), .B0(n616), .B1(n328), .Y(n655) );
  OAI22XL U469 ( .A0(n675), .A1(n99), .B0(n666), .B1(n884), .Y(n689) );
  CMPR32X1 U470 ( .A(n732), .B(n733), .C(n731), .CO(n708), .S(n760) );
  ADDFX2 U471 ( .A(n38), .B(n771), .CI(n770), .CO(n759), .S(n783) );
  OAI22XL U472 ( .A0(n743), .A1(n7), .B0(n739), .B1(n528), .Y(n771) );
  OAI22XL U473 ( .A0(n728), .A1(n99), .B0(n719), .B1(n884), .Y(n752) );
  CMPR32X1 U474 ( .A(n797), .B(n796), .C(n795), .CO(n784), .S(n808) );
  OAI22XL U475 ( .A0(n794), .A1(n257), .B0(n821), .B1(n258), .Y(n826) );
  OAI22XL U476 ( .A0(n863), .A1(n485), .B0(n836), .B1(n486), .Y(n909) );
  XOR2XL U477 ( .A(n50), .B(n840), .Y(n907) );
  OAI22XL U478 ( .A0(n931), .A1(n8), .B0(n911), .B1(n499), .Y(n952) );
  OAI22XL U479 ( .A0(n937), .A1(n329), .B0(n894), .B1(n328), .Y(n953) );
  OAI22XL U480 ( .A0(n298), .A1(n573), .B0(n936), .B1(n892), .Y(n976) );
  INVX1 U481 ( .A(n976), .Y(n57) );
  ADDFX2 U482 ( .A(n301), .B(n300), .CI(n299), .CO(n975), .S(n319) );
  OAI22XL U483 ( .A0(n297), .A1(n528), .B0(n296), .B1(n7), .Y(n300) );
  ADDFX2 U484 ( .A(n979), .B(n978), .CI(n977), .CO(n970), .S(n980) );
  NAND2XL U485 ( .A(n959), .B(n958), .Y(n979) );
  NAND2XL U486 ( .A(n955), .B(n954), .Y(n959) );
  OAI22XL U487 ( .A0(n853), .A1(n369), .B0(n822), .B1(n934), .Y(n850) );
  OAI2BB1X1 U488 ( .A0N(n838), .A1N(n36), .B0(n72), .Y(n851) );
  NAND2XL U489 ( .A(n464), .B(n463), .Y(n465) );
  ADDFX2 U490 ( .A(n586), .B(n585), .CI(n584), .CO(mult_x_1_n463), .S(
        mult_x_1_n464) );
  OAI2BB1XL U491 ( .A0N(n63), .A1N(n579), .B0(n62), .Y(n585) );
  NAND2XL U492 ( .A(n64), .B(n65), .Y(n63) );
  XOR2X1 U493 ( .A(n77), .B(n598), .Y(mult_x_1_n474) );
  NAND2XL U494 ( .A(n1028), .B(n1027), .Y(mult_x_1_n310) );
  NAND2XL U495 ( .A(n1026), .B(n1025), .Y(mult_x_1_n81) );
  INVXL U496 ( .A(n1024), .Y(n1026) );
  OAI22XL U497 ( .A0(n470), .A1(n102), .B0(n103), .B1(n529), .Y(n469) );
  INVXL U498 ( .A(n475), .Y(n479) );
  OAI22XL U499 ( .A0(n1046), .A1(n99), .B0(n482), .B1(n884), .Y(n492) );
  OAI22XL U500 ( .A0(n1044), .A1(n102), .B0(n483), .B1(n529), .Y(n491) );
  OAI22XL U501 ( .A0(n503), .A1(n258), .B0(n495), .B1(n257), .Y(n506) );
  INVXL U502 ( .A(n1048), .Y(n1049) );
  OAI22XL U503 ( .A0(n1045), .A1(n102), .B0(n1044), .B1(n529), .Y(n1051) );
  OAI22XL U504 ( .A0(n1047), .A1(n99), .B0(n1046), .B1(n884), .Y(n1050) );
  CMPR32X1 U505 ( .A(n537), .B(n536), .C(n535), .CO(mult_x_1_n443), .S(n532)
         );
  NAND2X1 U506 ( .A(n600), .B(n599), .Y(n75) );
  ADDFX2 U507 ( .A(n636), .B(n635), .CI(n634), .CO(mult_x_1_n487), .S(
        mult_x_1_n488) );
  ADDFX2 U508 ( .A(n982), .B(n981), .CI(n980), .CO(mult_x_1_n665), .S(
        mult_x_1_n666) );
  OAI2BB1X1 U509 ( .A0N(n55), .A1N(n975), .B0(n53), .Y(n981) );
  NAND2XL U510 ( .A(n58), .B(n57), .Y(n55) );
  NAND2XL U511 ( .A(n54), .B(n976), .Y(n53) );
  ADDFX2 U512 ( .A(n869), .B(n868), .CI(n867), .CO(mult_x_1_n611), .S(
        mult_x_1_n612) );
  NOR2BXL U513 ( .AN(n986), .B(n934), .Y(n1220) );
  XOR2XL U514 ( .A(n1093), .B(n1096), .Y(n1218) );
  NAND2XL U515 ( .A(n1092), .B(n1091), .Y(n1093) );
  INVXL U516 ( .A(n1090), .Y(n1092) );
  NAND2XL U517 ( .A(n411), .B(n1098), .Y(n1100) );
  NAND2XL U518 ( .A(n1113), .B(n1112), .Y(n1115) );
  INVXL U519 ( .A(n1111), .Y(n1113) );
  NAND2XL U520 ( .A(n403), .B(n1119), .Y(n1121) );
  NAND2XL U521 ( .A(n1087), .B(n1086), .Y(n1089) );
  NAND2XL U522 ( .A(n1053), .B(n1052), .Y(n1054) );
  CLKINVX3 U523 ( .A(A[5]), .Y(n74) );
  OR2X2 U524 ( .A(n839), .B(n840), .Y(n36) );
  INVX1 U525 ( .A(A[15]), .Y(n51) );
  INVXL U526 ( .A(n772), .Y(n37) );
  XOR2X1 U527 ( .A(B[13]), .B(n51), .Y(n571) );
  NAND2BX1 U528 ( .AN(n187), .B(n1014), .Y(n71) );
  AOI21X1 U529 ( .A0(n1014), .A1(n1013), .B0(n68), .Y(n67) );
  XNOR2X1 U530 ( .A(B[6]), .B(A[15]), .Y(n741) );
  XNOR2X1 U531 ( .A(B[6]), .B(A[9]), .Y(n879) );
  OAI22X1 U532 ( .A0(n773), .A1(n8), .B0(n740), .B1(n499), .Y(n778) );
  CMPR22X1 U533 ( .A(n692), .B(n691), .CO(n697), .S(n733) );
  OAI22X1 U534 ( .A0(n590), .A1(n258), .B0(n569), .B1(n257), .Y(n633) );
  CMPR22X1 U535 ( .A(n398), .B(n397), .CO(n428), .S(n434) );
  OAI22X1 U536 ( .A0(n389), .A1(n528), .B0(n7), .B1(n74), .Y(n398) );
  OAI22X1 U537 ( .A0(n49), .A1(n257), .B0(n664), .B1(n258), .Y(n649) );
  INVXL U538 ( .A(n594), .Y(n39) );
  INVX1 U539 ( .A(n39), .Y(n40) );
  INVXL U540 ( .A(n862), .Y(n41) );
  OAI22X1 U541 ( .A0(n489), .A1(n258), .B0(n97), .B1(n257), .Y(n475) );
  ADDFX2 U542 ( .A(n107), .B(n106), .CI(n105), .S(n997) );
  CMPR22X1 U543 ( .A(n855), .B(n854), .CO(n830), .S(n901) );
  INVXL U544 ( .A(n905), .Y(n43) );
  INVX1 U545 ( .A(n43), .Y(n44) );
  ADDFX2 U546 ( .A(n558), .B(n557), .CI(n556), .CO(n552), .S(n576) );
  OAI22X1 U547 ( .A0(n936), .A1(n369), .B0(n935), .B1(n934), .Y(n974) );
  XOR2X1 U548 ( .A(n838), .B(n839), .Y(n50) );
  OAI22X2 U549 ( .A0(n569), .A1(n258), .B0(n560), .B1(n257), .Y(n593) );
  INVXL U550 ( .A(n973), .Y(n47) );
  INVX1 U551 ( .A(n47), .Y(n48) );
  OAI22X1 U552 ( .A0(n932), .A1(n7), .B0(n889), .B1(n528), .Y(n944) );
  OAI22X1 U553 ( .A0(n889), .A1(n7), .B0(n888), .B1(n528), .Y(n906) );
  CLKINVX3 U554 ( .A(n488), .Y(n858) );
  OAI22X1 U555 ( .A0(n519), .A1(n8), .B0(n500), .B1(n499), .Y(n511) );
  OAI22X1 U556 ( .A0(n618), .A1(n617), .B0(n616), .B1(n329), .Y(n630) );
  XOR2X2 U557 ( .A(n67), .B(n1018), .Y(PRODUCT[26]) );
  NAND2X1 U558 ( .A(n210), .B(n209), .Y(n211) );
  XOR2X2 U559 ( .A(n219), .B(n218), .Y(PRODUCT[23]) );
  NAND2X1 U560 ( .A(n224), .B(n223), .Y(n225) );
  XNOR2X2 U561 ( .A(n183), .B(n182), .Y(PRODUCT[29]) );
  NAND2X1 U562 ( .A(n190), .B(n189), .Y(n191) );
  XNOR2X2 U563 ( .A(n200), .B(n199), .Y(PRODUCT[27]) );
  OAI22X1 U564 ( .A0(n640), .A1(n486), .B0(n652), .B1(n485), .Y(n672) );
  OAI22X1 U565 ( .A0(n836), .A1(n485), .B0(n802), .B1(n486), .Y(n848) );
  OAI22X1 U566 ( .A0(n614), .A1(n257), .B0(n49), .B1(n258), .Y(n620) );
  OAI22X1 U567 ( .A0(n886), .A1(n257), .B0(n287), .B1(n258), .Y(n929) );
  OAI22X1 U568 ( .A0(n675), .A1(n884), .B0(n99), .B1(n719), .Y(n691) );
  OAI22X1 U569 ( .A0(n666), .A1(n99), .B0(n639), .B1(n884), .Y(n673) );
  XNOR2XL U570 ( .A(B[25]), .B(A[15]), .Y(n104) );
  XNOR2XL U571 ( .A(B[20]), .B(A[15]), .Y(n1044) );
  XNOR2XL U572 ( .A(B[19]), .B(A[15]), .Y(n1045) );
  OAI22X1 U573 ( .A0(n648), .A1(n892), .B0(n678), .B1(n369), .Y(n681) );
  XNOR2XL U574 ( .A(B[24]), .B(A[9]), .Y(n524) );
  XNOR2XL U575 ( .A(B[17]), .B(A[9]), .Y(n640) );
  XNOR2X1 U576 ( .A(B[15]), .B(A[9]), .Y(n700) );
  NAND2X4 U577 ( .A(n52), .B(n884), .Y(n882) );
  XOR2X1 U578 ( .A(n975), .B(n56), .Y(n983) );
  XNOR2X1 U579 ( .A(B[15]), .B(n856), .Y(n589) );
  NAND2BXL U580 ( .AN(n65), .B(n580), .Y(n62) );
  INVXL U581 ( .A(n580), .Y(n64) );
  XNOR3X2 U582 ( .A(n580), .B(n65), .C(n579), .Y(n596) );
  NOR2X1 U583 ( .A(n565), .B(n882), .Y(n66) );
  NAND2X1 U584 ( .A(n214), .B(n123), .Y(n70) );
  AOI21X4 U585 ( .A0(n114), .A1(n113), .B0(n112), .Y(n204) );
  XNOR2X1 U586 ( .A(B[23]), .B(A[1]), .Y(n693) );
  XOR2X1 U587 ( .A(B[14]), .B(n51), .Y(n563) );
  OAI21XL U588 ( .A0(n250), .A1(n1127), .B0(n251), .Y(n81) );
  NAND2XL U589 ( .A(n1198), .B(n1197), .Y(n251) );
  NOR2X1 U590 ( .A(n1198), .B(n1197), .Y(n250) );
  CLKINVX3 U591 ( .A(n1014), .Y(n202) );
  OAI22X1 U592 ( .A0(n563), .A1(n102), .B0(n562), .B1(n529), .Y(n578) );
  XNOR2X1 U593 ( .A(B[15]), .B(A[15]), .Y(n562) );
  OAI22X1 U594 ( .A0(n699), .A1(n7), .B0(n663), .B1(n528), .Y(n705) );
  OAI22X1 U595 ( .A0(n648), .A1(n369), .B0(n605), .B1(n934), .Y(n646) );
  NOR2X1 U596 ( .A(n131), .B(n130), .Y(n188) );
  ADDFHX4 U597 ( .A(n1182), .B(n1183), .CI(n1181), .CO(n117), .S(n116) );
  XOR2X1 U598 ( .A(B[6]), .B(n73), .Y(n791) );
  OAI2BB1XL U599 ( .A0N(n76), .A1N(n598), .B0(n75), .Y(mult_x_1_n473) );
  OR2X2 U600 ( .A(n600), .B(n599), .Y(n76) );
  CMPR22X1 U601 ( .A(n621), .B(n620), .CO(n628), .S(n654) );
  OAI22X1 U602 ( .A0(n729), .A1(n329), .B0(n716), .B1(n617), .Y(n746) );
  XNOR2X1 U603 ( .A(B[21]), .B(A[3]), .Y(n716) );
  XNOR2X1 U604 ( .A(B[6]), .B(A[3]), .Y(n368) );
  XNOR2X1 U605 ( .A(B[7]), .B(A[3]), .Y(n354) );
  OAI22X1 U606 ( .A0(n748), .A1(n485), .B0(n718), .B1(n486), .Y(n753) );
  XNOR2X1 U607 ( .A(B[14]), .B(A[9]), .Y(n718) );
  NOR2X1 U608 ( .A(n168), .B(n173), .Y(n160) );
  XNOR2X2 U609 ( .A(n234), .B(n233), .Y(PRODUCT[19]) );
  OAI21XL U610 ( .A0(n173), .A1(n180), .B0(n174), .Y(n159) );
  AOI21X1 U611 ( .A0(n207), .A1(n230), .B0(n206), .Y(n212) );
  XNOR2X1 U612 ( .A(B[26]), .B(n9), .Y(n538) );
  XNOR2X1 U613 ( .A(B[21]), .B(A[5]), .Y(n663) );
  XNOR2X1 U614 ( .A(B[17]), .B(n856), .Y(n566) );
  OAI22X1 U615 ( .A0(n587), .A1(n8), .B0(n568), .B1(n499), .Y(n579) );
  OAI22X1 U616 ( .A0(n702), .A1(n258), .B0(n701), .B1(n257), .Y(n725) );
  XNOR2X1 U617 ( .A(B[13]), .B(n858), .Y(n701) );
  OAI22X1 U618 ( .A0(n764), .A1(n329), .B0(n729), .B1(n617), .Y(n755) );
  AOI21X1 U619 ( .A0(n82), .A1(n249), .B0(n81), .Y(n239) );
  ADDFHX1 U620 ( .A(n1160), .B(n1158), .CI(n1157), .CO(n136), .S(n135) );
  OAI22X1 U621 ( .A0(n765), .A1(n884), .B0(n791), .B1(n882), .Y(n792) );
  AOI21XL U622 ( .A0(n1035), .A1(n1034), .B0(n1033), .Y(n1036) );
  OAI22X2 U623 ( .A0(n352), .A1(n499), .B0(n351), .B1(n8), .Y(n377) );
  NOR2XL U624 ( .A(n250), .B(n1126), .Y(n82) );
  NAND2XL U625 ( .A(n1122), .B(n1123), .Y(n80) );
  INVXL U626 ( .A(n1128), .Y(n78) );
  OAI21XL U627 ( .A0(n1131), .A1(n80), .B0(n79), .Y(n249) );
  NOR2XL U628 ( .A(n1193), .B(n1194), .Y(n83) );
  INVXL U629 ( .A(n83), .Y(n242) );
  OR2X2 U630 ( .A(n1195), .B(n1196), .Y(n246) );
  NAND2XL U631 ( .A(n242), .B(n246), .Y(n86) );
  NAND2XL U632 ( .A(n1195), .B(n1196), .Y(n245) );
  INVXL U633 ( .A(n245), .Y(n240) );
  NAND2XL U634 ( .A(n1193), .B(n1194), .Y(n241) );
  INVXL U635 ( .A(n241), .Y(n84) );
  AOI21XL U636 ( .A0(n242), .A1(n240), .B0(n84), .Y(n85) );
  OAI21X2 U637 ( .A0(n239), .A1(n86), .B0(n85), .Y(n114) );
  NOR2XL U638 ( .A(n1190), .B(n1192), .Y(n231) );
  NAND2XL U639 ( .A(n1190), .B(n1192), .Y(n235) );
  INVXL U640 ( .A(n235), .Y(n88) );
  OAI21XL U641 ( .A0(n238), .A1(n108), .B0(n111), .Y(n93) );
  INVXL U642 ( .A(n110), .Y(n91) );
  XNOR2XL U643 ( .A(B[23]), .B(A[15]), .Y(n470) );
  XNOR2XL U644 ( .A(A[13]), .B(A[14]), .Y(n288) );
  XOR2XL U645 ( .A(A[15]), .B(A[14]), .Y(n94) );
  XNOR2X1 U646 ( .A(B[24]), .B(A[15]), .Y(n103) );
  XNOR2X1 U647 ( .A(B[25]), .B(A[13]), .Y(n98) );
  XNOR2X2 U648 ( .A(A[11]), .B(A[12]), .Y(n884) );
  XNOR2X1 U649 ( .A(B[26]), .B(A[13]), .Y(n100) );
  OAI22X1 U650 ( .A0(n98), .A1(n99), .B0(n100), .B1(n884), .Y(n106) );
  INVXL U651 ( .A(n106), .Y(n468) );
  XNOR2XL U652 ( .A(A[9]), .B(A[10]), .Y(n832) );
  XOR2XL U653 ( .A(A[11]), .B(A[10]), .Y(n95) );
  XNOR2X1 U654 ( .A(B[24]), .B(n856), .Y(n473) );
  OAI22XL U655 ( .A0(n98), .A1(n884), .B0(n473), .B1(n882), .Y(n471) );
  NAND2XL U656 ( .A(n998), .B(n997), .Y(mult_x_1_n100) );
  CMPR32X1 U657 ( .A(n1164), .B(n1165), .C(n1163), .CO(n130), .S(n129) );
  NOR2X1 U658 ( .A(n184), .B(n188), .Y(n133) );
  ADDFHX1 U659 ( .A(n1167), .B(n1168), .CI(n1166), .CO(n128), .S(n127) );
  NOR2X1 U660 ( .A(n127), .B(n126), .Y(n1015) );
  ADDFHX1 U661 ( .A(n1170), .B(n1171), .CI(n1169), .CO(n126), .S(n125) );
  ADDFHX1 U662 ( .A(n1161), .B(n1162), .CI(n1159), .CO(n134), .S(n131) );
  CMPR32X1 U663 ( .A(n1155), .B(n1156), .C(n1153), .CO(n138), .S(n137) );
  NOR2XL U664 ( .A(n163), .B(n154), .Y(n143) );
  NAND2XL U665 ( .A(n160), .B(n143), .Y(n144) );
  ADDFHX4 U666 ( .A(n1179), .B(n1180), .CI(n1178), .CO(n119), .S(n118) );
  NOR2X2 U667 ( .A(n108), .B(n110), .Y(n113) );
  NAND2X1 U668 ( .A(n118), .B(n117), .Y(n223) );
  NAND2XL U669 ( .A(n127), .B(n126), .Y(n1016) );
  NAND2XL U670 ( .A(n131), .B(n130), .Y(n189) );
  AOI21X2 U671 ( .A0(n133), .A1(n194), .B0(n132), .Y(n178) );
  NAND2XL U672 ( .A(n141), .B(n140), .Y(n155) );
  OAI21XL U673 ( .A0(n154), .A1(n164), .B0(n155), .Y(n142) );
  XOR2X2 U674 ( .A(n1029), .B(n147), .Y(PRODUCT[33]) );
  INVXL U675 ( .A(n160), .Y(n148) );
  NOR2XL U676 ( .A(n148), .B(n163), .Y(n151) );
  NAND2XL U677 ( .A(n151), .B(n11), .Y(n153) );
  INVXL U678 ( .A(n178), .Y(n170) );
  INVXL U679 ( .A(n159), .Y(n149) );
  OAI21XL U680 ( .A0(n149), .A1(n163), .B0(n164), .Y(n150) );
  AOI21XL U681 ( .A0(n170), .A1(n151), .B0(n150), .Y(n152) );
  NAND2X1 U682 ( .A(n156), .B(n155), .Y(n157) );
  XNOR2X4 U683 ( .A(n158), .B(n157), .Y(PRODUCT[32]) );
  NAND2XL U684 ( .A(n11), .B(n160), .Y(n162) );
  OAI21X1 U685 ( .A0(n202), .A1(n162), .B0(n161), .Y(n167) );
  NAND2X1 U686 ( .A(n165), .B(n164), .Y(n166) );
  NAND2XL U687 ( .A(n11), .B(n181), .Y(n172) );
  INVXL U688 ( .A(n180), .Y(n169) );
  INVXL U689 ( .A(n173), .Y(n175) );
  INVXL U690 ( .A(n184), .Y(n198) );
  NAND2XL U691 ( .A(n193), .B(n198), .Y(n187) );
  INVXL U692 ( .A(n197), .Y(n185) );
  AOI21XL U693 ( .A0(n194), .A1(n198), .B0(n185), .Y(n186) );
  INVXL U694 ( .A(n188), .Y(n190) );
  XNOR2X2 U695 ( .A(n192), .B(n191), .Y(PRODUCT[28]) );
  INVXL U696 ( .A(n193), .Y(n196) );
  INVXL U697 ( .A(n214), .Y(n203) );
  NOR2XL U698 ( .A(n203), .B(n215), .Y(n207) );
  CLKINVX3 U699 ( .A(n204), .Y(n230) );
  INVXL U700 ( .A(n213), .Y(n205) );
  INVXL U701 ( .A(n208), .Y(n210) );
  XOR2X2 U702 ( .A(n212), .B(n211), .Y(PRODUCT[24]) );
  INVXL U703 ( .A(n215), .Y(n217) );
  AOI21X1 U704 ( .A0(n230), .A1(n228), .B0(n221), .Y(n226) );
  INVXL U705 ( .A(n222), .Y(n224) );
  OAI21XL U706 ( .A0(n238), .A1(n231), .B0(n235), .Y(n234) );
  NAND2XL U707 ( .A(n236), .B(n235), .Y(n237) );
  XOR2X1 U708 ( .A(n238), .B(n237), .Y(PRODUCT[18]) );
  AOI21XL U709 ( .A0(n248), .A1(n246), .B0(n240), .Y(n244) );
  NAND2XL U710 ( .A(n242), .B(n241), .Y(n243) );
  XOR2X1 U711 ( .A(n244), .B(n243), .Y(PRODUCT[17]) );
  NAND2XL U712 ( .A(n246), .B(n245), .Y(n247) );
  INVXL U713 ( .A(n249), .Y(n1118) );
  OAI21XL U714 ( .A0(n1118), .A1(n1126), .B0(n1127), .Y(n254) );
  INVXL U715 ( .A(n250), .Y(n252) );
  NAND2XL U716 ( .A(n252), .B(n251), .Y(n253) );
  XOR2XL U717 ( .A(n9), .B(A[4]), .Y(n255) );
  XNOR2XL U718 ( .A(B[12]), .B(A[3]), .Y(n938) );
  OAI22XL U719 ( .A0(n269), .A1(n329), .B0(n938), .B1(n617), .Y(n964) );
  XNOR2X1 U720 ( .A(B[1]), .B(n858), .Y(n261) );
  XNOR2XL U721 ( .A(n986), .B(n858), .Y(n260) );
  XNOR2XL U722 ( .A(B[2]), .B(n858), .Y(n266) );
  XNOR2X1 U723 ( .A(B[7]), .B(n895), .Y(n283) );
  XOR2XL U724 ( .A(A[7]), .B(A[6]), .Y(n262) );
  OAI22XL U725 ( .A0(n283), .A1(n497), .B0(n282), .B1(n8), .Y(n271) );
  OAI22X2 U726 ( .A0(n263), .A1(n884), .B0(n882), .B1(n264), .Y(n290) );
  OAI22XL U727 ( .A0(n287), .A1(n257), .B0(n266), .B1(n258), .Y(n285) );
  XNOR2XL U728 ( .A(B[5]), .B(A[9]), .Y(n292) );
  XNOR2XL U729 ( .A(A[7]), .B(A[8]), .Y(n267) );
  XNOR2XL U730 ( .A(B[4]), .B(A[9]), .Y(n277) );
  XOR2XL U731 ( .A(A[9]), .B(A[8]), .Y(n268) );
  OAI22XL U732 ( .A0(n292), .A1(n486), .B0(n277), .B1(n485), .Y(n284) );
  XNOR2XL U733 ( .A(B[10]), .B(A[3]), .Y(n303) );
  OAI22XL U734 ( .A0(n303), .A1(n329), .B0(n269), .B1(n617), .Y(n314) );
  CMPR32X1 U735 ( .A(n272), .B(n271), .C(n270), .CO(n963), .S(n313) );
  XNOR2XL U736 ( .A(B[2]), .B(A[9]), .Y(n307) );
  XNOR2XL U737 ( .A(B[5]), .B(n895), .Y(n281) );
  XNOR2XL U738 ( .A(B[4]), .B(n895), .Y(n323) );
  OAI22XL U739 ( .A0(n281), .A1(n499), .B0(n323), .B1(n8), .Y(n309) );
  XNOR2X1 U740 ( .A(B[7]), .B(n9), .Y(n308) );
  OAI22XL U741 ( .A0(n296), .A1(n528), .B0(n308), .B1(n7), .Y(n321) );
  OAI22XL U742 ( .A0(n282), .A1(n499), .B0(n281), .B1(n8), .Y(n293) );
  XNOR2X1 U743 ( .A(B[13]), .B(A[1]), .Y(n298) );
  XNOR2XL U744 ( .A(B[14]), .B(A[1]), .Y(n936) );
  CLKINVX3 U745 ( .A(A[0]), .Y(n892) );
  CMPR32X1 U746 ( .A(n286), .B(n285), .C(n284), .CO(n957), .S(n270) );
  NOR2BX1 U747 ( .AN(n986), .B(n288), .Y(n878) );
  XNOR2XL U748 ( .A(B[2]), .B(n856), .Y(n883) );
  OAI22XL U749 ( .A0(n883), .A1(n884), .B0(n291), .B1(n882), .Y(n876) );
  OAI22XL U750 ( .A0(n879), .A1(n486), .B0(n292), .B1(n485), .Y(n927) );
  ADDFHX1 U751 ( .A(n295), .B(n294), .CI(n293), .CO(n301), .S(n320) );
  XNOR2XL U752 ( .A(B[12]), .B(A[1]), .Y(n302) );
  OAI22XL U753 ( .A0(n302), .A1(n369), .B0(n298), .B1(n934), .Y(n299) );
  XNOR2XL U754 ( .A(B[11]), .B(A[1]), .Y(n331) );
  OAI22XL U755 ( .A0(n331), .A1(n369), .B0(n302), .B1(n934), .Y(n334) );
  XNOR2X1 U756 ( .A(B[9]), .B(A[3]), .Y(n330) );
  OAI22XL U757 ( .A0(n330), .A1(n329), .B0(n303), .B1(n328), .Y(n333) );
  XNOR2XL U758 ( .A(n986), .B(A[9]), .Y(n305) );
  OAI22XL U759 ( .A0(n307), .A1(n486), .B0(n306), .B1(n485), .Y(n324) );
  CMPR32X1 U760 ( .A(n311), .B(n310), .C(n309), .CO(n322), .S(n335) );
  CMPR32X1 U761 ( .A(n314), .B(n313), .C(n312), .CO(n984), .S(n317) );
  NOR2XL U762 ( .A(n316), .B(n315), .Y(mult_x_1_n296) );
  CMPR32X1 U763 ( .A(n319), .B(n318), .C(n317), .CO(n315), .S(n988) );
  OAI22XL U764 ( .A0(n323), .A1(n499), .B0(n340), .B1(n8), .Y(n345) );
  ADDFHX1 U765 ( .A(n325), .B(n326), .CI(n324), .CO(n337), .S(n344) );
  XNOR2XL U766 ( .A(B[5]), .B(n9), .Y(n341) );
  OAI22XL U767 ( .A0(n327), .A1(n528), .B0(n341), .B1(n7), .Y(n343) );
  CMPR32X1 U768 ( .A(n334), .B(n333), .C(n332), .CO(n318), .S(n990) );
  NAND2XL U769 ( .A(n988), .B(n987), .Y(mult_x_1_n305) );
  OAI22XL U770 ( .A0(n341), .A1(n528), .B0(n364), .B1(n7), .Y(n355) );
  OAI22XL U771 ( .A0(n342), .A1(n328), .B0(n354), .B1(n329), .Y(n359) );
  ADDFHX1 U772 ( .A(n345), .B(n344), .CI(n343), .CO(n348), .S(n358) );
  CMPR32X1 U773 ( .A(n348), .B(n347), .C(n346), .CO(n991), .S(n993) );
  OAI22X1 U774 ( .A0(n370), .A1(n369), .B0(n349), .B1(n892), .Y(n363) );
  NOR2BX1 U775 ( .AN(n986), .B(n486), .Y(n367) );
  OAI22X2 U776 ( .A0(n350), .A1(n499), .B0(n8), .B1(n518), .Y(n378) );
  XNOR2XL U777 ( .A(B[1]), .B(n895), .Y(n352) );
  XNOR2XL U778 ( .A(n986), .B(n895), .Y(n351) );
  CMPR32X1 U779 ( .A(n6), .B(n356), .C(n355), .CO(n360), .S(n371) );
  CMPR32X1 U780 ( .A(n360), .B(n359), .C(n358), .CO(n994), .S(n361) );
  OAI22X1 U781 ( .A0(n364), .A1(n528), .B0(n379), .B1(n7), .Y(n384) );
  XNOR2XL U782 ( .A(B[5]), .B(A[3]), .Y(n380) );
  OAI22XL U783 ( .A0(n368), .A1(n328), .B0(n380), .B1(n329), .Y(n382) );
  XNOR2XL U784 ( .A(B[8]), .B(A[1]), .Y(n381) );
  CMPR32X1 U785 ( .A(n373), .B(n372), .C(n371), .CO(n362), .S(n374) );
  NOR2X1 U786 ( .A(n455), .B(n454), .Y(n1019) );
  NOR2XL U787 ( .A(n1024), .B(n1019), .Y(n459) );
  ADDHX2 U788 ( .A(n378), .B(n377), .CO(n366), .S(n396) );
  XNOR2XL U789 ( .A(B[2]), .B(n9), .Y(n392) );
  OAI22XL U790 ( .A0(n379), .A1(n528), .B0(n392), .B1(n7), .Y(n395) );
  XNOR2X1 U791 ( .A(B[4]), .B(A[3]), .Y(n426) );
  OAI22XL U792 ( .A0(n380), .A1(n328), .B0(n426), .B1(n329), .Y(n394) );
  XNOR2XL U793 ( .A(B[7]), .B(A[1]), .Y(n393) );
  OAI22XL U794 ( .A0(n381), .A1(n892), .B0(n393), .B1(n369), .Y(n387) );
  NOR2X1 U795 ( .A(n450), .B(n449), .Y(n385) );
  CMPR32X1 U796 ( .A(n388), .B(n387), .C(n386), .CO(n449), .S(n448) );
  XNOR2X1 U797 ( .A(B[1]), .B(n9), .Y(n391) );
  XNOR2X1 U798 ( .A(n986), .B(n9), .Y(n390) );
  XNOR2XL U799 ( .A(B[6]), .B(A[1]), .Y(n431) );
  OAI22XL U800 ( .A0(n393), .A1(n892), .B0(n431), .B1(n369), .Y(n438) );
  CMPR32X1 U801 ( .A(n396), .B(n395), .C(n394), .CO(n388), .S(n437) );
  OR2X2 U802 ( .A(n448), .B(n447), .Y(n1053) );
  XNOR2XL U803 ( .A(B[3]), .B(A[3]), .Y(n425) );
  XNOR2XL U804 ( .A(B[2]), .B(A[3]), .Y(n402) );
  OAI22XL U805 ( .A0(n425), .A1(n328), .B0(n402), .B1(n329), .Y(n433) );
  XNOR2XL U806 ( .A(B[5]), .B(A[1]), .Y(n430) );
  XNOR2XL U807 ( .A(B[4]), .B(A[1]), .Y(n419) );
  OAI22XL U808 ( .A0(n430), .A1(n892), .B0(n419), .B1(n369), .Y(n432) );
  OAI22X1 U809 ( .A0(n399), .A1(n328), .B0(n329), .B1(n19), .Y(n410) );
  XNOR2X1 U810 ( .A(B[1]), .B(A[3]), .Y(n401) );
  XNOR2XL U811 ( .A(n986), .B(A[3]), .Y(n400) );
  OAI22X1 U812 ( .A0(n401), .A1(n328), .B0(n400), .B1(n329), .Y(n409) );
  OAI21XL U813 ( .A0(n1090), .A1(n1096), .B0(n1091), .Y(n1099) );
  NOR2XL U814 ( .A(n421), .B(n420), .Y(n1111) );
  OAI21XL U815 ( .A0(n1114), .A1(n1111), .B0(n1112), .Y(n1120) );
  NAND2XL U816 ( .A(n423), .B(n422), .Y(n1119) );
  INVXL U817 ( .A(n1119), .Y(n424) );
  AOI21XL U818 ( .A0(n403), .A1(n1120), .B0(n424), .Y(n1088) );
  CMPR32X1 U819 ( .A(n429), .B(n428), .C(n427), .CO(n439), .S(n441) );
  CMPR32X1 U820 ( .A(n434), .B(n433), .C(n432), .CO(n435), .S(n423) );
  NOR2X1 U821 ( .A(n436), .B(n435), .Y(n1085) );
  OAI21XL U822 ( .A0(n1088), .A1(n1085), .B0(n1086), .Y(n1078) );
  CMPR32X1 U823 ( .A(n439), .B(n438), .C(n437), .CO(n447), .S(n445) );
  CMPR32X1 U824 ( .A(n442), .B(n441), .C(n440), .CO(n444), .S(n436) );
  NOR2XL U825 ( .A(n445), .B(n444), .Y(n443) );
  INVXL U826 ( .A(n443), .Y(n1077) );
  NAND2XL U827 ( .A(n445), .B(n444), .Y(n1076) );
  INVXL U828 ( .A(n1076), .Y(n446) );
  AOI21XL U829 ( .A0(n1078), .A1(n1077), .B0(n446), .Y(n461) );
  NAND2XL U830 ( .A(n448), .B(n447), .Y(n1052) );
  INVXL U831 ( .A(n1052), .Y(n462) );
  NAND2XL U832 ( .A(n450), .B(n449), .Y(n463) );
  INVXL U833 ( .A(n463), .Y(n451) );
  OAI21XL U834 ( .A0(n1024), .A1(n1020), .B0(n1025), .Y(n458) );
  AOI21XL U835 ( .A0(n459), .A1(n460), .B0(n458), .Y(mult_x_1_n312) );
  OAI21XL U836 ( .A0(n1023), .A1(n1019), .B0(n1020), .Y(mult_x_1_n317) );
  INVXL U837 ( .A(n461), .Y(n1055) );
  AOI21XL U838 ( .A0(n1055), .A1(n1053), .B0(n462), .Y(n466) );
  XOR2X1 U839 ( .A(n466), .B(n465), .Y(n1211) );
  CMPR32X1 U840 ( .A(n469), .B(n468), .C(n467), .CO(n998), .S(mult_x_1_n404)
         );
  XNOR2XL U841 ( .A(B[22]), .B(A[15]), .Y(n474) );
  CMPR32X1 U842 ( .A(n472), .B(n475), .C(n471), .CO(n467), .S(n477) );
  OAI22XL U843 ( .A0(n482), .A1(n99), .B0(n473), .B1(n884), .Y(n481) );
  XNOR2XL U844 ( .A(B[21]), .B(A[15]), .Y(n483) );
  OAI22XL U845 ( .A0(n483), .A1(n102), .B0(n474), .B1(n529), .Y(n480) );
  CMPR32X1 U846 ( .A(n481), .B(n480), .C(n479), .CO(n476), .S(mult_x_1_n414)
         );
  XNOR2X1 U847 ( .A(B[22]), .B(n856), .Y(n1046) );
  OAI22XL U848 ( .A0(n502), .A1(n485), .B0(n487), .B1(n486), .Y(n1048) );
  CMPR32X1 U849 ( .A(n492), .B(n491), .C(n490), .CO(mult_x_1_n419), .S(
        mult_x_1_n420) );
  CMPR32X1 U850 ( .A(n494), .B(n493), .C(n1048), .CO(mult_x_1_n421), .S(n490)
         );
  INVXL U851 ( .A(n500), .Y(n496) );
  OAI22XL U852 ( .A0(n502), .A1(n486), .B0(n524), .B1(n485), .Y(n507) );
  XNOR2XL U853 ( .A(B[20]), .B(n856), .Y(n509) );
  XNOR2X1 U854 ( .A(B[21]), .B(n856), .Y(n1047) );
  OAI22XL U855 ( .A0(n509), .A1(n99), .B0(n1047), .B1(n884), .Y(n513) );
  XNOR2XL U856 ( .A(B[22]), .B(n858), .Y(n525) );
  CMPR32X1 U857 ( .A(n506), .B(n505), .C(n504), .CO(mult_x_1_n425), .S(
        mult_x_1_n426) );
  CMPR32X1 U858 ( .A(n508), .B(n511), .C(n507), .CO(n505), .S(n517) );
  XNOR2X1 U859 ( .A(B[19]), .B(n856), .Y(n520) );
  OAI22XL U860 ( .A0(n520), .A1(n99), .B0(n509), .B1(n884), .Y(n523) );
  XNOR2XL U861 ( .A(B[17]), .B(A[15]), .Y(n531) );
  INVXL U862 ( .A(n511), .Y(n521) );
  CMPR32X1 U863 ( .A(n514), .B(n513), .C(n512), .CO(n504), .S(n515) );
  CMPR32X1 U864 ( .A(n517), .B(n516), .C(n515), .CO(mult_x_1_n433), .S(
        mult_x_1_n434) );
  XNOR2XL U865 ( .A(B[20]), .B(n858), .Y(n549) );
  XNOR2XL U866 ( .A(B[21]), .B(n858), .Y(n526) );
  OAI22XL U867 ( .A0(n549), .A1(n258), .B0(n526), .B1(n257), .Y(n542) );
  XNOR2X1 U868 ( .A(B[18]), .B(n856), .Y(n548) );
  OAI22XL U869 ( .A0(n548), .A1(n99), .B0(n520), .B1(n884), .Y(n540) );
  OAI22XL U870 ( .A0(n543), .A1(n485), .B0(n524), .B1(n486), .Y(n537) );
  OAI22XL U871 ( .A0(n526), .A1(n258), .B0(n525), .B1(n257), .Y(n536) );
  INVXL U872 ( .A(n538), .Y(n527) );
  OAI2BB1X1 U873 ( .A0N(n528), .A1N(n7), .B0(n527), .Y(n546) );
  XNOR2X1 U874 ( .A(B[16]), .B(A[15]), .Y(n530) );
  OAI22X2 U875 ( .A0(n530), .A1(n529), .B0(n562), .B1(n102), .Y(n547) );
  OAI22XL U876 ( .A0(n531), .A1(n529), .B0(n530), .B1(n102), .Y(n545) );
  CMPR32X1 U877 ( .A(n534), .B(n533), .C(n532), .CO(mult_x_1_n441), .S(
        mult_x_1_n442) );
  OAI22XL U878 ( .A0(n567), .A1(n7), .B0(n538), .B1(n528), .Y(n558) );
  OAI22X1 U879 ( .A0(n559), .A1(n485), .B0(n544), .B1(n486), .Y(n557) );
  OAI22XL U880 ( .A0(n568), .A1(n8), .B0(n539), .B1(n499), .Y(n556) );
  CMPR32X1 U881 ( .A(n542), .B(n541), .C(n540), .CO(n534), .S(n551) );
  OAI22XL U882 ( .A0(n544), .A1(n485), .B0(n543), .B1(n486), .Y(n555) );
  OAI22XL U883 ( .A0(n566), .A1(n99), .B0(n548), .B1(n884), .Y(n582) );
  XNOR2XL U884 ( .A(B[19]), .B(A[11]), .Y(n560) );
  OAI22XL U885 ( .A0(n560), .A1(n258), .B0(n549), .B1(n257), .Y(n581) );
  CMPR32X1 U886 ( .A(n555), .B(n554), .C(n553), .CO(mult_x_1_n453), .S(n550)
         );
  XNOR2XL U887 ( .A(B[20]), .B(A[9]), .Y(n588) );
  OAI22XL U888 ( .A0(n588), .A1(n485), .B0(n559), .B1(n486), .Y(n594) );
  INVXL U889 ( .A(n564), .Y(n561) );
  XNOR2X1 U890 ( .A(B[16]), .B(n856), .Y(n565) );
  INVXL U891 ( .A(n577), .Y(n626) );
  XNOR2XL U892 ( .A(B[25]), .B(A[3]), .Y(n618) );
  OAI22XL U893 ( .A0(n618), .A1(n329), .B0(n564), .B1(n617), .Y(n625) );
  XNOR2XL U894 ( .A(B[23]), .B(n9), .Y(n601) );
  OAI22XL U895 ( .A0(n613), .A1(n572), .B0(n571), .B1(n529), .Y(n603) );
  CMPR32X1 U896 ( .A(n583), .B(n582), .C(n581), .CO(n553), .S(n584) );
  XNOR2XL U897 ( .A(B[19]), .B(A[9]), .Y(n591) );
  OAI22XL U898 ( .A0(n591), .A1(n485), .B0(n588), .B1(n486), .Y(n608) );
  XNOR2XL U899 ( .A(B[18]), .B(A[9]), .Y(n606) );
  OAI22XL U900 ( .A0(n606), .A1(n485), .B0(n591), .B1(n486), .Y(n610) );
  ADDFHX4 U901 ( .A(n40), .B(n593), .CI(n592), .CO(n575), .S(n599) );
  CMPR32X1 U902 ( .A(n597), .B(n596), .C(n595), .CO(n574), .S(n598) );
  XNOR2XL U903 ( .A(B[22]), .B(A[5]), .Y(n637) );
  OAI22XL U904 ( .A0(n637), .A1(n7), .B0(n601), .B1(n528), .Y(n644) );
  XNOR2X1 U905 ( .A(n603), .B(n602), .Y(n643) );
  OAI22XL U906 ( .A0(n639), .A1(n99), .B0(n604), .B1(n884), .Y(n647) );
  OAI22XL U907 ( .A0(n640), .A1(n485), .B0(n606), .B1(n486), .Y(n645) );
  CMPR32X1 U908 ( .A(n609), .B(n608), .C(n607), .CO(n600), .S(n623) );
  CMPR32X1 U909 ( .A(n612), .B(n611), .C(n610), .CO(n607), .S(n661) );
  XNOR2XL U910 ( .A(B[23]), .B(A[3]), .Y(n662) );
  OAI22X1 U911 ( .A0(n651), .A1(n102), .B0(n615), .B1(n529), .Y(n650) );
  OAI22X1 U912 ( .A0(n638), .A1(n8), .B0(n619), .B1(n499), .Y(n629) );
  CMPR32X1 U913 ( .A(n624), .B(n623), .C(n622), .CO(mult_x_1_n485), .S(
        mult_x_1_n486) );
  CMPR32X1 U914 ( .A(n627), .B(n626), .C(n625), .CO(n597), .S(n636) );
  XNOR2XL U915 ( .A(B[19]), .B(A[7]), .Y(n641) );
  XNOR2XL U916 ( .A(B[12]), .B(n856), .Y(n666) );
  XNOR2XL U917 ( .A(B[18]), .B(A[7]), .Y(n667) );
  OAI22XL U918 ( .A0(n667), .A1(n8), .B0(n641), .B1(n499), .Y(n671) );
  CMPR32X1 U919 ( .A(n644), .B(n643), .C(n642), .CO(n624), .S(n657) );
  CMPR22X1 U920 ( .A(n650), .B(n649), .CO(n653), .S(n680) );
  CMPR32X1 U921 ( .A(n655), .B(n654), .C(n653), .CO(n660), .S(n685) );
  OAI22XL U922 ( .A0(n698), .A1(n329), .B0(n662), .B1(n617), .Y(n706) );
  XNOR2X1 U923 ( .A(B[20]), .B(A[5]), .Y(n699) );
  OAI22XL U924 ( .A0(n701), .A1(n665), .B0(n664), .B1(n257), .Y(n690) );
  XNOR2XL U925 ( .A(B[17]), .B(A[7]), .Y(n703) );
  OAI22XL U926 ( .A0(n703), .A1(n8), .B0(n667), .B1(n499), .Y(n688) );
  OAI22XL U927 ( .A0(n693), .A1(n369), .B0(n678), .B1(n892), .Y(n695) );
  CMPR32X1 U928 ( .A(n690), .B(n689), .C(n688), .CO(n704), .S(n709) );
  OAI22X1 U929 ( .A0(n730), .A1(n369), .B0(n693), .B1(n892), .Y(n732) );
  XNOR2XL U930 ( .A(B[7]), .B(A[15]), .Y(n727) );
  OAI22XL U931 ( .A0(n694), .A1(n529), .B0(n727), .B1(n102), .Y(n738) );
  XNOR2XL U932 ( .A(B[11]), .B(n858), .Y(n747) );
  XNOR2XL U933 ( .A(B[12]), .B(n858), .Y(n702) );
  OAI22XL U934 ( .A0(n716), .A1(n329), .B0(n698), .B1(n617), .Y(n723) );
  OAI22X1 U935 ( .A0(n718), .A1(n485), .B0(n700), .B1(n486), .Y(n726) );
  XNOR2XL U936 ( .A(B[16]), .B(A[7]), .Y(n720) );
  OAI22XL U937 ( .A0(n703), .A1(n499), .B0(n720), .B1(n8), .Y(n724) );
  CMPR32X1 U938 ( .A(n706), .B(n705), .C(n704), .CO(n684), .S(n711) );
  CMPR32X1 U939 ( .A(n712), .B(n711), .C(n710), .CO(mult_x_1_n527), .S(
        mult_x_1_n528) );
  XNOR2XL U940 ( .A(B[18]), .B(n9), .Y(n739) );
  XNOR2XL U941 ( .A(B[9]), .B(n856), .Y(n728) );
  OAI22XL U942 ( .A0(n720), .A1(n499), .B0(n740), .B1(n8), .Y(n751) );
  CMPR32X1 U943 ( .A(n723), .B(n722), .C(n721), .CO(n712), .S(n735) );
  CMPR32X1 U944 ( .A(n726), .B(n725), .C(n724), .CO(n721), .S(n762) );
  OAI22XL U945 ( .A0(n727), .A1(n529), .B0(n741), .B1(n102), .Y(n750) );
  OAI22XL U946 ( .A0(n728), .A1(n884), .B0(n766), .B1(n882), .Y(n749) );
  XNOR2XL U947 ( .A(B[19]), .B(A[3]), .Y(n764) );
  XNOR2XL U948 ( .A(B[21]), .B(A[1]), .Y(n763) );
  OAI22XL U949 ( .A0(n763), .A1(n369), .B0(n730), .B1(n892), .Y(n754) );
  CMPR32X1 U950 ( .A(n736), .B(n735), .C(n734), .CO(mult_x_1_n541), .S(
        mult_x_1_n542) );
  ADDHXL U951 ( .A(n738), .B(n737), .CO(n731), .S(n772) );
  XNOR2XL U952 ( .A(B[17]), .B(A[5]), .Y(n743) );
  XNOR2XL U953 ( .A(B[5]), .B(A[15]), .Y(n742) );
  XNOR2XL U954 ( .A(B[16]), .B(A[5]), .Y(n775) );
  OAI22XL U955 ( .A0(n743), .A1(n528), .B0(n775), .B1(n7), .Y(n776) );
  XNOR2XL U956 ( .A(B[10]), .B(n858), .Y(n774) );
  OAI22XL U957 ( .A0(n774), .A1(n258), .B0(n747), .B1(n257), .Y(n781) );
  XNOR2XL U958 ( .A(B[12]), .B(A[9]), .Y(n769) );
  OAI22XL U959 ( .A0(n769), .A1(n485), .B0(n748), .B1(n486), .Y(n780) );
  ADDHXL U960 ( .A(n750), .B(n749), .CO(n756), .S(n779) );
  CMPR32X1 U961 ( .A(n753), .B(n752), .C(n751), .CO(n744), .S(n786) );
  ADDFHX1 U962 ( .A(n756), .B(n755), .CI(n754), .CO(n761), .S(n785) );
  CMPR32X1 U963 ( .A(n759), .B(n758), .C(n757), .CO(mult_x_1_n555), .S(
        mult_x_1_n556) );
  XNOR2XL U964 ( .A(B[20]), .B(A[1]), .Y(n788) );
  OAI22XL U965 ( .A0(n788), .A1(n369), .B0(n763), .B1(n934), .Y(n797) );
  XNOR2XL U966 ( .A(B[18]), .B(A[3]), .Y(n789) );
  OAI22XL U967 ( .A0(n789), .A1(n329), .B0(n764), .B1(n328), .Y(n796) );
  OAI22XL U968 ( .A0(n802), .A1(n485), .B0(n769), .B1(n486), .Y(n798) );
  OAI22XL U969 ( .A0(n801), .A1(n8), .B0(n773), .B1(n499), .Y(n806) );
  OAI22XL U970 ( .A0(n794), .A1(n258), .B0(n774), .B1(n257), .Y(n805) );
  XNOR2XL U971 ( .A(B[15]), .B(A[5]), .Y(n813) );
  OAI22XL U972 ( .A0(n775), .A1(n528), .B0(n813), .B1(n7), .Y(n804) );
  CMPR32X1 U973 ( .A(n781), .B(n780), .C(n779), .CO(n787), .S(n810) );
  XNOR2XL U974 ( .A(B[19]), .B(A[1]), .Y(n822) );
  XNOR2XL U975 ( .A(B[17]), .B(A[3]), .Y(n803) );
  OAI22XL U976 ( .A0(n803), .A1(n329), .B0(n789), .B1(n617), .Y(n824) );
  XNOR2XL U977 ( .A(B[3]), .B(A[15]), .Y(n814) );
  OAI22X1 U978 ( .A0(n790), .A1(n529), .B0(n814), .B1(n102), .Y(n820) );
  XNOR2XL U979 ( .A(B[12]), .B(n895), .Y(n837) );
  OAI22X1 U980 ( .A0(n837), .A1(n8), .B0(n801), .B1(n499), .Y(n849) );
  XNOR2XL U981 ( .A(B[10]), .B(A[9]), .Y(n836) );
  XNOR2XL U982 ( .A(B[16]), .B(A[3]), .Y(n835) );
  OAI22XL U983 ( .A0(n803), .A1(n328), .B0(n835), .B1(n329), .Y(n847) );
  CMPR32X1 U984 ( .A(n806), .B(n805), .C(n804), .CO(n812), .S(n844) );
  XNOR2XL U985 ( .A(B[14]), .B(n9), .Y(n834) );
  OAI22XL U986 ( .A0(n834), .A1(n7), .B0(n813), .B1(n528), .Y(n852) );
  XNOR2XL U987 ( .A(B[2]), .B(A[15]), .Y(n818) );
  XNOR2XL U988 ( .A(n986), .B(A[15]), .Y(n816) );
  CMPR22X1 U989 ( .A(n820), .B(n819), .CO(n828), .S(n839) );
  CMPR32X1 U990 ( .A(n825), .B(n824), .C(n823), .CO(n809), .S(n842) );
  CMPR32X1 U991 ( .A(n828), .B(n826), .C(n827), .CO(n823), .S(n872) );
  XNOR2XL U992 ( .A(B[4]), .B(n856), .Y(n857) );
  OAI22XL U993 ( .A0(n829), .A1(n884), .B0(n857), .B1(n882), .Y(n862) );
  OAI22XL U994 ( .A0(n833), .A1(n832), .B0(n859), .B1(n258), .Y(n860) );
  XNOR2XL U995 ( .A(B[13]), .B(n9), .Y(n888) );
  OAI22XL U996 ( .A0(n888), .A1(n7), .B0(n834), .B1(n528), .Y(n865) );
  OAI22XL U997 ( .A0(n835), .A1(n328), .B0(n890), .B1(n329), .Y(n864) );
  XNOR2XL U998 ( .A(B[11]), .B(A[7]), .Y(n910) );
  OAI22XL U999 ( .A0(n910), .A1(n8), .B0(n837), .B1(n499), .Y(n908) );
  CMPR32X1 U1000 ( .A(n843), .B(n842), .C(n841), .CO(mult_x_1_n597), .S(
        mult_x_1_n598) );
  CMPR32X1 U1001 ( .A(n846), .B(n845), .C(n844), .CO(n807), .S(mult_x_1_n600)
         );
  CMPR32X1 U1002 ( .A(n849), .B(n848), .C(n847), .CO(n845), .S(n869) );
  CMPR32X1 U1003 ( .A(n852), .B(n851), .C(n850), .CO(n843), .S(n868) );
  XNOR2XL U1004 ( .A(B[17]), .B(A[1]), .Y(n893) );
  OAI22X1 U1005 ( .A0(n893), .A1(n369), .B0(n853), .B1(n934), .Y(n875) );
  XNOR2XL U1006 ( .A(B[3]), .B(n856), .Y(n885) );
  OAI22X1 U1007 ( .A0(n857), .A1(n884), .B0(n885), .B1(n882), .Y(n900) );
  XNOR2XL U1008 ( .A(B[5]), .B(n858), .Y(n887) );
  OAI22XL U1009 ( .A0(n859), .A1(n257), .B0(n887), .B1(n258), .Y(n899) );
  CMPR32X1 U1010 ( .A(n866), .B(n865), .C(n864), .CO(n871), .S(n873) );
  ADDFHX1 U1011 ( .A(n872), .B(n871), .CI(n870), .CO(n841), .S(mult_x_1_n614)
         );
  XNOR2XL U1012 ( .A(B[16]), .B(A[1]), .Y(n891) );
  OAI22X2 U1013 ( .A0(n891), .A1(n892), .B0(n935), .B1(n369), .Y(n943) );
  OAI22XL U1014 ( .A0(n885), .A1(n884), .B0(n883), .B1(n882), .Y(n897) );
  OAI22XL U1015 ( .A0(n887), .A1(n257), .B0(n886), .B1(n258), .Y(n896) );
  XNOR2XL U1016 ( .A(B[14]), .B(A[3]), .Y(n894) );
  OAI22XL U1017 ( .A0(n893), .A1(n892), .B0(n891), .B1(n369), .Y(n904) );
  XNOR2XL U1018 ( .A(B[13]), .B(A[3]), .Y(n937) );
  CMPR32X1 U1019 ( .A(n898), .B(n897), .C(n896), .CO(n914), .S(n939) );
  CMPR32X1 U1020 ( .A(n909), .B(n908), .C(n907), .CO(n870), .S(n922) );
  OAI22X1 U1021 ( .A0(n911), .A1(n8), .B0(n910), .B1(n499), .Y(n926) );
  OAI22X1 U1022 ( .A0(n931), .A1(n499), .B0(n930), .B1(n8), .Y(n961) );
  OAI22X1 U1023 ( .A0(n933), .A1(n7), .B0(n932), .B1(n528), .Y(n960) );
  OAI22XL U1024 ( .A0(n938), .A1(n329), .B0(n937), .B1(n328), .Y(n973) );
  CMPR32X1 U1025 ( .A(n941), .B(n940), .C(n939), .CO(n942), .S(n972) );
  CMPR32X1 U1026 ( .A(n953), .B(n952), .C(n951), .CO(n945), .S(n971) );
  OR2X2 U1027 ( .A(n957), .B(n956), .Y(n954) );
  NAND2XL U1028 ( .A(n957), .B(n956), .Y(n958) );
  CMPR32X1 U1029 ( .A(n965), .B(n964), .C(n963), .CO(n977), .S(n985) );
  CMPR32X1 U1030 ( .A(n985), .B(n984), .C(n983), .CO(mult_x_1_n679), .S(n316)
         );
  NOR2XL U1031 ( .A(n988), .B(n987), .Y(n989) );
  INVXL U1032 ( .A(n989), .Y(mult_x_1_n387) );
  CMPR32X1 U1033 ( .A(n992), .B(n991), .C(n990), .CO(n987), .S(n1028) );
  CMPR32X1 U1034 ( .A(n995), .B(n994), .C(n993), .CO(n1027), .S(n457) );
  INVXL U1035 ( .A(n996), .Y(mult_x_1_n388) );
  NOR2XL U1036 ( .A(n998), .B(n997), .Y(n999) );
  INVXL U1037 ( .A(n999), .Y(mult_x_1_n361) );
  CMPR32X1 U1038 ( .A(n1148), .B(n1145), .C(n1146), .CO(n1001), .S(n145) );
  OR2X2 U1039 ( .A(n1001), .B(n1000), .Y(n1030) );
  AND2X2 U1040 ( .A(n1030), .B(n1003), .Y(n1002) );
  NAND2XL U1041 ( .A(n12), .B(n1030), .Y(n1006) );
  INVXL U1042 ( .A(n1037), .Y(n1004) );
  AOI21XL U1043 ( .A0(n1030), .A1(n1004), .B0(n1034), .Y(n1005) );
  CMPR32X1 U1044 ( .A(n1143), .B(n1141), .C(n1144), .CO(n1008), .S(n1000) );
  OR2X2 U1045 ( .A(n1008), .B(n1007), .Y(n1035) );
  INVXL U1046 ( .A(n1015), .Y(n1017) );
  INVXL U1047 ( .A(n1019), .Y(n1021) );
  NAND2XL U1048 ( .A(n1021), .B(n1020), .Y(n1022) );
  CMPR32X1 U1049 ( .A(n1142), .B(n1138), .C(n1140), .CO(n1041), .S(n1007) );
  OR2X2 U1050 ( .A(n1041), .B(n1040), .Y(n1103) );
  CMPR32X1 U1051 ( .A(n1051), .B(n1050), .C(n1049), .CO(mult_x_1_n427), .S(
        mult_x_1_n428) );
  XNOR2X1 U1052 ( .A(n1055), .B(n1054), .Y(n1212) );
  CMPR32X1 U1053 ( .A(n1139), .B(n1136), .C(n1137), .CO(n1057), .S(n1040) );
  OR2X2 U1054 ( .A(n1057), .B(n1135), .Y(n1108) );
  NAND2XL U1055 ( .A(n1101), .B(n1060), .Y(n1062) );
  OAI21XL U1056 ( .A0(n1066), .A1(n1071), .B0(n1072), .Y(n1059) );
  AOI21XL U1057 ( .A0(n1104), .A1(n1060), .B0(n1059), .Y(n1061) );
  OAI21XL U1058 ( .A0(n1029), .A1(n1062), .B0(n1061), .Y(n1064) );
  OAI21XL U1059 ( .A0(n1029), .A1(n1070), .B0(n1069), .Y(n1075) );
  NAND2XL U1060 ( .A(n1077), .B(n1076), .Y(n1079) );
  XNOR2XL U1061 ( .A(n1079), .B(n1078), .Y(n1213) );
  AOI21XL U1062 ( .A0(n1084), .A1(n1123), .B0(n1080), .Y(n1082) );
  INVXL U1063 ( .A(n1085), .Y(n1087) );
  XOR2XL U1064 ( .A(n1089), .B(n1088), .Y(n1214) );
  XNOR2XL U1065 ( .A(n1100), .B(n1099), .Y(n1217) );
  XOR2XL U1066 ( .A(n1115), .B(n1114), .Y(n1216) );
  NAND2XL U1067 ( .A(n1116), .B(n1127), .Y(n1117) );
  XNOR2XL U1068 ( .A(n1121), .B(n1120), .Y(n1215) );
endmodule


module FFT2048_DW02_mult_2_stage_J1_17 ( A, B, TC, CLK, PRODUCT );
  input [15:0] A;
  input [26:0] B;
  output [42:0] PRODUCT;
  input TC, CLK;
  wire   n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, mult_x_1_n335, mult_x_1_n327, mult_x_1_n320,
         mult_x_1_n317, mult_x_1_n316, mult_x_1_n313, mult_x_1_n312,
         mult_x_1_n306, mult_x_1_n305, mult_x_1_n303, mult_x_1_n302,
         mult_x_1_n300, mult_x_1_n299, mult_x_1_n297, mult_x_1_n292,
         mult_x_1_n291, mult_x_1_n289, mult_x_1_n288, mult_x_1_n278,
         mult_x_1_n277, mult_x_1_n271, mult_x_1_n270, mult_x_1_n260,
         mult_x_1_n259, mult_x_1_n253, mult_x_1_n252, mult_x_1_n242,
         mult_x_1_n241, mult_x_1_n233, mult_x_1_n232, mult_x_1_n224,
         mult_x_1_n223, mult_x_1_n221, mult_x_1_n220, mult_x_1_n210,
         mult_x_1_n209, mult_x_1_n203, mult_x_1_n202, mult_x_1_n192,
         mult_x_1_n191, mult_x_1_n185, mult_x_1_n184, mult_x_1_n174,
         mult_x_1_n173, mult_x_1_n163, mult_x_1_n162, mult_x_1_n150,
         mult_x_1_n149, mult_x_1_n135, mult_x_1_n134, mult_x_1_n126,
         mult_x_1_n125, mult_x_1_n115, mult_x_1_n114, mult_x_1_n106,
         mult_x_1_n105, mult_x_1_n81, mult_x_1_n80, mult_x_1_n78, mult_x_1_n54,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262;

  DFFHQXL mult_x_1_clk_r_REG22_S1 ( .D(mult_x_1_n220), .CK(CLK), .Q(n1226) );
  DFFHQXL mult_x_1_clk_r_REG40_S1 ( .D(mult_x_1_n173), .CK(CLK), .Q(n1216) );
  DFFHQXL mult_x_1_clk_r_REG24_S1 ( .D(mult_x_1_n209), .CK(CLK), .Q(n1224) );
  DFFHQXL mult_x_1_clk_r_REG42_S1 ( .D(mult_x_1_n162), .CK(CLK), .Q(n1214) );
  DFFHQX4 mult_x_1_clk_r_REG61_S1 ( .D(mult_x_1_n335), .CK(CLK), .Q(n1262) );
  DFFHQX4 mult_x_1_clk_r_REG54_S1 ( .D(mult_x_1_n317), .CK(CLK), .Q(n1259) );
  DFFHQX4 mult_x_1_clk_r_REG1_S1 ( .D(mult_x_1_n306), .CK(CLK), .Q(n1258) );
  DFFHQX4 mult_x_1_clk_r_REG55_S1 ( .D(mult_x_1_n316), .CK(CLK), .Q(n1255) );
  DFFHQX1 mult_x_1_clk_r_REG0_S1 ( .D(mult_x_1_n313), .CK(CLK), .Q(n1254) );
  DFFHQX4 mult_x_1_clk_r_REG3_S1 ( .D(mult_x_1_n305), .CK(CLK), .Q(n1251) );
  DFFHQX4 mult_x_1_clk_r_REG5_S1 ( .D(mult_x_1_n303), .CK(CLK), .Q(n1250) );
  DFFHQX4 mult_x_1_clk_r_REG7_S1 ( .D(mult_x_1_n297), .CK(CLK), .Q(n1246) );
  DFFHQX4 mult_x_1_clk_r_REG10_S1 ( .D(mult_x_1_n292), .CK(CLK), .Q(n1245) );
  DFFHQX4 mult_x_1_clk_r_REG32_S1 ( .D(mult_x_1_n288), .CK(CLK), .Q(n1242) );
  DFFHQX4 mult_x_1_clk_r_REG29_S1 ( .D(mult_x_1_n278), .CK(CLK), .Q(n1241) );
  DFFHQX4 mult_x_1_clk_r_REG30_S1 ( .D(mult_x_1_n277), .CK(CLK), .Q(n1240) );
  DFFHQX4 mult_x_1_clk_r_REG25_S1 ( .D(mult_x_1_n260), .CK(CLK), .Q(n1237) );
  DFFHQX4 mult_x_1_clk_r_REG26_S1 ( .D(mult_x_1_n259), .CK(CLK), .Q(n1236) );
  DFFHQX1 mult_x_1_clk_r_REG17_S1 ( .D(mult_x_1_n233), .CK(CLK), .Q(n1231) );
  DFFHQX4 mult_x_1_clk_r_REG18_S1 ( .D(mult_x_1_n232), .CK(CLK), .Q(n1230) );
  DFFHQXL clk_r_REG58_S1 ( .D(n1276), .CK(CLK), .Q(PRODUCT[12]) );
  DFFHQXL mult_x_1_clk_r_REG20_S1 ( .D(mult_x_1_n223), .CK(CLK), .Q(n1228) );
  DFFHQXL clk_r_REG60_S1 ( .D(n1277), .CK(CLK), .Q(PRODUCT[11]) );
  DFFHQXL mult_x_1_clk_r_REG37_S1 ( .D(mult_x_1_n185), .CK(CLK), .Q(n1219) );
  DFFHQX4 mult_x_1_clk_r_REG31_S1 ( .D(mult_x_1_n289), .CK(CLK), .Q(n1243) );
  DFFHQXL mult_x_1_clk_r_REG34_S1 ( .D(mult_x_1_n202), .CK(CLK), .Q(n1222) );
  DFFHQXL mult_x_1_clk_r_REG36_S1 ( .D(mult_x_1_n191), .CK(CLK), .Q(n1220) );
  DFFHQX1 mult_x_1_clk_r_REG56_S1 ( .D(mult_x_1_n81), .CK(CLK), .Q(n1257) );
  DFFHQXL clk_r_REG62_S1 ( .D(n1278), .CK(CLK), .Q(PRODUCT[10]) );
  DFFHQXL mult_x_1_clk_r_REG35_S1 ( .D(mult_x_1_n192), .CK(CLK), .Q(n1221) );
  DFFHQXL mult_x_1_clk_r_REG59_S1 ( .D(mult_x_1_n327), .CK(CLK), .Q(n1261) );
  DFFHQXL mult_x_1_clk_r_REG41_S1 ( .D(mult_x_1_n163), .CK(CLK), .Q(n1215) );
  DFFHQXL mult_x_1_clk_r_REG33_S1 ( .D(mult_x_1_n203), .CK(CLK), .Q(n1223) );
  DFFHQXL clk_r_REG63_S1 ( .D(n1279), .CK(CLK), .Q(PRODUCT[9]) );
  DFFHQXL mult_x_1_clk_r_REG4_S1 ( .D(mult_x_1_n78), .CK(CLK), .Q(n1252) );
  DFFHQXL mult_x_1_clk_r_REG23_S1 ( .D(mult_x_1_n210), .CK(CLK), .Q(n1225) );
  DFFHQXL clk_r_REG64_S1 ( .D(n1280), .CK(CLK), .Q(PRODUCT[8]) );
  DFFHQXL mult_x_1_clk_r_REG44_S1 ( .D(mult_x_1_n149), .CK(CLK), .Q(n1212) );
  DFFHQXL mult_x_1_clk_r_REG19_S1 ( .D(mult_x_1_n224), .CK(CLK), .Q(n1229) );
  DFFHQXL mult_x_1_clk_r_REG39_S1 ( .D(mult_x_1_n174), .CK(CLK), .Q(n1217) );
  DFFHQX1 mult_x_1_clk_r_REG11_S1 ( .D(mult_x_1_n291), .CK(CLK), .Q(n1244) );
  DFFHQXL clk_r_REG65_S1 ( .D(n1281), .CK(CLK), .Q(PRODUCT[7]) );
  DFFHQXL clk_r_REG66_S1 ( .D(n1282), .CK(CLK), .Q(PRODUCT[6]) );
  DFFHQXL clk_r_REG67_S1 ( .D(n1283), .CK(CLK), .Q(PRODUCT[5]) );
  DFFHQXL clk_r_REG68_S1 ( .D(n1284), .CK(CLK), .Q(PRODUCT[4]) );
  DFFHQXL clk_r_REG69_S1 ( .D(n1285), .CK(CLK), .Q(PRODUCT[3]) );
  DFFHQXL clk_r_REG70_S1 ( .D(n1286), .CK(CLK), .Q(PRODUCT[2]) );
  DFFHQXL clk_r_REG71_S1 ( .D(n1287), .CK(CLK), .Q(PRODUCT[1]) );
  DFFHQXL clk_r_REG72_S1 ( .D(n1288), .CK(CLK), .Q(PRODUCT[0]) );
  DFFHQXL mult_x_1_clk_r_REG6_S1 ( .D(mult_x_1_n302), .CK(CLK), .Q(n1249) );
  DFFHQX1 mult_x_1_clk_r_REG57_S1 ( .D(mult_x_1_n320), .CK(CLK), .Q(n1260) );
  DFFHQX1 mult_x_1_clk_r_REG53_S1 ( .D(mult_x_1_n80), .CK(CLK), .Q(n1256) );
  DFFHQXL mult_x_1_clk_r_REG21_S1 ( .D(mult_x_1_n221), .CK(CLK), .Q(n1227) );
  DFFHQXL mult_x_1_clk_r_REG38_S1 ( .D(mult_x_1_n184), .CK(CLK), .Q(n1218) );
  DFFHQXL mult_x_1_clk_r_REG43_S1 ( .D(mult_x_1_n150), .CK(CLK), .Q(n1213) );
  DFFHQXL mult_x_1_clk_r_REG45_S1 ( .D(mult_x_1_n135), .CK(CLK), .Q(n1211) );
  DFFHQXL mult_x_1_clk_r_REG46_S1 ( .D(mult_x_1_n134), .CK(CLK), .Q(n1210) );
  DFFHQXL mult_x_1_clk_r_REG47_S1 ( .D(mult_x_1_n126), .CK(CLK), .Q(n1209) );
  DFFHQXL mult_x_1_clk_r_REG48_S1 ( .D(mult_x_1_n125), .CK(CLK), .Q(n1208) );
  DFFHQXL mult_x_1_clk_r_REG49_S1 ( .D(mult_x_1_n115), .CK(CLK), .Q(n1207) );
  DFFHQXL mult_x_1_clk_r_REG50_S1 ( .D(mult_x_1_n114), .CK(CLK), .Q(n1206) );
  DFFHQXL mult_x_1_clk_r_REG51_S1 ( .D(mult_x_1_n106), .CK(CLK), .Q(n1205) );
  DFFHQXL mult_x_1_clk_r_REG52_S1 ( .D(mult_x_1_n105), .CK(CLK), .Q(n1204) );
  DFFHQXL mult_x_1_clk_r_REG12_S1 ( .D(mult_x_1_n54), .CK(CLK), .Q(n1203) );
  DFFHQX1 mult_x_1_clk_r_REG2_S1 ( .D(mult_x_1_n312), .CK(CLK), .Q(n1253) );
  DFFHQX2 mult_x_1_clk_r_REG16_S1 ( .D(mult_x_1_n241), .CK(CLK), .Q(n1232) );
  DFFHQX2 mult_x_1_clk_r_REG8_S1 ( .D(mult_x_1_n300), .CK(CLK), .Q(n1248) );
  DFFHQX1 mult_x_1_clk_r_REG15_S1 ( .D(mult_x_1_n242), .CK(CLK), .Q(n1233) );
  DFFHQX2 mult_x_1_clk_r_REG27_S1 ( .D(mult_x_1_n271), .CK(CLK), .Q(n1239) );
  DFFHQX2 mult_x_1_clk_r_REG28_S1 ( .D(mult_x_1_n270), .CK(CLK), .Q(n1238) );
  DFFHQX2 mult_x_1_clk_r_REG9_S1 ( .D(mult_x_1_n299), .CK(CLK), .Q(n1247) );
  DFFHQX2 mult_x_1_clk_r_REG14_S1 ( .D(mult_x_1_n252), .CK(CLK), .Q(n1234) );
  DFFHQX1 mult_x_1_clk_r_REG13_S1 ( .D(mult_x_1_n253), .CK(CLK), .Q(n1235) );
  CMPR32X1 U1 ( .A(n1056), .B(n1055), .C(n1054), .CO(n1072), .S(n404) );
  ADDFHX1 U2 ( .A(n548), .B(n547), .CI(n546), .CO(n537), .S(n574) );
  ADDFHX1 U3 ( .A(n747), .B(n746), .CI(n745), .CO(n720), .S(n754) );
  ADDFHX1 U4 ( .A(n572), .B(n571), .CI(n570), .CO(n547), .S(n576) );
  ADDFHX1 U5 ( .A(n946), .B(n945), .CI(n944), .CO(n926), .S(n951) );
  ADDFHX1 U6 ( .A(n949), .B(n948), .CI(n947), .CO(n950), .S(n954) );
  ADDFHX1 U7 ( .A(n940), .B(n939), .CI(n938), .CO(n945), .S(n947) );
  ADDFHX1 U8 ( .A(n696), .B(n695), .CI(n694), .CO(n709), .S(n746) );
  ADDFHX1 U9 ( .A(n937), .B(n936), .CI(n935), .CO(n948), .S(n941) );
  CMPR32X1 U10 ( .A(n770), .B(n769), .C(n768), .CO(n782), .S(n824) );
  INVXL U11 ( .A(n943), .Y(n46) );
  ADDFHX1 U12 ( .A(n992), .B(n991), .CI(n990), .CO(n1000), .S(n350) );
  XNOR2X1 U13 ( .A(B[17]), .B(n82), .Y(n766) );
  ADDFHX1 U14 ( .A(n337), .B(n336), .CI(n335), .CO(n342), .S(n344) );
  INVX1 U15 ( .A(n438), .Y(n437) );
  BUFX3 U16 ( .A(A[5]), .Y(n812) );
  BUFX3 U17 ( .A(A[1]), .Y(n484) );
  NAND2X1 U18 ( .A(n1045), .B(n17), .Y(n1198) );
  XNOR2X1 U19 ( .A(n1201), .B(n607), .Y(PRODUCT[27]) );
  XOR2X1 U20 ( .A(n7), .B(n753), .Y(PRODUCT[23]) );
  OAI21XL U21 ( .A0(n98), .A1(n789), .B0(n788), .Y(n792) );
  XOR2X1 U22 ( .A(n952), .B(n25), .Y(PRODUCT[17]) );
  OAI21XL U23 ( .A0(n1234), .A1(n1237), .B0(n1235), .Y(n641) );
  NOR2X2 U24 ( .A(n1234), .B(n1236), .Y(n638) );
  OAI21X2 U25 ( .A0(n1245), .A1(n1242), .B0(n1243), .Y(n112) );
  OAI22X1 U26 ( .A0(n1060), .A1(n173), .B0(n1061), .B1(n157), .Y(n172) );
  XNOR2XL U27 ( .A(n907), .B(n47), .Y(PRODUCT[19]) );
  XOR2X1 U28 ( .A(n472), .B(n61), .Y(PRODUCT[31]) );
  XNOR2XL U29 ( .A(n438), .B(n807), .Y(n233) );
  XNOR2XL U30 ( .A(n815), .B(n807), .Y(n326) );
  BUFX3 U31 ( .A(A[3]), .Y(n438) );
  XNOR2XL U32 ( .A(B[18]), .B(n82), .Y(n730) );
  XNOR2XL U33 ( .A(A[13]), .B(B[6]), .Y(n808) );
  XNOR2XL U34 ( .A(n6), .B(B[0]), .Y(n124) );
  XNOR2XL U35 ( .A(n1062), .B(B[3]), .Y(n136) );
  XNOR2XL U36 ( .A(n1129), .B(n812), .Y(n33) );
  XNOR2XL U37 ( .A(n1062), .B(n1129), .Y(n1082) );
  XNOR2XL U38 ( .A(A[10]), .B(A[9]), .Y(n1109) );
  XNOR2XL U39 ( .A(A[13]), .B(n1146), .Y(n1131) );
  ADDFX2 U40 ( .A(n706), .B(n705), .CI(n704), .CO(n724), .S(n757) );
  XOR2XL U41 ( .A(n32), .B(n419), .Y(n462) );
  XOR2XL U42 ( .A(n1160), .B(n1159), .Y(n1280) );
  AND2X4 U43 ( .A(n1258), .B(n1246), .Y(n5) );
  AOI21XL U44 ( .A0(n217), .A1(n540), .B0(n216), .Y(n218) );
  NOR2X1 U45 ( .A(n538), .B(n537), .Y(mult_x_1_n202) );
  INVX1 U46 ( .A(n1026), .Y(n1160) );
  INVX1 U47 ( .A(n993), .Y(n1015) );
  NOR2X1 U48 ( .A(n1006), .B(n1005), .Y(n1007) );
  NAND2X1 U49 ( .A(n1001), .B(n1000), .Y(n1013) );
  NAND2XL U50 ( .A(n31), .B(n30), .Y(n467) );
  XNOR2X1 U51 ( .A(n1170), .B(n1169), .Y(n1282) );
  INVX1 U52 ( .A(n349), .Y(n34) );
  NAND2X1 U53 ( .A(n350), .B(n349), .Y(n1019) );
  OAI21XL U54 ( .A0(n419), .A1(n420), .B0(n418), .Y(n31) );
  XOR2X1 U55 ( .A(n77), .B(n985), .Y(n987) );
  NAND2XL U56 ( .A(n42), .B(n172), .Y(n41) );
  CLKBUFX2 U57 ( .A(n918), .Y(n63) );
  XNOR2X1 U58 ( .A(n484), .B(n1146), .Y(n514) );
  XNOR2X1 U59 ( .A(n1202), .B(n1203), .Y(PRODUCT[40]) );
  XNOR2X1 U60 ( .A(n812), .B(B[13]), .Y(n852) );
  NAND2BXL U61 ( .AN(n1051), .B(n20), .Y(n19) );
  AOI21X1 U62 ( .A0(n1198), .A1(n1094), .B0(n1093), .Y(n1095) );
  INVXL U63 ( .A(n1201), .Y(n20) );
  AOI21X1 U64 ( .A0(n1198), .A1(n1089), .B0(n1092), .Y(n16) );
  XNOR2X1 U65 ( .A(n484), .B(B[3]), .Y(n278) );
  NAND2X1 U66 ( .A(n29), .B(n113), .Y(n116) );
  NAND2BXL U67 ( .AN(n640), .B(n47), .Y(n8) );
  INVXL U68 ( .A(n844), .Y(n36) );
  AND2X2 U69 ( .A(n352), .B(n1217), .Y(n60) );
  INVX1 U70 ( .A(n112), .Y(n113) );
  AND2X2 U71 ( .A(n575), .B(n1227), .Y(n58) );
  AOI2BB1X2 U72 ( .A0N(n1238), .A1N(n1241), .B0(n104), .Y(n14) );
  OAI21XL U73 ( .A0(n1230), .A1(n1233), .B0(n1231), .Y(n10) );
  INVXL U74 ( .A(n1211), .Y(n1092) );
  NOR2X1 U75 ( .A(n1224), .B(n1222), .Y(n217) );
  INVX1 U76 ( .A(n1251), .Y(n26) );
  XOR2X1 U77 ( .A(n92), .B(n1021), .Y(n1277) );
  XNOR2X1 U78 ( .A(n1031), .B(n1030), .Y(n1279) );
  OAI2BB1X1 U79 ( .A0N(n943), .A1N(n942), .B0(n83), .Y(n953) );
  NAND2X1 U80 ( .A(n1006), .B(n1005), .Y(n1008) );
  XOR2X1 U81 ( .A(n535), .B(n536), .Y(n40) );
  NOR2X1 U82 ( .A(n1001), .B(n1000), .Y(n993) );
  NAND2XL U83 ( .A(n637), .B(n636), .Y(mult_x_1_n224) );
  NAND2XL U84 ( .A(n85), .B(n1164), .Y(n298) );
  ADDFHX1 U85 ( .A(n999), .B(n998), .CI(n997), .CO(n1005), .S(n1003) );
  NOR2X1 U86 ( .A(n303), .B(n302), .Y(n1027) );
  NAND2XL U87 ( .A(n419), .B(n420), .Y(n30) );
  INVX1 U88 ( .A(n347), .Y(n73) );
  INVX1 U89 ( .A(n457), .Y(n491) );
  XOR2X1 U90 ( .A(n418), .B(n420), .Y(n32) );
  NAND2X1 U91 ( .A(n301), .B(n300), .Y(n1157) );
  INVX1 U92 ( .A(n44), .Y(n42) );
  NOR2X1 U93 ( .A(n301), .B(n300), .Y(n1156) );
  OAI22X1 U94 ( .A0(n33), .A1(n853), .B0(n855), .B1(n452), .Y(n461) );
  NAND2BXL U95 ( .AN(n519), .B(n103), .Y(n102) );
  NAND2X1 U96 ( .A(n19), .B(n16), .Y(n1053) );
  BUFX3 U97 ( .A(B[5]), .Y(n807) );
  NAND2X1 U98 ( .A(n751), .B(n8), .Y(n7) );
  INVXL U99 ( .A(n1046), .Y(n18) );
  INVXL U100 ( .A(n713), .Y(n751) );
  NAND2X2 U101 ( .A(n15), .B(n14), .Y(n713) );
  INVX1 U102 ( .A(n214), .Y(n12) );
  INVXL U103 ( .A(n67), .Y(n66) );
  NAND2X1 U104 ( .A(n433), .B(n1219), .Y(n434) );
  AND2X2 U105 ( .A(n471), .B(n1221), .Y(n61) );
  NAND2X1 U106 ( .A(n505), .B(n1223), .Y(n506) );
  NAND2X1 U107 ( .A(n873), .B(n1243), .Y(n874) );
  AOI21X1 U108 ( .A0(n641), .A1(n13), .B0(n10), .Y(n9) );
  NAND2X1 U109 ( .A(n638), .B(n13), .Y(n214) );
  NAND2X1 U110 ( .A(n217), .B(n539), .Y(n1035) );
  INVX1 U111 ( .A(n1208), .Y(n1091) );
  INVX1 U112 ( .A(n1212), .Y(n1039) );
  INVX1 U113 ( .A(n1214), .Y(n1033) );
  NAND2X1 U114 ( .A(n1251), .B(n1246), .Y(n28) );
  INVX4 U115 ( .A(n369), .Y(n6) );
  BUFX3 U116 ( .A(A[13]), .Y(n1100) );
  NOR2X1 U117 ( .A(n954), .B(n953), .Y(mult_x_1_n302) );
  NAND2XL U118 ( .A(n537), .B(n538), .Y(mult_x_1_n203) );
  NAND3X1 U119 ( .A(n1025), .B(n1020), .C(n1023), .Y(n69) );
  ADDFHX2 U120 ( .A(n510), .B(n509), .CI(n508), .CO(n500), .S(n538) );
  XNOR2X1 U121 ( .A(n1025), .B(n1024), .Y(n1278) );
  NAND2XL U122 ( .A(n872), .B(n871), .Y(mult_x_1_n278) );
  INVXL U123 ( .A(n474), .Y(n100) );
  XOR2X1 U124 ( .A(n534), .B(n40), .Y(n546) );
  OAI2BB1X1 U125 ( .A0N(n304), .A1N(n1026), .B0(n70), .Y(n1025) );
  OR2X2 U126 ( .A(n535), .B(n536), .Y(n39) );
  INVXL U127 ( .A(n1018), .Y(n1022) );
  ADDFHX2 U128 ( .A(n194), .B(n193), .CI(n192), .CO(n942), .S(n208) );
  ADDFHX1 U129 ( .A(n467), .B(n466), .CI(n465), .CO(n428), .S(n468) );
  INVXL U130 ( .A(n475), .Y(n101) );
  INVXL U131 ( .A(n829), .Y(n95) );
  INVXL U132 ( .A(n877), .Y(n106) );
  INVXL U133 ( .A(n1028), .Y(n71) );
  ADDFHX1 U134 ( .A(n610), .B(n609), .CI(n608), .CO(n604), .S(n637) );
  OAI2BB1X1 U135 ( .A0N(n171), .A1N(n43), .B0(n41), .Y(n166) );
  NAND2BXL U136 ( .AN(n1162), .B(n1163), .Y(n85) );
  ADDFHX2 U137 ( .A(n603), .B(n602), .CI(n601), .CO(n577), .S(n608) );
  ADDFX2 U138 ( .A(n524), .B(n523), .CI(n522), .CO(n536), .S(n571) );
  NAND2XL U139 ( .A(n80), .B(n79), .Y(n923) );
  ADDFHX2 U140 ( .A(n673), .B(n672), .CI(n671), .CO(n646), .S(n681) );
  OR2XL U141 ( .A(n1153), .B(n1152), .Y(n1155) );
  INVXL U142 ( .A(n878), .Y(n107) );
  INVXL U143 ( .A(n830), .Y(n96) );
  ADDFHX2 U144 ( .A(n782), .B(n781), .CI(n780), .CO(n755), .S(n793) );
  NAND2BXL U145 ( .AN(n810), .B(n55), .Y(n54) );
  XOR2X1 U146 ( .A(n809), .B(n56), .Y(n869) );
  NAND2XL U147 ( .A(n933), .B(n934), .Y(n79) );
  INVXL U148 ( .A(n933), .Y(n81) );
  NAND2XL U149 ( .A(n985), .B(n986), .Y(n75) );
  NAND2XL U150 ( .A(n111), .B(n981), .Y(n110) );
  XNOR3X2 U151 ( .A(n172), .B(n44), .C(n171), .Y(n976) );
  INVXL U152 ( .A(n296), .Y(n86) );
  INVXL U153 ( .A(n986), .Y(n78) );
  OAI21X1 U154 ( .A0(n37), .A1(n846), .B0(n35), .Y(n457) );
  ADDFHX1 U155 ( .A(n776), .B(n775), .CI(n774), .CO(n768), .S(n832) );
  NAND2XL U156 ( .A(n810), .B(n811), .Y(n53) );
  ADDFHX2 U157 ( .A(n735), .B(n734), .CI(n733), .CO(n747), .S(n781) );
  OAI22X1 U158 ( .A0(n33), .A1(n855), .B0(n372), .B1(n853), .Y(n416) );
  OAI21XL U159 ( .A0(n37), .A1(n520), .B0(n102), .Y(n533) );
  NAND2BX1 U160 ( .AN(n439), .B(n36), .Y(n35) );
  OAI22X1 U161 ( .A0(n1060), .A1(n411), .B0(n1061), .B1(n406), .Y(n420) );
  XNOR2X1 U162 ( .A(n1142), .B(n1141), .Y(PRODUCT[39]) );
  XNOR2X1 U163 ( .A(n1099), .B(n1098), .Y(PRODUCT[38]) );
  OR2X2 U164 ( .A(n275), .B(n274), .Y(n273) );
  XNOR2X1 U165 ( .A(n361), .B(n360), .Y(PRODUCT[35]) );
  AND2XL U166 ( .A(n1186), .B(n1185), .Y(n1287) );
  OR2XL U167 ( .A(n1184), .B(n1183), .Y(n1186) );
  NAND2BX1 U168 ( .AN(n218), .B(n18), .Y(n17) );
  NAND2BX1 U169 ( .AN(n114), .B(n47), .Y(n29) );
  INVXL U170 ( .A(n846), .Y(n103) );
  NAND2X2 U171 ( .A(n11), .B(n9), .Y(n23) );
  AND2XL U172 ( .A(n1191), .B(n1193), .Y(n1197) );
  NAND2X1 U173 ( .A(n713), .B(n12), .Y(n11) );
  INVX1 U174 ( .A(n640), .Y(n750) );
  NAND2BXL U175 ( .AN(n676), .B(n639), .Y(n52) );
  NAND2X1 U176 ( .A(n119), .B(n1109), .Y(n1108) );
  NAND2X1 U177 ( .A(n125), .B(n126), .Y(n1133) );
  NAND2X1 U178 ( .A(n127), .B(n128), .Y(n306) );
  NAND2X1 U179 ( .A(n112), .B(n213), .Y(n15) );
  AND2X2 U180 ( .A(n752), .B(n1237), .Y(n753) );
  XOR2X1 U181 ( .A(A[2]), .B(n438), .Y(n120) );
  NAND2X1 U182 ( .A(n117), .B(n118), .Y(n656) );
  AND2X2 U183 ( .A(n606), .B(n1229), .Y(n607) );
  INVXL U184 ( .A(n1247), .Y(n929) );
  INVXL U185 ( .A(n1233), .Y(n50) );
  INVX1 U186 ( .A(n1240), .Y(n787) );
  XNOR2X1 U187 ( .A(A[8]), .B(A[7]), .Y(n118) );
  INVX1 U188 ( .A(n1210), .Y(n1089) );
  INVX1 U189 ( .A(A[0]), .Y(n131) );
  OAI21X4 U190 ( .A0(n928), .A1(n28), .B0(n27), .Y(n47) );
  NOR2X1 U191 ( .A(n1230), .B(n1232), .Y(n13) );
  NOR2X1 U192 ( .A(n1238), .B(n1240), .Y(n213) );
  NOR2X4 U193 ( .A(n21), .B(n5), .Y(n27) );
  OAI21X4 U194 ( .A0(n1247), .A1(n1250), .B0(n1248), .Y(n21) );
  XOR2X2 U195 ( .A(n22), .B(n58), .Y(PRODUCT[28]) );
  OAI21X1 U196 ( .A0(n1201), .A1(n1228), .B0(n1229), .Y(n22) );
  NOR2X4 U197 ( .A(n24), .B(n23), .Y(n1201) );
  NOR2BX4 U198 ( .AN(n215), .B(n98), .Y(n24) );
  NAND2BX1 U199 ( .AN(n1249), .B(n1250), .Y(n25) );
  AOI2BB1X4 U200 ( .A0N(n928), .A1N(n26), .B0(n1258), .Y(n952) );
  AOI21X4 U201 ( .A0(n1255), .A1(n1262), .B0(n1259), .Y(n928) );
  CLKINVX3 U202 ( .A(n47), .Y(n98) );
  AOI21X1 U203 ( .A0(n470), .A1(n1034), .B0(n1044), .Y(n219) );
  OAI22X1 U204 ( .A0(n846), .A1(n806), .B0(n844), .B1(n766), .Y(n818) );
  NAND2BX1 U205 ( .AN(n350), .B(n34), .Y(n1020) );
  XOR2X1 U206 ( .A(n1129), .B(n437), .Y(n37) );
  OAI2BB1X2 U207 ( .A0N(n39), .A1N(n534), .B0(n38), .Y(n509) );
  NAND2X1 U208 ( .A(n535), .B(n536), .Y(n38) );
  NAND2BX1 U209 ( .AN(n172), .B(n44), .Y(n43) );
  AOI2BB1X1 U210 ( .A0N(n158), .A1N(n844), .B0(n45), .Y(n44) );
  NOR2X1 U211 ( .A(n159), .B(n846), .Y(n45) );
  XOR2X1 U212 ( .A(n942), .B(n46), .Y(n84) );
  NAND2X1 U213 ( .A(n785), .B(n213), .Y(n640) );
  NAND3X1 U214 ( .A(n52), .B(n49), .C(n48), .Y(n644) );
  NAND3XL U215 ( .A(n47), .B(n750), .C(n51), .Y(n48) );
  AOI21X1 U216 ( .A0(n713), .A1(n51), .B0(n50), .Y(n49) );
  NOR2BX1 U217 ( .AN(n638), .B(n1232), .Y(n51) );
  OAI2BB1X1 U218 ( .A0N(n54), .A1N(n809), .B0(n53), .Y(n825) );
  INVXL U219 ( .A(n811), .Y(n55) );
  XOR2X1 U220 ( .A(n810), .B(n811), .Y(n56) );
  XNOR2X1 U221 ( .A(B[17]), .B(n803), .Y(n555) );
  XNOR2X1 U222 ( .A(B[17]), .B(n812), .Y(n697) );
  XNOR2X1 U223 ( .A(B[17]), .B(n484), .Y(n836) );
  XNOR2X1 U224 ( .A(B[17]), .B(n1062), .Y(n489) );
  XNOR2X1 U225 ( .A(B[17]), .B(n815), .Y(n626) );
  XNOR2X1 U226 ( .A(B[17]), .B(n1100), .Y(n447) );
  XNOR2X1 U227 ( .A(B[17]), .B(n6), .Y(n370) );
  OAI22X1 U228 ( .A0(n1060), .A1(n765), .B0(n1061), .B1(n729), .Y(n776) );
  OAI22X1 U229 ( .A0(n846), .A1(n145), .B0(n844), .B1(n187), .Y(n185) );
  OAI21XL U230 ( .A0(n958), .A1(mult_x_1_n313), .B0(n959), .Y(mult_x_1_n306)
         );
  NOR2X1 U231 ( .A(n212), .B(n211), .Y(n958) );
  NAND2X1 U232 ( .A(n956), .B(n957), .Y(mult_x_1_n313) );
  OAI22X1 U233 ( .A0(n801), .A1(n174), .B0(n142), .B1(n1032), .Y(n178) );
  XNOR2X2 U234 ( .A(n484), .B(B[12]), .Y(n142) );
  OAI22X1 U235 ( .A0(n846), .A1(n619), .B0(n844), .B1(n587), .Y(n628) );
  XNOR2X1 U236 ( .A(B[22]), .B(n82), .Y(n587) );
  OAI22X1 U237 ( .A0(n861), .A1(n448), .B0(n859), .B1(n408), .Y(n445) );
  ADDFX2 U238 ( .A(n916), .B(n915), .CI(n914), .CO(n940), .S(n936) );
  OAI22X1 U239 ( .A0(n656), .A1(n121), .B0(n1061), .B1(n186), .Y(n200) );
  XNOR2X1 U240 ( .A(n803), .B(B[18]), .Y(n518) );
  XNOR2X1 U241 ( .A(n84), .B(n941), .Y(n212) );
  NAND2XL U242 ( .A(n1091), .B(n1209), .Y(n1052) );
  NAND2XL U243 ( .A(n1036), .B(n1089), .Y(n1051) );
  NAND2XL U244 ( .A(n1039), .B(n1213), .Y(n360) );
  XNOR2XL U245 ( .A(n815), .B(B[6]), .Y(n144) );
  NAND2XL U246 ( .A(n1034), .B(n1043), .Y(n1046) );
  NAND2XL U247 ( .A(n1097), .B(n1207), .Y(n1098) );
  INVXL U248 ( .A(n1206), .Y(n1097) );
  AOI21XL U249 ( .A0(n713), .A1(n752), .B0(n712), .Y(n714) );
  INVXL U250 ( .A(n1237), .Y(n712) );
  XNOR2X1 U251 ( .A(B[11]), .B(n484), .Y(n174) );
  XNOR2XL U252 ( .A(n812), .B(B[8]), .Y(n161) );
  XNOR2XL U253 ( .A(n815), .B(B[4]), .Y(n327) );
  XNOR2XL U254 ( .A(n438), .B(B[8]), .Y(n331) );
  XNOR2XL U255 ( .A(n815), .B(n1146), .Y(n377) );
  XNOR2X1 U256 ( .A(n803), .B(n1129), .Y(n393) );
  XNOR2XL U257 ( .A(n6), .B(B[16]), .Y(n409) );
  XNOR2XL U258 ( .A(n803), .B(B[24]), .Y(n381) );
  XNOR2XL U259 ( .A(n1100), .B(B[20]), .Y(n379) );
  CLKINVX3 U260 ( .A(n437), .Y(n82) );
  NOR2XL U261 ( .A(n1137), .B(n1206), .Y(n1191) );
  INVXL U262 ( .A(n1204), .Y(n1193) );
  OR2X2 U263 ( .A(n982), .B(n983), .Y(n111) );
  XNOR2XL U264 ( .A(n6), .B(B[21]), .Y(n1080) );
  OAI22XL U265 ( .A0(n1060), .A1(n307), .B0(n1061), .B1(n173), .Y(n980) );
  XNOR2XL U266 ( .A(n1100), .B(B[22]), .Y(n1064) );
  XNOR2XL U267 ( .A(n6), .B(B[19]), .Y(n392) );
  XNOR2XL U268 ( .A(n1100), .B(B[21]), .Y(n391) );
  XNOR2XL U269 ( .A(n1062), .B(B[24]), .Y(n1063) );
  XNOR2XL U270 ( .A(n6), .B(B[18]), .Y(n376) );
  XNOR2XL U271 ( .A(n1062), .B(B[22]), .Y(n380) );
  XNOR2XL U272 ( .A(n815), .B(B[9]), .Y(n191) );
  ADDFX2 U273 ( .A(n919), .B(n63), .CI(n917), .CO(n925), .S(n939) );
  ADDFX2 U274 ( .A(n242), .B(n241), .CI(n240), .CO(n302), .S(n301) );
  OAI21XL U275 ( .A0(n90), .A1(n89), .B0(n88), .Y(n241) );
  INVXL U276 ( .A(n246), .Y(n89) );
  INVXL U277 ( .A(n91), .Y(n90) );
  XNOR2X1 U278 ( .A(n6), .B(n1129), .Y(n1149) );
  XNOR2XL U279 ( .A(n6), .B(B[24]), .Y(n1130) );
  XNOR2X1 U280 ( .A(n1100), .B(n1129), .Y(n1111) );
  XNOR2XL U281 ( .A(n1100), .B(B[24]), .Y(n1101) );
  OAI21XL U282 ( .A0(n299), .A1(n1161), .B0(n298), .Y(n1026) );
  ADDFX2 U283 ( .A(n260), .B(n62), .CI(n258), .CO(n296), .S(n295) );
  OAI22XL U284 ( .A0(n846), .A1(n261), .B0(n844), .B1(n252), .Y(n260) );
  AOI21XL U285 ( .A0(n1189), .A1(n1188), .B0(n293), .Y(n1161) );
  INVXL U286 ( .A(n1187), .Y(n293) );
  NAND2XL U287 ( .A(n303), .B(n302), .Y(n1028) );
  INVXL U288 ( .A(n1044), .Y(n363) );
  INVXL U289 ( .A(n1198), .Y(n1047) );
  NAND2X1 U290 ( .A(n47), .B(n906), .Y(n97) );
  INVXL U291 ( .A(n1220), .Y(n471) );
  AOI21XL U292 ( .A0(n470), .A1(n471), .B0(n430), .Y(n431) );
  INVXL U293 ( .A(n1221), .Y(n430) );
  XNOR2XL U294 ( .A(n6), .B(B[8]), .Y(n654) );
  XNOR2XL U295 ( .A(n6), .B(n807), .Y(n763) );
  XNOR2X1 U296 ( .A(B[18]), .B(n484), .Y(n108) );
  XNOR2X1 U297 ( .A(B[23]), .B(n484), .Y(n616) );
  XNOR2XL U298 ( .A(n68), .B(n6), .Y(n74) );
  INVXL U299 ( .A(n1253), .Y(n961) );
  NAND2BX1 U300 ( .AN(n1252), .B(n66), .Y(n65) );
  INVX1 U301 ( .A(n1254), .Y(n955) );
  NAND2XL U302 ( .A(n790), .B(n1239), .Y(n791) );
  XNOR2X1 U303 ( .A(n718), .B(n717), .Y(PRODUCT[24]) );
  NAND2XL U304 ( .A(n716), .B(n1235), .Y(n717) );
  INVXL U305 ( .A(n1234), .Y(n716) );
  XNOR2X1 U306 ( .A(n680), .B(n679), .Y(PRODUCT[25]) );
  NAND2XL U307 ( .A(n639), .B(n1233), .Y(n679) );
  INVXL U308 ( .A(n1232), .Y(n639) );
  XNOR2X1 U309 ( .A(n644), .B(n643), .Y(PRODUCT[26]) );
  NAND2XL U310 ( .A(n642), .B(n1231), .Y(n643) );
  INVXL U311 ( .A(n1230), .Y(n642) );
  XOR2X1 U312 ( .A(n368), .B(n59), .Y(PRODUCT[34]) );
  AND2XL U313 ( .A(n1033), .B(n1215), .Y(n59) );
  XNOR2X1 U314 ( .A(B[24]), .B(n82), .Y(n519) );
  XNOR2X1 U315 ( .A(B[23]), .B(n82), .Y(n556) );
  XNOR2XL U316 ( .A(n815), .B(B[18]), .Y(n594) );
  XNOR2X1 U317 ( .A(n1062), .B(B[13]), .Y(n625) );
  XNOR2XL U318 ( .A(n815), .B(B[16]), .Y(n664) );
  XNOR2XL U319 ( .A(n815), .B(n805), .Y(n699) );
  XNOR2XL U320 ( .A(n815), .B(B[14]), .Y(n738) );
  XNOR2XL U321 ( .A(n815), .B(B[13]), .Y(n773) );
  XNOR2XL U322 ( .A(n815), .B(B[12]), .Y(n816) );
  XOR2XL U323 ( .A(B[16]), .B(n437), .Y(n806) );
  XNOR2XL U324 ( .A(n815), .B(B[7]), .Y(n134) );
  NOR2BXL U325 ( .AN(B[0]), .B(n1134), .Y(n179) );
  OAI22XL U326 ( .A0(n1083), .A1(n328), .B0(n1081), .B1(n143), .Y(n177) );
  INVXL U327 ( .A(n1100), .Y(n133) );
  XNOR2X1 U328 ( .A(B[9]), .B(n484), .Y(n313) );
  XNOR2XL U329 ( .A(n438), .B(B[7]), .Y(n325) );
  XNOR2XL U330 ( .A(n438), .B(n1146), .Y(n439) );
  XNOR2XL U331 ( .A(n803), .B(B[21]), .Y(n449) );
  XNOR2XL U332 ( .A(n1100), .B(B[19]), .Y(n383) );
  XNOR2XL U333 ( .A(n815), .B(B[19]), .Y(n563) );
  XNOR2XL U334 ( .A(n1100), .B(B[16]), .Y(n479) );
  XNOR2XL U335 ( .A(n1062), .B(B[4]), .Y(n146) );
  NAND2BXL U336 ( .AN(B[0]), .B(n812), .Y(n254) );
  NAND2BXL U337 ( .AN(B[0]), .B(n815), .Y(n224) );
  XNOR2XL U338 ( .A(n803), .B(n1146), .Y(n1058) );
  OAI22XL U339 ( .A0(n861), .A1(n326), .B0(n859), .B1(n144), .Y(n974) );
  OAI22XL U340 ( .A0(n846), .A1(n331), .B0(n844), .B1(n330), .Y(n966) );
  XNOR2XL U341 ( .A(n6), .B(B[20]), .Y(n1057) );
  XNOR2XL U342 ( .A(n1062), .B(B[21]), .Y(n384) );
  OAI2BB1XL U343 ( .A0N(n859), .A1N(n700), .B0(n378), .Y(n395) );
  OAI22XL U344 ( .A0(n1150), .A1(n376), .B0(n1148), .B1(n392), .Y(n397) );
  INVXL U345 ( .A(n377), .Y(n378) );
  OAI22XL U346 ( .A0(n1060), .A1(n381), .B0(n1061), .B1(n393), .Y(n398) );
  OAI22XL U347 ( .A0(n1112), .A1(n379), .B0(n1134), .B1(n391), .Y(n400) );
  XNOR2XL U348 ( .A(n803), .B(B[22]), .Y(n411) );
  OAI2BB1XL U349 ( .A0N(n853), .A1N(n855), .B0(n373), .Y(n415) );
  OAI22XL U350 ( .A0(n1150), .A1(n409), .B0(n1148), .B1(n370), .Y(n417) );
  INVXL U351 ( .A(n372), .Y(n373) );
  CMPR32X1 U352 ( .A(n530), .B(n529), .C(n528), .CO(n522), .S(n580) );
  OAI2BB1XL U353 ( .A0N(n1032), .A1N(n801), .B0(n485), .Y(n528) );
  OAI22XL U354 ( .A0(n1112), .A1(n188), .B0(n1134), .B1(n848), .Y(n886) );
  INVXL U355 ( .A(n1195), .Y(n1196) );
  AOI21XL U356 ( .A0(n1194), .A1(n1193), .B0(n1192), .Y(n1195) );
  INVXL U357 ( .A(n1205), .Y(n1192) );
  NAND2XL U358 ( .A(n1193), .B(n1205), .Y(n1141) );
  NAND2XL U359 ( .A(n1036), .B(n1191), .Y(n1140) );
  NAND2X1 U360 ( .A(n110), .B(n109), .Y(n988) );
  NAND2XL U361 ( .A(n982), .B(n983), .Y(n109) );
  OAI2BB1XL U362 ( .A0N(n1109), .A1N(n1108), .B0(n1107), .Y(n1113) );
  OAI22XL U363 ( .A0(n1150), .A1(n1105), .B0(n1148), .B1(n1110), .Y(n1114) );
  INVXL U364 ( .A(n1106), .Y(n1107) );
  OAI22XL U365 ( .A0(n1112), .A1(n1079), .B0(n1134), .B1(n1101), .Y(n1104) );
  INVXL U366 ( .A(n1115), .Y(n1102) );
  OAI22XL U367 ( .A0(n1150), .A1(n1080), .B0(n1148), .B1(n1105), .Y(n1103) );
  OAI22XL U368 ( .A0(n1112), .A1(n1064), .B0(n1134), .B1(n1079), .Y(n1085) );
  OAI22XL U369 ( .A0(n1083), .A1(n1063), .B0(n1109), .B1(n1082), .Y(n1086) );
  OAI22XL U370 ( .A0(n861), .A1(n860), .B0(n859), .B1(n858), .Y(n898) );
  OAI22XL U371 ( .A0(n1083), .A1(n857), .B0(n1081), .B1(n856), .Y(n899) );
  OAI22XL U372 ( .A0(n861), .A1(n191), .B0(n859), .B1(n860), .Y(n892) );
  OAI22XL U373 ( .A0(n1083), .A1(n190), .B0(n1081), .B1(n857), .Y(n893) );
  OAI22XL U374 ( .A0(n1112), .A1(n848), .B0(n1134), .B1(n847), .Y(n895) );
  NOR2BXL U375 ( .AN(B[0]), .B(n853), .Y(n290) );
  OAI22XL U376 ( .A0(n846), .A1(n280), .B0(n844), .B1(n279), .Y(n288) );
  OAI22XL U377 ( .A0(n801), .A1(n278), .B0(n277), .B1(n1032), .Y(n289) );
  OAI22XL U378 ( .A0(n306), .A1(n263), .B0(n853), .B1(n262), .Y(n286) );
  OAI22XL U379 ( .A0(n846), .A1(n279), .B0(n844), .B1(n261), .Y(n287) );
  OAI22XL U380 ( .A0(n1150), .A1(n1149), .B0(n1148), .B1(n1147), .Y(n1151) );
  OAI2BB1XL U381 ( .A0N(n1134), .A1N(n1133), .B0(n1132), .Y(n1143) );
  OAI22XL U382 ( .A0(n1150), .A1(n1130), .B0(n1148), .B1(n1149), .Y(n1144) );
  INVXL U383 ( .A(n1131), .Y(n1132) );
  NAND2BX1 U384 ( .AN(n348), .B(n73), .Y(n1023) );
  AOI2BB1X1 U385 ( .A0N(n1027), .A1N(n1157), .B0(n71), .Y(n70) );
  OAI22XL U386 ( .A0(n801), .A1(B[0]), .B0(n266), .B1(n1032), .Y(n1184) );
  NAND2XL U387 ( .A(n267), .B(n801), .Y(n1183) );
  NAND2BXL U388 ( .AN(B[0]), .B(n484), .Y(n267) );
  NAND2XL U389 ( .A(n1184), .B(n1183), .Y(n1185) );
  NOR2XL U390 ( .A(n284), .B(n283), .Y(n1171) );
  AOI21XL U391 ( .A0(n1177), .A1(n273), .B0(n276), .Y(n1174) );
  INVXL U392 ( .A(n1176), .Y(n276) );
  NAND2XL U393 ( .A(n284), .B(n283), .Y(n1172) );
  NAND2XL U394 ( .A(n292), .B(n291), .Y(n1187) );
  NAND2X1 U395 ( .A(n296), .B(n297), .Y(n1163) );
  INVXL U396 ( .A(n1161), .Y(n1169) );
  INVXL U397 ( .A(n1137), .Y(n1094) );
  NOR2X1 U398 ( .A(n928), .B(n1253), .Y(n67) );
  INVXL U399 ( .A(n1241), .Y(n786) );
  INVXL U400 ( .A(n1217), .Y(n353) );
  XNOR2XL U401 ( .A(n6), .B(B[7]), .Y(n690) );
  XNOR2XL U402 ( .A(n6), .B(B[6]), .Y(n728) );
  NAND2BXL U403 ( .AN(B[0]), .B(A[13]), .Y(n132) );
  NAND2BXL U404 ( .AN(B[0]), .B(n1062), .Y(n175) );
  NAND2BXL U405 ( .AN(B[0]), .B(n803), .Y(n226) );
  XNOR2XL U406 ( .A(n6), .B(B[3]), .Y(n839) );
  INVXL U407 ( .A(n1215), .Y(n1038) );
  AOI21XL U408 ( .A0(n1092), .A1(n1091), .B0(n1090), .Y(n1138) );
  INVXL U409 ( .A(n1209), .Y(n1090) );
  INVXL U410 ( .A(n1138), .Y(n1093) );
  NAND2XL U411 ( .A(n1036), .B(n1094), .Y(n1096) );
  NAND2XL U412 ( .A(n1089), .B(n1091), .Y(n1137) );
  NAND2XL U413 ( .A(n1089), .B(n1211), .Y(n1049) );
  INVXL U414 ( .A(n1036), .Y(n1048) );
  XNOR2X2 U415 ( .A(n875), .B(n874), .Y(PRODUCT[20]) );
  NAND2X1 U416 ( .A(n97), .B(n1245), .Y(n875) );
  XOR2X2 U417 ( .A(n221), .B(n60), .Y(PRODUCT[33]) );
  OAI21XL U418 ( .A0(n1201), .A1(n220), .B0(n219), .Y(n221) );
  OAI21XL U419 ( .A0(n1201), .A1(n432), .B0(n431), .Y(n435) );
  INVXL U420 ( .A(n1218), .Y(n433) );
  XNOR2XL U421 ( .A(n812), .B(B[4]), .Y(n223) );
  OAI22X1 U422 ( .A0(n1032), .A1(n616), .B0(n653), .B1(n801), .Y(n652) );
  XNOR2X1 U423 ( .A(n68), .B(n1062), .Y(n698) );
  OAI22X1 U424 ( .A0(n762), .A1(n1032), .B0(n801), .B1(n108), .Y(n800) );
  XNOR2XL U425 ( .A(n1062), .B(B[0]), .Y(n329) );
  XNOR2XL U426 ( .A(n1062), .B(B[1]), .Y(n328) );
  XNOR2XL U427 ( .A(n812), .B(B[7]), .Y(n305) );
  XNOR2XL U428 ( .A(n803), .B(B[3]), .Y(n307) );
  XNOR2XL U429 ( .A(n438), .B(B[6]), .Y(n225) );
  XNOR2XL U430 ( .A(n6), .B(B[12]), .Y(n515) );
  XNOR2XL U431 ( .A(n815), .B(B[22]), .Y(n453) );
  XNOR2XL U432 ( .A(n803), .B(B[20]), .Y(n455) );
  XNOR2XL U433 ( .A(n6), .B(B[13]), .Y(n483) );
  OAI22X1 U434 ( .A0(n585), .A1(n1150), .B0(n74), .B1(n1148), .Y(n582) );
  OAI22X1 U435 ( .A0(n150), .A1(n801), .B0(n1032), .B1(n203), .Y(n202) );
  NAND2BXL U436 ( .AN(B[0]), .B(n6), .Y(n149) );
  OAI22XL U437 ( .A0(n1150), .A1(n204), .B0(n1148), .B1(n840), .Y(n884) );
  NAND2XL U438 ( .A(n1033), .B(n1039), .Y(n1041) );
  AOI21XL U439 ( .A0(n1039), .A1(n1038), .B0(n1037), .Y(n1040) );
  INVXL U440 ( .A(n1213), .Y(n1037) );
  NOR2XL U441 ( .A(n1216), .B(n1041), .Y(n1043) );
  INVX1 U442 ( .A(n1239), .Y(n104) );
  AOI21XL U443 ( .A0(n1198), .A1(n1191), .B0(n1194), .Y(n1139) );
  CMPR32X1 U444 ( .A(n318), .B(n317), .C(n316), .CO(n338), .S(n346) );
  OAI22XL U445 ( .A0(n855), .A1(n223), .B0(n853), .B1(n324), .Y(n316) );
  OAI22X1 U446 ( .A0(n1060), .A1(n222), .B0(n1061), .B1(n315), .Y(n317) );
  OAI22XL U447 ( .A0(n861), .A1(n229), .B0(n859), .B1(n322), .Y(n318) );
  NOR2BXL U448 ( .AN(B[0]), .B(n1061), .Y(n232) );
  OAI22XL U449 ( .A0(n861), .A1(n234), .B0(n859), .B1(n229), .Y(n230) );
  XNOR2X1 U450 ( .A(n984), .B(n78), .Y(n77) );
  XNOR2XL U451 ( .A(n1062), .B(n1146), .Y(n1106) );
  XNOR2XL U452 ( .A(n6), .B(B[22]), .Y(n1105) );
  XNOR2XL U453 ( .A(B[23]), .B(n1100), .Y(n1079) );
  ADDFX2 U454 ( .A(n566), .B(n565), .CI(n564), .CO(n558), .S(n612) );
  OAI22XL U455 ( .A0(n1112), .A1(n557), .B0(n1134), .B1(n521), .Y(n564) );
  OAI22XL U456 ( .A0(n846), .A1(n556), .B0(n520), .B1(n519), .Y(n565) );
  OAI22XL U457 ( .A0(n1060), .A1(n555), .B0(n1061), .B1(n518), .Y(n566) );
  OAI22XL U458 ( .A0(n861), .A1(n594), .B0(n859), .B1(n563), .Y(n598) );
  OAI22XL U459 ( .A0(n855), .A1(n592), .B0(n853), .B1(n561), .Y(n600) );
  ADDFX2 U460 ( .A(n597), .B(n596), .CI(n595), .CO(n589), .S(n649) );
  OAI22XL U461 ( .A0(n1112), .A1(n588), .B0(n1134), .B1(n557), .Y(n595) );
  OAI22X1 U462 ( .A0(n846), .A1(n587), .B0(n844), .B1(n556), .Y(n596) );
  CMPR32X1 U463 ( .A(n632), .B(n631), .C(n630), .CO(n650), .S(n684) );
  OAI22XL U464 ( .A0(n1083), .A1(n625), .B0(n1081), .B1(n593), .Y(n631) );
  OAI22XL U465 ( .A0(n855), .A1(n624), .B0(n853), .B1(n592), .Y(n632) );
  ADDFX2 U466 ( .A(n629), .B(n628), .CI(n627), .CO(n621), .S(n685) );
  OAI22XL U467 ( .A0(n1112), .A1(n620), .B0(n1134), .B1(n588), .Y(n627) );
  ADDFX2 U468 ( .A(n661), .B(n660), .CI(n659), .CO(n673), .S(n708) );
  CMPR32X1 U469 ( .A(n670), .B(n669), .C(n668), .CO(n686), .S(n722) );
  OAI22XL U470 ( .A0(n1083), .A1(n663), .B0(n1081), .B1(n625), .Y(n669) );
  OAI22XL U471 ( .A0(n855), .A1(n662), .B0(n853), .B1(n624), .Y(n670) );
  OAI22XL U472 ( .A0(n861), .A1(n699), .B0(n859), .B1(n664), .Y(n704) );
  ADDFX2 U473 ( .A(n703), .B(n702), .CI(n701), .CO(n694), .S(n758) );
  OAI22XL U474 ( .A0(n1112), .A1(n693), .B0(n1134), .B1(n658), .Y(n701) );
  OAI22X1 U475 ( .A0(n846), .A1(n692), .B0(n844), .B1(n657), .Y(n702) );
  OAI22XL U476 ( .A0(n656), .A1(n691), .B0(n1061), .B1(n655), .Y(n703) );
  OAI22XL U477 ( .A0(n1112), .A1(n732), .B0(n1134), .B1(n693), .Y(n739) );
  OAI22XL U478 ( .A0(n846), .A1(n730), .B0(n844), .B1(n692), .Y(n740) );
  OAI22XL U479 ( .A0(n861), .A1(n773), .B0(n859), .B1(n738), .Y(n777) );
  OAI22XL U480 ( .A0(n1112), .A1(n767), .B0(n1134), .B1(n732), .Y(n774) );
  CMPR32X1 U481 ( .A(n819), .B(n818), .C(n817), .CO(n809), .S(n880) );
  OAI22XL U482 ( .A0(n1112), .A1(n808), .B0(n1134), .B1(n767), .Y(n817) );
  OAI22XL U483 ( .A0(n1060), .A1(n804), .B0(n1061), .B1(n765), .Y(n819) );
  OAI22XL U484 ( .A0(n861), .A1(n816), .B0(n859), .B1(n773), .Y(n820) );
  OAI22XL U485 ( .A0(n861), .A1(n858), .B0(n859), .B1(n816), .Y(n865) );
  OAI22XL U486 ( .A0(n1083), .A1(n856), .B0(n1081), .B1(n814), .Y(n866) );
  OAI22XL U487 ( .A0(n1112), .A1(n847), .B0(n1134), .B1(n808), .Y(n862) );
  OAI22XL U488 ( .A0(n1112), .A1(n152), .B0(n1134), .B1(n188), .Y(n198) );
  OAI22XL U489 ( .A0(n1150), .A1(n124), .B0(n1148), .B1(n204), .Y(n199) );
  NOR2BXL U490 ( .AN(B[0]), .B(n1148), .Y(n156) );
  OAI22XL U491 ( .A0(n1112), .A1(n153), .B0(n1134), .B1(n152), .Y(n154) );
  OAI22X1 U492 ( .A0(n801), .A1(n151), .B0(n150), .B1(n1032), .Y(n155) );
  ADDFX2 U493 ( .A(n164), .B(n163), .CI(n162), .CO(n207), .S(n165) );
  OAI22X1 U494 ( .A0(n1083), .A1(n136), .B0(n1081), .B1(n146), .Y(n163) );
  OAI22XL U495 ( .A0(n656), .A1(n157), .B0(n1061), .B1(n121), .Y(n164) );
  CMPR32X1 U496 ( .A(n139), .B(n138), .C(n137), .CO(n205), .S(n181) );
  OAI22XL U497 ( .A0(n1083), .A1(n143), .B0(n1081), .B1(n136), .Y(n168) );
  OAI22XL U498 ( .A0(n1112), .A1(n135), .B0(n1134), .B1(n153), .Y(n169) );
  OAI22XL U499 ( .A0(n861), .A1(n144), .B0(n859), .B1(n134), .Y(n170) );
  NOR2BXL U500 ( .AN(B[0]), .B(n1081), .Y(n321) );
  OAI22XL U501 ( .A0(n656), .A1(n315), .B0(n1061), .B1(n314), .Y(n319) );
  OAI22X1 U502 ( .A0(n801), .A1(n313), .B0(n312), .B1(n1032), .Y(n320) );
  ADDFX2 U503 ( .A(n334), .B(n333), .CI(n332), .CO(n982), .S(n343) );
  OAI22XL U504 ( .A0(n846), .A1(n325), .B0(n844), .B1(n331), .Y(n332) );
  OAI22XL U505 ( .A0(n855), .A1(n324), .B0(n853), .B1(n323), .Y(n333) );
  OAI2BB1XL U506 ( .A0N(n520), .A1N(n731), .B0(n440), .Y(n456) );
  OAI22XL U507 ( .A0(n1060), .A1(n449), .B0(n1061), .B1(n411), .Y(n441) );
  OAI22XL U508 ( .A0(n1083), .A1(n407), .B0(n1081), .B1(n384), .Y(n412) );
  OAI22XL U509 ( .A0(n1133), .A1(n410), .B0(n1134), .B1(n383), .Y(n413) );
  OAI22XL U510 ( .A0(n861), .A1(n408), .B0(n859), .B1(n382), .Y(n414) );
  OAI22XL U511 ( .A0(n1133), .A1(n383), .B0(n1134), .B1(n379), .Y(n387) );
  OAI22XL U512 ( .A0(n861), .A1(n563), .B0(n859), .B1(n527), .Y(n567) );
  OAI22XL U513 ( .A0(n855), .A1(n561), .B0(n853), .B1(n525), .Y(n569) );
  CMPR32X1 U514 ( .A(n623), .B(n622), .C(n621), .CO(n635), .S(n672) );
  CMPR32X1 U515 ( .A(n496), .B(n495), .C(n494), .CO(n513), .S(n549) );
  OAI22XL U516 ( .A0(n1060), .A1(n482), .B0(n1061), .B1(n455), .Y(n494) );
  OAI22XL U517 ( .A0(n1150), .A1(n483), .B0(n1148), .B1(n454), .Y(n495) );
  OAI22XL U518 ( .A0(n861), .A1(n480), .B0(n859), .B1(n453), .Y(n496) );
  OAI22X1 U519 ( .A0(n1083), .A1(n489), .B0(n1081), .B1(n451), .Y(n493) );
  OAI22XL U520 ( .A0(n855), .A1(n490), .B0(n853), .B1(n452), .Y(n492) );
  OAI22XL U521 ( .A0(n1108), .A1(n526), .B0(n1081), .B1(n489), .Y(n532) );
  OAI22XL U522 ( .A0(n1133), .A1(n481), .B0(n1134), .B1(n479), .Y(n524) );
  OR2XL U523 ( .A(n516), .B(n517), .Y(n523) );
  XNOR2XL U524 ( .A(n1062), .B(B[7]), .Y(n856) );
  XNOR2XL U525 ( .A(n68), .B(n815), .Y(n858) );
  XNOR2XL U526 ( .A(n1062), .B(B[6]), .Y(n857) );
  XNOR2X1 U527 ( .A(n815), .B(B[10]), .Y(n860) );
  XNOR2X1 U528 ( .A(n68), .B(n812), .Y(n189) );
  XNOR2XL U529 ( .A(n805), .B(n82), .Y(n843) );
  XNOR2XL U530 ( .A(n803), .B(B[9]), .Y(n841) );
  XNOR2XL U531 ( .A(n803), .B(B[8]), .Y(n842) );
  OAI22XL U532 ( .A0(n861), .A1(n147), .B0(n859), .B1(n191), .Y(n183) );
  OAI22XL U533 ( .A0(n1083), .A1(n146), .B0(n1081), .B1(n190), .Y(n184) );
  XNOR2X1 U534 ( .A(A[2]), .B(A[1]), .Y(n520) );
  OAI22XL U535 ( .A0(n855), .A1(n371), .B0(n853), .B1(n254), .Y(n264) );
  XNOR2XL U536 ( .A(n438), .B(B[3]), .Y(n261) );
  NOR2BXL U537 ( .AN(B[0]), .B(n859), .Y(n257) );
  OAI22XL U538 ( .A0(n855), .A1(n262), .B0(n853), .B1(n248), .Y(n255) );
  XNOR2XL U539 ( .A(n815), .B(B[0]), .Y(n235) );
  OAI22XL U540 ( .A0(n861), .A1(n375), .B0(n859), .B1(n224), .Y(n243) );
  INVXL U541 ( .A(n815), .Y(n375) );
  OAI2BB1XL U542 ( .A0N(n1061), .A1N(n1060), .B0(n1059), .Y(n1076) );
  OAI22XL U543 ( .A0(n1150), .A1(n1057), .B0(n1148), .B1(n1080), .Y(n1078) );
  INVXL U544 ( .A(n1058), .Y(n1059) );
  ADDFX2 U545 ( .A(n499), .B(n498), .CI(n497), .CO(n474), .S(n508) );
  ADDFX2 U546 ( .A(n686), .B(n685), .CI(n684), .CO(n671), .S(n721) );
  OR2X2 U547 ( .A(n829), .B(n830), .Y(n94) );
  ADDFX2 U548 ( .A(n870), .B(n869), .CI(n868), .CO(n829), .S(n876) );
  ADDFX2 U549 ( .A(n833), .B(n832), .CI(n831), .CO(n823), .S(n878) );
  ADDFX2 U550 ( .A(n881), .B(n880), .CI(n879), .CO(n868), .S(n910) );
  ADDFX2 U551 ( .A(n903), .B(n902), .CI(n901), .CO(n877), .S(n908) );
  OAI21XL U552 ( .A0(n933), .A1(n934), .B0(n932), .Y(n80) );
  ADDFX2 U553 ( .A(n167), .B(n166), .CI(n165), .CO(n192), .S(n996) );
  NAND2X1 U554 ( .A(n76), .B(n75), .Y(n998) );
  OAI21XL U555 ( .A0(n985), .A1(n986), .B0(n984), .Y(n76) );
  OAI22XL U556 ( .A0(n1112), .A1(n391), .B0(n1134), .B1(n1064), .Y(n1067) );
  OAI22XL U557 ( .A0(n1150), .A1(n392), .B0(n1148), .B1(n1057), .Y(n1066) );
  INVXL U558 ( .A(n1077), .Y(n1065) );
  OAI22XL U559 ( .A0(n1083), .A1(n394), .B0(n1109), .B1(n1063), .Y(n1070) );
  OAI22XL U560 ( .A0(n1083), .A1(n384), .B0(n1081), .B1(n380), .Y(n390) );
  OAI22XL U561 ( .A0(n1150), .A1(n370), .B0(n1148), .B1(n376), .Y(n389) );
  ADDFX2 U562 ( .A(n464), .B(n463), .CI(n462), .CO(n466), .S(n473) );
  CMPR32X1 U563 ( .A(n423), .B(n422), .C(n421), .CO(n424), .S(n465) );
  OAI22XL U564 ( .A0(n801), .A1(n266), .B0(n270), .B1(n1032), .Y(n269) );
  NOR2BXL U565 ( .AN(B[0]), .B(n844), .Y(n268) );
  OAI22XL U566 ( .A0(n846), .A1(n437), .B0(n520), .B1(n272), .Y(n274) );
  NAND2BXL U567 ( .AN(B[0]), .B(n438), .Y(n272) );
  NAND2XL U568 ( .A(n1036), .B(n1197), .Y(n1200) );
  AOI21XL U569 ( .A0(n1198), .A1(n1197), .B0(n1196), .Y(n1199) );
  XOR3X2 U570 ( .A(n475), .B(n473), .C(n474), .Y(n501) );
  OAI22XL U571 ( .A0(n1150), .A1(n1110), .B0(n1148), .B1(n1130), .Y(n1128) );
  INVXL U572 ( .A(n1145), .Y(n1127) );
  OAI22XL U573 ( .A0(n1112), .A1(n1101), .B0(n1134), .B1(n1111), .Y(n1123) );
  ADDFX2 U574 ( .A(n1075), .B(n1074), .CI(n1073), .CO(n1088), .S(n1071) );
  OAI21XL U575 ( .A0(n101), .A1(n100), .B0(n99), .Y(n469) );
  OAI21XL U576 ( .A0(n474), .A1(n475), .B0(n473), .Y(n99) );
  OAI21XL U577 ( .A0(n96), .A1(n95), .B0(n93), .Y(n826) );
  NAND2X1 U578 ( .A(n94), .B(n828), .Y(n93) );
  XOR3X2 U579 ( .A(n830), .B(n829), .C(n828), .Y(n872) );
  OAI21XL U580 ( .A0(n107), .A1(n106), .B0(n105), .Y(n871) );
  OAI21XL U581 ( .A0(n877), .A1(n878), .B0(n876), .Y(n105) );
  OAI2BB1X1 U582 ( .A0N(n910), .A1N(n909), .B0(n87), .Y(n904) );
  OAI21XL U583 ( .A0(n909), .A1(n910), .B0(n908), .Y(n87) );
  XOR3X2 U584 ( .A(n878), .B(n876), .C(n877), .Y(n905) );
  XOR3X2 U585 ( .A(n910), .B(n908), .C(n909), .Y(n927) );
  ADDFX2 U586 ( .A(n996), .B(n995), .CI(n994), .CO(n956), .S(n1006) );
  NAND2XL U587 ( .A(n212), .B(n211), .Y(n959) );
  AOI21X1 U588 ( .A0(n57), .A1(n1016), .B0(n1004), .Y(n1010) );
  XNOR3X2 U589 ( .A(n934), .B(n932), .C(n81), .Y(n949) );
  OAI21XL U590 ( .A0(n942), .A1(n943), .B0(n941), .Y(n83) );
  NOR2XL U591 ( .A(n269), .B(n268), .Y(n1179) );
  NAND2XL U592 ( .A(n269), .B(n268), .Y(n1180) );
  NAND2XL U593 ( .A(n275), .B(n274), .Y(n1176) );
  NOR2X1 U594 ( .A(n957), .B(n956), .Y(mult_x_1_n312) );
  NOR2XL U595 ( .A(n1072), .B(n1071), .Y(mult_x_1_n149) );
  NAND2XL U596 ( .A(n1158), .B(n1157), .Y(n1159) );
  INVXL U597 ( .A(n1156), .Y(n1158) );
  NAND2XL U598 ( .A(n1029), .B(n1028), .Y(n1030) );
  NAND2XL U599 ( .A(n1020), .B(n1019), .Y(n1021) );
  AOI21XL U600 ( .A0(n1025), .A1(n1023), .B0(n1018), .Y(n92) );
  NAND2XL U601 ( .A(n1155), .B(n1154), .Y(mult_x_1_n54) );
  NAND2XL U602 ( .A(n1153), .B(n1152), .Y(n1154) );
  INVXL U603 ( .A(n1151), .Y(n1152) );
  NOR2XL U604 ( .A(n1136), .B(n1135), .Y(mult_x_1_n105) );
  NAND2XL U605 ( .A(n1136), .B(n1135), .Y(mult_x_1_n106) );
  NOR2XL U606 ( .A(n1117), .B(n1116), .Y(mult_x_1_n114) );
  NAND2XL U607 ( .A(n1117), .B(n1116), .Y(mult_x_1_n115) );
  NOR2XL U608 ( .A(n1125), .B(n1124), .Y(mult_x_1_n125) );
  NAND2XL U609 ( .A(n1125), .B(n1124), .Y(mult_x_1_n126) );
  NOR2XL U610 ( .A(n1088), .B(n1087), .Y(mult_x_1_n134) );
  NAND2XL U611 ( .A(n1088), .B(n1087), .Y(mult_x_1_n135) );
  NAND2XL U612 ( .A(n1072), .B(n1071), .Y(mult_x_1_n150) );
  NOR2X1 U613 ( .A(n951), .B(n950), .Y(mult_x_1_n299) );
  NAND2X1 U614 ( .A(n72), .B(n69), .Y(mult_x_1_n335) );
  AOI21XL U615 ( .A0(n1018), .A1(n1020), .B0(n351), .Y(n72) );
  NOR2BXL U616 ( .AN(B[0]), .B(n1032), .Y(n1288) );
  XOR2XL U617 ( .A(n1182), .B(n1185), .Y(n1286) );
  NAND2XL U618 ( .A(n1181), .B(n1180), .Y(n1182) );
  INVXL U619 ( .A(n1179), .Y(n1181) );
  XNOR2XL U620 ( .A(n1178), .B(n1177), .Y(n1285) );
  NAND2XL U621 ( .A(n273), .B(n1176), .Y(n1178) );
  XOR2XL U622 ( .A(n1175), .B(n1174), .Y(n1284) );
  NAND2XL U623 ( .A(n1173), .B(n1172), .Y(n1175) );
  INVXL U624 ( .A(n1171), .Y(n1173) );
  NAND2XL U625 ( .A(n1188), .B(n1187), .Y(n1190) );
  XOR2XL U626 ( .A(n1166), .B(n1165), .Y(n1281) );
  NAND2XL U627 ( .A(n1164), .B(n1163), .Y(n1165) );
  BUFX3 U628 ( .A(A[11]), .Y(n1062) );
  BUFX3 U629 ( .A(A[9]), .Y(n803) );
  OR2X2 U630 ( .A(n1003), .B(n1002), .Y(n57) );
  BUFX3 U631 ( .A(A[7]), .Y(n815) );
  OAI22X1 U632 ( .A0(n838), .A1(n554), .B0(n514), .B1(n1032), .Y(n553) );
  OAI22X1 U633 ( .A0(n764), .A1(n617), .B0(n1148), .B1(n585), .Y(n614) );
  OAI22X1 U634 ( .A0(n764), .A1(n654), .B0(n1148), .B1(n617), .Y(n651) );
  OAI22X1 U635 ( .A0(n764), .A1(n690), .B0(n1148), .B1(n654), .Y(n687) );
  OAI22X1 U636 ( .A0(n1150), .A1(n515), .B0(n1148), .B1(n483), .Y(n529) );
  ADDFX2 U637 ( .A(n744), .B(n743), .CI(n742), .CO(n759), .S(n796) );
  XNOR2X1 U638 ( .A(n815), .B(B[21]), .Y(n480) );
  XNOR2XL U639 ( .A(B[23]), .B(n6), .Y(n1110) );
  OAI22X1 U640 ( .A0(n700), .A1(n382), .B0(n859), .B1(n377), .Y(n396) );
  BUFX1 U641 ( .A(n259), .Y(n62) );
  CMPR22X1 U642 ( .A(n583), .B(n582), .CO(n590), .S(n623) );
  CMPR22X1 U643 ( .A(n553), .B(n552), .CO(n560), .S(n591) );
  OAI22X1 U644 ( .A0(n515), .A1(n1148), .B0(n1150), .B1(n74), .Y(n552) );
  CMPR22X1 U645 ( .A(n835), .B(n834), .CO(n850), .S(n891) );
  OAI22X1 U646 ( .A0(n836), .A1(n801), .B0(n1032), .B1(n108), .Y(n835) );
  XNOR2X1 U647 ( .A(n68), .B(n803), .Y(n765) );
  OAI22X1 U648 ( .A0(n846), .A1(n225), .B0(n844), .B1(n325), .Y(n337) );
  XNOR2X2 U649 ( .A(n545), .B(n544), .Y(PRODUCT[29]) );
  NAND2X1 U650 ( .A(n543), .B(n1225), .Y(n544) );
  XNOR2X1 U651 ( .A(n792), .B(n791), .Y(PRODUCT[22]) );
  OAI22X1 U652 ( .A0(n844), .A1(n619), .B0(n657), .B1(n731), .Y(n666) );
  OAI21XL U653 ( .A0(n955), .A1(n67), .B0(n1252), .Y(n64) );
  OAI21X2 U654 ( .A0(n955), .A1(n65), .B0(n64), .Y(PRODUCT[16]) );
  XNOR2X1 U655 ( .A(n68), .B(A[13]), .Y(n620) );
  BUFX4 U656 ( .A(B[11]), .Y(n68) );
  XNOR2X1 U657 ( .A(n68), .B(n438), .Y(n158) );
  NOR2BX1 U658 ( .AN(n348), .B(n73), .Y(n1018) );
  NAND2X1 U659 ( .A(n1003), .B(n1002), .Y(n1012) );
  XNOR2X1 U660 ( .A(B[20]), .B(n82), .Y(n657) );
  XNOR2X1 U661 ( .A(B[19]), .B(n82), .Y(n692) );
  XNOR2X1 U662 ( .A(B[21]), .B(n82), .Y(n619) );
  XNOR2X1 U663 ( .A(n805), .B(n484), .Y(n203) );
  XNOR2X1 U664 ( .A(B[25]), .B(n484), .Y(n554) );
  NAND2BX1 U665 ( .AN(n297), .B(n86), .Y(n1164) );
  OAI21XL U666 ( .A0(n246), .A1(n91), .B0(n245), .Y(n88) );
  XOR3X2 U667 ( .A(n246), .B(n91), .C(n245), .Y(n250) );
  OAI22X2 U668 ( .A0(n233), .A1(n844), .B0(n846), .B1(n252), .Y(n91) );
  XNOR2X1 U669 ( .A(B[22]), .B(n484), .Y(n653) );
  OAI21XL U670 ( .A0(n715), .A1(n98), .B0(n714), .Y(n718) );
  OAI21XL U671 ( .A0(n678), .A1(n98), .B0(n677), .Y(n680) );
  BUFX3 U672 ( .A(B[25]), .Y(n1129) );
  INVX1 U673 ( .A(mult_x_1_n335), .Y(n1017) );
  AOI21X1 U674 ( .A0(n112), .A1(n787), .B0(n786), .Y(n788) );
  INVX1 U675 ( .A(n218), .Y(n470) );
  XNOR2X1 U676 ( .A(B[23]), .B(n815), .Y(n448) );
  XNOR2X1 U677 ( .A(B[23]), .B(n812), .Y(n490) );
  XNOR2X1 U678 ( .A(B[23]), .B(n803), .Y(n406) );
  XNOR2X1 U679 ( .A(B[23]), .B(n1062), .Y(n394) );
  XOR2X1 U680 ( .A(n962), .B(n928), .Y(PRODUCT[15]) );
  XOR3X2 U681 ( .A(n983), .B(n982), .C(n981), .Y(n990) );
  OAI22X1 U682 ( .A0(n801), .A1(n228), .B0(n227), .B1(n1032), .Y(n231) );
  OAI22X1 U683 ( .A0(n1060), .A1(n655), .B0(n1061), .B1(n618), .Y(n667) );
  CMPR22X1 U684 ( .A(n141), .B(n140), .CO(n137), .S(n965) );
  OAI22X1 U685 ( .A0(n801), .A1(n142), .B0(n151), .B1(n1032), .Y(n141) );
  OAI22X1 U686 ( .A0(n846), .A1(n187), .B0(n844), .B1(n845), .Y(n887) );
  OAI22X1 U687 ( .A0(n838), .A1(n837), .B0(n836), .B1(n1032), .Y(n883) );
  NOR2X1 U688 ( .A(n640), .B(n214), .Y(n215) );
  OAI22X1 U689 ( .A0(n846), .A1(n845), .B0(n844), .B1(n843), .Y(n896) );
  OAI22X1 U690 ( .A0(n801), .A1(n312), .B0(n174), .B1(n1032), .Y(n309) );
  XNOR2X1 U691 ( .A(A[13]), .B(n807), .Y(n847) );
  NOR2X2 U692 ( .A(n1244), .B(n1242), .Y(n785) );
  INVXL U693 ( .A(n785), .Y(n114) );
  NAND2X1 U694 ( .A(n787), .B(n1241), .Y(n115) );
  XNOR2X2 U695 ( .A(n116), .B(n115), .Y(PRODUCT[21]) );
  XOR2XL U696 ( .A(A[8]), .B(A[9]), .Y(n117) );
  XNOR2X1 U697 ( .A(n803), .B(n807), .Y(n157) );
  BUFX3 U698 ( .A(n118), .Y(n1061) );
  XNOR2X1 U699 ( .A(n803), .B(B[6]), .Y(n121) );
  XOR2XL U700 ( .A(A[10]), .B(A[11]), .Y(n119) );
  BUFX3 U701 ( .A(n1108), .Y(n1083) );
  INVXL U702 ( .A(n1062), .Y(n176) );
  BUFX3 U703 ( .A(n1109), .Y(n1081) );
  NAND2X1 U704 ( .A(n120), .B(n520), .Y(n731) );
  BUFX3 U705 ( .A(n731), .Y(n846) );
  BUFX3 U706 ( .A(n520), .Y(n844) );
  XNOR2X1 U707 ( .A(n438), .B(B[12]), .Y(n145) );
  OAI22XL U708 ( .A0(n846), .A1(n158), .B0(n844), .B1(n145), .Y(n162) );
  XNOR2X1 U709 ( .A(n803), .B(B[7]), .Y(n186) );
  XOR2XL U710 ( .A(A[14]), .B(A[15]), .Y(n122) );
  XNOR2XL U711 ( .A(A[14]), .B(A[13]), .Y(n123) );
  NAND2X1 U712 ( .A(n122), .B(n123), .Y(n764) );
  BUFX3 U713 ( .A(n764), .Y(n1150) );
  INVX1 U714 ( .A(A[15]), .Y(n369) );
  BUFX3 U715 ( .A(n123), .Y(n1148) );
  XNOR2XL U716 ( .A(n6), .B(B[1]), .Y(n204) );
  XOR2XL U717 ( .A(A[12]), .B(A[13]), .Y(n125) );
  XNOR2XL U718 ( .A(A[12]), .B(A[11]), .Y(n126) );
  BUFX3 U719 ( .A(n1133), .Y(n1112) );
  XNOR2XL U720 ( .A(n1100), .B(B[2]), .Y(n152) );
  BUFX3 U721 ( .A(n126), .Y(n1134) );
  XNOR2X1 U722 ( .A(A[13]), .B(B[3]), .Y(n188) );
  XOR2XL U723 ( .A(A[4]), .B(A[5]), .Y(n127) );
  XNOR2XL U724 ( .A(A[4]), .B(A[3]), .Y(n128) );
  BUFX3 U725 ( .A(n306), .Y(n855) );
  XNOR2X1 U726 ( .A(n812), .B(B[9]), .Y(n160) );
  BUFX3 U727 ( .A(n128), .Y(n853) );
  XNOR2X1 U728 ( .A(n812), .B(B[10]), .Y(n148) );
  OAI22XL U729 ( .A0(n855), .A1(n160), .B0(n853), .B1(n148), .Y(n139) );
  XOR2XL U730 ( .A(A[6]), .B(A[7]), .Y(n129) );
  XNOR2XL U731 ( .A(A[6]), .B(A[5]), .Y(n130) );
  NAND2X1 U732 ( .A(n129), .B(n130), .Y(n700) );
  BUFX3 U733 ( .A(n700), .Y(n861) );
  BUFX3 U734 ( .A(n130), .Y(n859) );
  XNOR2X1 U735 ( .A(n815), .B(B[8]), .Y(n147) );
  OAI22XL U736 ( .A0(n861), .A1(n134), .B0(n859), .B1(n147), .Y(n138) );
  NAND2X1 U737 ( .A(A[1]), .B(n131), .Y(n838) );
  BUFX3 U738 ( .A(n838), .Y(n801) );
  XNOR2X1 U739 ( .A(n484), .B(B[13]), .Y(n151) );
  BUFX3 U740 ( .A(n131), .Y(n1032) );
  OAI22X1 U741 ( .A0(n1112), .A1(n133), .B0(n1134), .B1(n132), .Y(n140) );
  XNOR2XL U742 ( .A(n1100), .B(B[0]), .Y(n135) );
  XNOR2XL U743 ( .A(n1100), .B(B[1]), .Y(n153) );
  XNOR2XL U744 ( .A(n1062), .B(B[2]), .Y(n143) );
  XNOR2X1 U745 ( .A(n438), .B(B[9]), .Y(n330) );
  XNOR2X1 U746 ( .A(n438), .B(B[10]), .Y(n159) );
  OAI22XL U747 ( .A0(n846), .A1(n330), .B0(n844), .B1(n159), .Y(n973) );
  OAI22XL U748 ( .A0(n855), .A1(n305), .B0(n853), .B1(n161), .Y(n972) );
  XNOR2X1 U749 ( .A(n438), .B(B[13]), .Y(n187) );
  XNOR2X1 U750 ( .A(n1062), .B(n807), .Y(n190) );
  OAI22XL U751 ( .A0(n855), .A1(n148), .B0(n853), .B1(n189), .Y(n197) );
  XNOR2X1 U752 ( .A(n484), .B(B[14]), .Y(n150) );
  BUFX3 U753 ( .A(B[15]), .Y(n805) );
  OAI22X1 U754 ( .A0(n1150), .A1(n369), .B0(n1148), .B1(n149), .Y(n201) );
  ADDFHX1 U755 ( .A(n156), .B(n155), .CI(n154), .CO(n195), .S(n167) );
  BUFX3 U756 ( .A(n656), .Y(n1060) );
  XNOR2XL U757 ( .A(n803), .B(B[4]), .Y(n173) );
  OAI22XL U758 ( .A0(n306), .A1(n161), .B0(n853), .B1(n160), .Y(n171) );
  CMPR32X1 U759 ( .A(n170), .B(n169), .C(n168), .CO(n182), .S(n977) );
  XNOR2X1 U760 ( .A(n484), .B(B[10]), .Y(n312) );
  OAI22X1 U761 ( .A0(n1083), .A1(n176), .B0(n1081), .B1(n175), .Y(n308) );
  ADDFHX1 U762 ( .A(n179), .B(n178), .CI(n177), .CO(n964), .S(n978) );
  CMPR32X1 U763 ( .A(n182), .B(n181), .C(n180), .CO(n209), .S(n994) );
  CMPR32X1 U764 ( .A(n185), .B(n184), .C(n183), .CO(n922), .S(n194) );
  OAI22X1 U765 ( .A0(n1060), .A1(n186), .B0(n1061), .B1(n842), .Y(n888) );
  XNOR2X1 U766 ( .A(n438), .B(B[14]), .Y(n845) );
  XNOR2XL U767 ( .A(A[13]), .B(B[4]), .Y(n848) );
  XNOR2X1 U768 ( .A(n812), .B(B[12]), .Y(n854) );
  OAI22XL U769 ( .A0(n855), .A1(n189), .B0(n853), .B1(n854), .Y(n894) );
  CMPR32X1 U770 ( .A(n197), .B(n196), .C(n195), .CO(n937), .S(n193) );
  CMPR32X1 U771 ( .A(n200), .B(n199), .C(n198), .CO(n916), .S(n206) );
  CMPR22X1 U772 ( .A(n202), .B(n201), .CO(n915), .S(n196) );
  XNOR2X1 U773 ( .A(n484), .B(B[16]), .Y(n837) );
  OAI22XL U774 ( .A0(n838), .A1(n203), .B0(n837), .B1(n1032), .Y(n885) );
  XNOR2XL U775 ( .A(n6), .B(B[2]), .Y(n840) );
  CMPR32X1 U776 ( .A(n207), .B(n206), .C(n205), .CO(n935), .S(n210) );
  CMPR32X1 U777 ( .A(n210), .B(n209), .C(n208), .CO(n211), .S(n957) );
  NOR2X1 U778 ( .A(n1228), .B(n1226), .Y(n539) );
  INVX1 U779 ( .A(n1035), .Y(n429) );
  NOR2XL U780 ( .A(n1220), .B(n1218), .Y(n1034) );
  INVXL U781 ( .A(n1034), .Y(n362) );
  NAND2XL U782 ( .A(n429), .B(n1034), .Y(n220) );
  OAI21X1 U783 ( .A0(n1226), .A1(n1229), .B0(n1227), .Y(n540) );
  OAI21XL U784 ( .A0(n1222), .A1(n1225), .B0(n1223), .Y(n216) );
  OAI21XL U785 ( .A0(n1218), .A1(n1221), .B0(n1219), .Y(n1044) );
  INVXL U786 ( .A(n1216), .Y(n352) );
  XNOR2XL U787 ( .A(n815), .B(B[2]), .Y(n229) );
  XNOR2X1 U788 ( .A(n815), .B(B[3]), .Y(n322) );
  XNOR2XL U789 ( .A(n803), .B(B[0]), .Y(n222) );
  XNOR2XL U790 ( .A(n803), .B(B[1]), .Y(n315) );
  XNOR2X1 U791 ( .A(n812), .B(n807), .Y(n324) );
  OAI22XL U792 ( .A0(n846), .A1(n233), .B0(n844), .B1(n225), .Y(n239) );
  XNOR2X1 U793 ( .A(n812), .B(B[3]), .Y(n236) );
  OAI22XL U794 ( .A0(n306), .A1(n236), .B0(n853), .B1(n223), .Y(n238) );
  XNOR2X1 U795 ( .A(n484), .B(B[6]), .Y(n247) );
  XNOR2X1 U796 ( .A(n484), .B(B[7]), .Y(n228) );
  OAI22XL U797 ( .A0(n801), .A1(n247), .B0(n228), .B1(n1032), .Y(n244) );
  XNOR2X1 U798 ( .A(n484), .B(B[8]), .Y(n227) );
  OAI22X1 U799 ( .A0(n801), .A1(n227), .B0(n313), .B1(n1032), .Y(n311) );
  INVXL U800 ( .A(n803), .Y(n374) );
  OAI22X1 U801 ( .A0(n1060), .A1(n374), .B0(n1061), .B1(n226), .Y(n310) );
  XNOR2XL U802 ( .A(n815), .B(B[1]), .Y(n234) );
  CMPR32X1 U803 ( .A(n232), .B(n231), .C(n230), .CO(n335), .S(n242) );
  XNOR2XL U804 ( .A(n438), .B(B[4]), .Y(n252) );
  OAI22X1 U805 ( .A0(n861), .A1(n235), .B0(n859), .B1(n234), .Y(n246) );
  XNOR2XL U806 ( .A(n812), .B(B[2]), .Y(n248) );
  OAI22X1 U807 ( .A0(n855), .A1(n248), .B0(n853), .B1(n236), .Y(n245) );
  CMPR32X1 U808 ( .A(n239), .B(n238), .C(n237), .CO(n345), .S(n240) );
  ADDHXL U809 ( .A(n244), .B(n243), .CO(n237), .S(n251) );
  XNOR2X1 U810 ( .A(n484), .B(n807), .Y(n253) );
  OAI22XL U811 ( .A0(n801), .A1(n253), .B0(n247), .B1(n1032), .Y(n256) );
  XNOR2XL U812 ( .A(n812), .B(B[1]), .Y(n262) );
  NOR2XL U813 ( .A(n1027), .B(n1156), .Y(n304) );
  CMPR32X1 U814 ( .A(n249), .B(n250), .C(n251), .CO(n300), .S(n297) );
  XNOR2XL U815 ( .A(n484), .B(B[4]), .Y(n277) );
  OAI22XL U816 ( .A0(n801), .A1(n277), .B0(n253), .B1(n1032), .Y(n265) );
  INVXL U817 ( .A(n812), .Y(n371) );
  CMPR32X1 U818 ( .A(n257), .B(n256), .C(n255), .CO(n249), .S(n258) );
  XNOR2XL U819 ( .A(n438), .B(B[2]), .Y(n279) );
  XNOR2XL U820 ( .A(n812), .B(B[0]), .Y(n263) );
  ADDHXL U821 ( .A(n265), .B(n264), .CO(n259), .S(n285) );
  OR2X2 U822 ( .A(n295), .B(n294), .Y(n1168) );
  NAND2XL U823 ( .A(n1164), .B(n1168), .Y(n299) );
  XNOR2XL U824 ( .A(n484), .B(B[1]), .Y(n266) );
  XNOR2XL U825 ( .A(n484), .B(B[2]), .Y(n270) );
  OAI21XL U826 ( .A0(n1179), .A1(n1185), .B0(n1180), .Y(n1177) );
  OAI22X1 U827 ( .A0(n801), .A1(n270), .B0(n278), .B1(n1032), .Y(n282) );
  XNOR2XL U828 ( .A(n438), .B(B[0]), .Y(n271) );
  XNOR2XL U829 ( .A(n438), .B(B[1]), .Y(n280) );
  OAI22X1 U830 ( .A0(n846), .A1(n271), .B0(n844), .B1(n280), .Y(n281) );
  CMPR22X1 U831 ( .A(n282), .B(n281), .CO(n283), .S(n275) );
  OAI21XL U832 ( .A0(n1174), .A1(n1171), .B0(n1172), .Y(n1189) );
  CMPR32X1 U833 ( .A(n287), .B(n286), .C(n285), .CO(n294), .S(n292) );
  CMPR32X1 U834 ( .A(n290), .B(n289), .C(n288), .CO(n291), .S(n284) );
  OR2X2 U835 ( .A(n292), .B(n291), .Y(n1188) );
  NAND2XL U836 ( .A(n295), .B(n294), .Y(n1167) );
  INVXL U837 ( .A(n1167), .Y(n1162) );
  XNOR2X1 U838 ( .A(n812), .B(B[6]), .Y(n323) );
  OAI22XL U839 ( .A0(n306), .A1(n323), .B0(n853), .B1(n305), .Y(n971) );
  XNOR2XL U840 ( .A(n803), .B(B[2]), .Y(n314) );
  OAI22XL U841 ( .A0(n1060), .A1(n314), .B0(n1061), .B1(n307), .Y(n970) );
  CMPR22X1 U842 ( .A(n309), .B(n308), .CO(n979), .S(n969) );
  CMPR22X1 U843 ( .A(n311), .B(n310), .CO(n340), .S(n336) );
  ADDFHX1 U844 ( .A(n321), .B(n320), .CI(n319), .CO(n983), .S(n339) );
  OAI22XL U845 ( .A0(n861), .A1(n322), .B0(n859), .B1(n327), .Y(n334) );
  OAI22XL U846 ( .A0(n861), .A1(n327), .B0(n859), .B1(n326), .Y(n968) );
  OAI22XL U847 ( .A0(n1083), .A1(n329), .B0(n1081), .B1(n328), .Y(n967) );
  ADDFHX1 U848 ( .A(n340), .B(n339), .CI(n338), .CO(n991), .S(n341) );
  CMPR32X1 U849 ( .A(n343), .B(n342), .C(n341), .CO(n349), .S(n348) );
  CMPR32X1 U850 ( .A(n346), .B(n345), .C(n344), .CO(n347), .S(n303) );
  INVXL U851 ( .A(n1019), .Y(n351) );
  NAND2XL U852 ( .A(n352), .B(n1033), .Y(n355) );
  NOR2XL U853 ( .A(n362), .B(n355), .Y(n357) );
  NAND2XL U854 ( .A(n429), .B(n357), .Y(n359) );
  AOI21XL U855 ( .A0(n353), .A1(n1033), .B0(n1038), .Y(n354) );
  OAI21XL U856 ( .A0(n363), .A1(n355), .B0(n354), .Y(n356) );
  AOI21XL U857 ( .A0(n470), .A1(n357), .B0(n356), .Y(n358) );
  OAI21XL U858 ( .A0(n1201), .A1(n359), .B0(n358), .Y(n361) );
  NOR2XL U859 ( .A(n362), .B(n1216), .Y(n365) );
  NAND2XL U860 ( .A(n429), .B(n365), .Y(n367) );
  OAI21XL U861 ( .A0(n363), .A1(n1216), .B0(n1217), .Y(n364) );
  AOI21XL U862 ( .A0(n470), .A1(n365), .B0(n364), .Y(n366) );
  OAI21XL U863 ( .A0(n1201), .A1(n367), .B0(n366), .Y(n368) );
  BUFX3 U864 ( .A(B[26]), .Y(n1146) );
  XNOR2X1 U865 ( .A(n812), .B(n1146), .Y(n372) );
  OAI22XL U866 ( .A0(n1060), .A1(n406), .B0(n1061), .B1(n381), .Y(n386) );
  XNOR2X1 U867 ( .A(n815), .B(n1129), .Y(n382) );
  INVXL U868 ( .A(n396), .Y(n385) );
  OAI22XL U869 ( .A0(n1108), .A1(n380), .B0(n1081), .B1(n394), .Y(n399) );
  XNOR2X1 U870 ( .A(n815), .B(B[24]), .Y(n408) );
  XNOR2X1 U871 ( .A(n1100), .B(B[18]), .Y(n410) );
  XNOR2X1 U872 ( .A(n1062), .B(B[20]), .Y(n407) );
  CMPR32X1 U873 ( .A(n387), .B(n386), .C(n385), .CO(n403), .S(n422) );
  CMPR32X1 U874 ( .A(n390), .B(n389), .C(n388), .CO(n426), .S(n421) );
  OAI22X1 U875 ( .A0(n1060), .A1(n393), .B0(n1061), .B1(n1058), .Y(n1077) );
  CMPR32X1 U876 ( .A(n397), .B(n396), .C(n395), .CO(n1069), .S(n402) );
  CMPR32X1 U877 ( .A(n400), .B(n399), .C(n398), .CO(n1068), .S(n401) );
  CMPR32X1 U878 ( .A(n403), .B(n402), .C(n401), .CO(n1054), .S(n425) );
  NOR2XL U879 ( .A(n405), .B(n404), .Y(mult_x_1_n162) );
  NAND2XL U880 ( .A(n405), .B(n404), .Y(mult_x_1_n163) );
  XNOR2X1 U881 ( .A(n1062), .B(B[19]), .Y(n450) );
  OAI22XL U882 ( .A0(n1108), .A1(n450), .B0(n1081), .B1(n407), .Y(n446) );
  INVXL U883 ( .A(n416), .Y(n444) );
  XNOR2X1 U884 ( .A(n6), .B(n805), .Y(n436) );
  OAI22XL U885 ( .A0(n1150), .A1(n436), .B0(n1148), .B1(n409), .Y(n443) );
  OAI22XL U886 ( .A0(n1133), .A1(n447), .B0(n1134), .B1(n410), .Y(n442) );
  CMPR32X1 U887 ( .A(n414), .B(n413), .C(n412), .CO(n423), .S(n464) );
  CMPR32X1 U888 ( .A(n417), .B(n416), .C(n415), .CO(n388), .S(n463) );
  CMPR32X1 U889 ( .A(n426), .B(n425), .C(n424), .CO(n405), .S(n427) );
  NOR2XL U890 ( .A(n428), .B(n427), .Y(mult_x_1_n173) );
  NAND2XL U891 ( .A(n428), .B(n427), .Y(mult_x_1_n174) );
  NAND2XL U892 ( .A(n429), .B(n471), .Y(n432) );
  XNOR2X2 U893 ( .A(n435), .B(n434), .Y(PRODUCT[32]) );
  XNOR2X1 U894 ( .A(n6), .B(B[14]), .Y(n454) );
  OAI22XL U895 ( .A0(n1150), .A1(n454), .B0(n1148), .B1(n436), .Y(n458) );
  INVXL U896 ( .A(n439), .Y(n440) );
  CMPR32X1 U897 ( .A(n443), .B(n442), .C(n441), .CO(n418), .S(n477) );
  CMPR32X1 U898 ( .A(n446), .B(n445), .C(n444), .CO(n419), .S(n476) );
  XNOR2X1 U899 ( .A(n812), .B(B[24]), .Y(n452) );
  OAI22XL U900 ( .A0(n1112), .A1(n479), .B0(n1134), .B1(n447), .Y(n460) );
  OAI22XL U901 ( .A0(n861), .A1(n453), .B0(n859), .B1(n448), .Y(n459) );
  OAI22XL U902 ( .A0(n1060), .A1(n455), .B0(n1061), .B1(n449), .Y(n488) );
  XNOR2X1 U903 ( .A(n1062), .B(B[18]), .Y(n451) );
  OAI22XL U904 ( .A0(n1108), .A1(n451), .B0(n1081), .B1(n450), .Y(n487) );
  XNOR2X1 U905 ( .A(n803), .B(B[19]), .Y(n482) );
  ADDFHX1 U906 ( .A(n458), .B(n457), .CI(n456), .CO(n478), .S(n512) );
  CMPR32X1 U907 ( .A(n461), .B(n460), .C(n459), .CO(n499), .S(n511) );
  NOR2XL U908 ( .A(n469), .B(n468), .Y(mult_x_1_n184) );
  NAND2XL U909 ( .A(n469), .B(n468), .Y(mult_x_1_n185) );
  OAI21XL U910 ( .A0(n1201), .A1(n1035), .B0(n218), .Y(n472) );
  CMPR32X1 U911 ( .A(n478), .B(n477), .C(n476), .CO(n475), .S(n510) );
  XNOR2X1 U912 ( .A(n1100), .B(n805), .Y(n481) );
  XNOR2X1 U913 ( .A(n815), .B(B[20]), .Y(n527) );
  OAI22X1 U914 ( .A0(n861), .A1(n527), .B0(n859), .B1(n480), .Y(n516) );
  XNOR2X1 U915 ( .A(n1100), .B(B[14]), .Y(n521) );
  OAI22XL U916 ( .A0(n1112), .A1(n521), .B0(n1134), .B1(n481), .Y(n517) );
  OAI22X1 U917 ( .A0(n1060), .A1(n518), .B0(n1061), .B1(n482), .Y(n530) );
  INVXL U918 ( .A(n514), .Y(n485) );
  CMPR32X1 U919 ( .A(n488), .B(n487), .C(n486), .CO(n498), .S(n535) );
  XNOR2X1 U920 ( .A(n1062), .B(B[16]), .Y(n526) );
  XNOR2X1 U921 ( .A(n812), .B(B[22]), .Y(n525) );
  OAI22XL U922 ( .A0(n855), .A1(n525), .B0(n853), .B1(n490), .Y(n531) );
  CMPR32X1 U923 ( .A(n493), .B(n492), .C(n491), .CO(n486), .S(n550) );
  NOR2XL U924 ( .A(n501), .B(n500), .Y(mult_x_1_n191) );
  NAND2XL U925 ( .A(n501), .B(n500), .Y(mult_x_1_n192) );
  INVXL U926 ( .A(n1224), .Y(n543) );
  NAND2XL U927 ( .A(n539), .B(n543), .Y(n504) );
  INVXL U928 ( .A(n1225), .Y(n502) );
  AOI21XL U929 ( .A0(n540), .A1(n543), .B0(n502), .Y(n503) );
  OAI21XL U930 ( .A0(n1201), .A1(n504), .B0(n503), .Y(n507) );
  INVXL U931 ( .A(n1222), .Y(n505) );
  XNOR2X2 U932 ( .A(n507), .B(n506), .Y(PRODUCT[30]) );
  CMPR32X1 U933 ( .A(n513), .B(n512), .C(n511), .CO(n497), .S(n548) );
  XNOR2X1 U934 ( .A(n517), .B(n516), .Y(n559) );
  XNOR2X1 U935 ( .A(A[13]), .B(B[13]), .Y(n557) );
  XNOR2X1 U936 ( .A(n812), .B(B[21]), .Y(n561) );
  XNOR2X1 U937 ( .A(n1062), .B(n805), .Y(n562) );
  OAI22XL U938 ( .A0(n1083), .A1(n562), .B0(n1081), .B1(n526), .Y(n568) );
  CMPR32X1 U939 ( .A(n533), .B(n532), .C(n531), .CO(n551), .S(n579) );
  INVXL U940 ( .A(n539), .Y(n542) );
  INVXL U941 ( .A(n540), .Y(n541) );
  OAI21XL U942 ( .A0(n1201), .A1(n542), .B0(n541), .Y(n545) );
  CMPR32X1 U943 ( .A(n551), .B(n550), .C(n549), .CO(n534), .S(n578) );
  XNOR2X1 U944 ( .A(n484), .B(B[24]), .Y(n584) );
  OAI22X1 U945 ( .A0(n838), .A1(n584), .B0(n554), .B1(n1032), .Y(n583) );
  XNOR2X1 U946 ( .A(n6), .B(B[10]), .Y(n585) );
  XNOR2X1 U947 ( .A(n803), .B(B[16]), .Y(n586) );
  OAI22X1 U948 ( .A0(n1060), .A1(n586), .B0(n1061), .B1(n555), .Y(n597) );
  XNOR2X1 U949 ( .A(A[13]), .B(B[12]), .Y(n588) );
  CMPR32X1 U950 ( .A(n560), .B(n559), .C(n558), .CO(n572), .S(n602) );
  XNOR2X1 U951 ( .A(n812), .B(B[20]), .Y(n592) );
  XNOR2X1 U952 ( .A(n1062), .B(B[14]), .Y(n593) );
  OAI22XL U953 ( .A0(n1083), .A1(n593), .B0(n1081), .B1(n562), .Y(n599) );
  CMPR32X1 U954 ( .A(n569), .B(n568), .C(n567), .CO(n581), .S(n611) );
  NOR2XL U955 ( .A(n574), .B(n573), .Y(mult_x_1_n209) );
  NAND2XL U956 ( .A(n574), .B(n573), .Y(mult_x_1_n210) );
  INVXL U957 ( .A(n1226), .Y(n575) );
  CMPR32X1 U958 ( .A(n578), .B(n577), .C(n576), .CO(n573), .S(n605) );
  CMPR32X1 U959 ( .A(n581), .B(n580), .C(n579), .CO(n570), .S(n610) );
  OAI22X1 U960 ( .A0(n801), .A1(n616), .B0(n584), .B1(n1032), .Y(n615) );
  XNOR2X1 U961 ( .A(n6), .B(B[9]), .Y(n617) );
  XNOR2X1 U962 ( .A(n803), .B(n805), .Y(n618) );
  OAI22XL U963 ( .A0(n1060), .A1(n618), .B0(n1061), .B1(n586), .Y(n629) );
  CMPR32X1 U964 ( .A(n591), .B(n590), .C(n589), .CO(n603), .S(n634) );
  XNOR2X1 U965 ( .A(n812), .B(B[19]), .Y(n624) );
  OAI22XL U966 ( .A0(n700), .A1(n626), .B0(n859), .B1(n594), .Y(n630) );
  CMPR32X1 U967 ( .A(n600), .B(n599), .C(n598), .CO(n613), .S(n648) );
  NOR2XL U968 ( .A(n605), .B(n604), .Y(mult_x_1_n220) );
  NAND2XL U969 ( .A(n605), .B(n604), .Y(mult_x_1_n221) );
  INVXL U970 ( .A(n1228), .Y(n606) );
  CMPR32X1 U971 ( .A(n613), .B(n612), .C(n611), .CO(n601), .S(n647) );
  CMPR22X1 U972 ( .A(n615), .B(n614), .CO(n622), .S(n661) );
  XNOR2X1 U973 ( .A(n803), .B(B[14]), .Y(n655) );
  XNOR2X1 U974 ( .A(A[13]), .B(B[10]), .Y(n658) );
  OAI22X1 U975 ( .A0(n1112), .A1(n658), .B0(n1134), .B1(n620), .Y(n665) );
  XNOR2X1 U976 ( .A(n812), .B(B[18]), .Y(n662) );
  XNOR2X1 U977 ( .A(n1062), .B(B[12]), .Y(n663) );
  OAI22XL U978 ( .A0(n700), .A1(n664), .B0(n859), .B1(n626), .Y(n668) );
  CMPR32X1 U979 ( .A(n635), .B(n634), .C(n633), .CO(n609), .S(n645) );
  NOR2XL U980 ( .A(n637), .B(n636), .Y(mult_x_1_n223) );
  INVXL U981 ( .A(n641), .Y(n676) );
  CMPR32X1 U982 ( .A(n647), .B(n646), .C(n645), .CO(n636), .S(n675) );
  CMPR32X1 U983 ( .A(n650), .B(n649), .C(n648), .CO(n633), .S(n683) );
  CMPR22X1 U984 ( .A(n652), .B(n651), .CO(n660), .S(n696) );
  XNOR2X1 U985 ( .A(n484), .B(B[21]), .Y(n689) );
  OAI22X1 U986 ( .A0(n801), .A1(n689), .B0(n653), .B1(n1032), .Y(n688) );
  XNOR2X1 U987 ( .A(n803), .B(B[13]), .Y(n691) );
  XNOR2X1 U988 ( .A(A[13]), .B(B[9]), .Y(n693) );
  OAI22X1 U989 ( .A0(n855), .A1(n697), .B0(n853), .B1(n662), .Y(n706) );
  OAI22X1 U990 ( .A0(n1083), .A1(n698), .B0(n1081), .B1(n663), .Y(n705) );
  ADDFHX1 U991 ( .A(n667), .B(n666), .CI(n665), .CO(n659), .S(n723) );
  NOR2XL U992 ( .A(n675), .B(n674), .Y(mult_x_1_n232) );
  NAND2XL U993 ( .A(n675), .B(n674), .Y(mult_x_1_n233) );
  NAND2XL U994 ( .A(n750), .B(n638), .Y(n678) );
  AOI21XL U995 ( .A0(n713), .A1(n638), .B0(n641), .Y(n677) );
  CMPR32X1 U996 ( .A(n683), .B(n682), .C(n681), .CO(n674), .S(n711) );
  CMPR22X1 U997 ( .A(n688), .B(n687), .CO(n695), .S(n735) );
  XNOR2X1 U998 ( .A(n484), .B(B[20]), .Y(n727) );
  OAI22X1 U999 ( .A0(n801), .A1(n727), .B0(n689), .B1(n1032), .Y(n726) );
  OAI22X1 U1000 ( .A0(n1150), .A1(n728), .B0(n1148), .B1(n690), .Y(n725) );
  XNOR2X1 U1001 ( .A(n803), .B(B[12]), .Y(n729) );
  OAI22XL U1002 ( .A0(n1060), .A1(n729), .B0(n1061), .B1(n691), .Y(n741) );
  XNOR2X1 U1003 ( .A(A[13]), .B(B[8]), .Y(n732) );
  XNOR2X1 U1004 ( .A(n812), .B(B[16]), .Y(n736) );
  OAI22X1 U1005 ( .A0(n855), .A1(n736), .B0(n853), .B1(n697), .Y(n744) );
  XNOR2X1 U1006 ( .A(n1062), .B(B[10]), .Y(n737) );
  OAI22X1 U1007 ( .A0(n1083), .A1(n737), .B0(n1081), .B1(n698), .Y(n743) );
  OAI22X1 U1008 ( .A0(n700), .A1(n738), .B0(n859), .B1(n699), .Y(n742) );
  CMPR32X1 U1009 ( .A(n709), .B(n708), .C(n707), .CO(n682), .S(n719) );
  NOR2XL U1010 ( .A(n711), .B(n710), .Y(mult_x_1_n241) );
  NAND2XL U1011 ( .A(n711), .B(n710), .Y(mult_x_1_n242) );
  NAND2XL U1012 ( .A(n750), .B(n752), .Y(n715) );
  CMPR32X1 U1013 ( .A(n721), .B(n720), .C(n719), .CO(n710), .S(n749) );
  CMPR32X1 U1014 ( .A(n724), .B(n723), .C(n722), .CO(n707), .S(n756) );
  CMPR22X1 U1015 ( .A(n726), .B(n725), .CO(n734), .S(n770) );
  XNOR2X1 U1016 ( .A(n484), .B(B[19]), .Y(n762) );
  OAI22X1 U1017 ( .A0(n801), .A1(n762), .B0(n727), .B1(n1032), .Y(n761) );
  OAI22X1 U1018 ( .A0(n1150), .A1(n763), .B0(n1148), .B1(n728), .Y(n760) );
  OAI22X1 U1019 ( .A0(n731), .A1(n766), .B0(n844), .B1(n730), .Y(n775) );
  XNOR2X1 U1020 ( .A(A[13]), .B(B[7]), .Y(n767) );
  XNOR2X1 U1021 ( .A(n805), .B(n812), .Y(n771) );
  OAI22XL U1022 ( .A0(n855), .A1(n771), .B0(n853), .B1(n736), .Y(n779) );
  XNOR2X1 U1023 ( .A(n1062), .B(B[9]), .Y(n772) );
  OAI22XL U1024 ( .A0(n1083), .A1(n772), .B0(n1081), .B1(n737), .Y(n778) );
  CMPR32X1 U1025 ( .A(n741), .B(n740), .C(n739), .CO(n733), .S(n797) );
  NOR2XL U1026 ( .A(n749), .B(n748), .Y(mult_x_1_n252) );
  NAND2XL U1027 ( .A(n749), .B(n748), .Y(mult_x_1_n253) );
  INVX1 U1028 ( .A(n1236), .Y(n752) );
  CMPR32X1 U1029 ( .A(n756), .B(n755), .C(n754), .CO(n748), .S(n784) );
  CMPR32X1 U1030 ( .A(n759), .B(n758), .C(n757), .CO(n745), .S(n795) );
  CMPR22X1 U1031 ( .A(n761), .B(n760), .CO(n769), .S(n811) );
  XNOR2XL U1032 ( .A(n6), .B(B[4]), .Y(n802) );
  OAI22X1 U1033 ( .A0(n764), .A1(n802), .B0(n1148), .B1(n763), .Y(n799) );
  XNOR2X1 U1034 ( .A(n803), .B(B[10]), .Y(n804) );
  XNOR2X1 U1035 ( .A(n812), .B(B[14]), .Y(n813) );
  OAI22XL U1036 ( .A0(n855), .A1(n813), .B0(n853), .B1(n771), .Y(n822) );
  XNOR2X1 U1037 ( .A(n1062), .B(B[8]), .Y(n814) );
  OAI22XL U1038 ( .A0(n1083), .A1(n814), .B0(n1081), .B1(n772), .Y(n821) );
  CMPR32X1 U1039 ( .A(n779), .B(n778), .C(n777), .CO(n798), .S(n831) );
  NOR2XL U1040 ( .A(n784), .B(n783), .Y(mult_x_1_n259) );
  NAND2XL U1041 ( .A(n784), .B(n783), .Y(mult_x_1_n260) );
  NAND2XL U1042 ( .A(n785), .B(n787), .Y(n789) );
  INVXL U1043 ( .A(n1238), .Y(n790) );
  CMPR32X1 U1044 ( .A(n795), .B(n794), .C(n793), .CO(n783), .S(n827) );
  CMPR32X1 U1045 ( .A(n798), .B(n797), .C(n796), .CO(n780), .S(n830) );
  CMPR22X1 U1046 ( .A(n800), .B(n799), .CO(n810), .S(n851) );
  OAI22X1 U1047 ( .A0(n1150), .A1(n839), .B0(n1148), .B1(n802), .Y(n834) );
  OAI22XL U1048 ( .A0(n1060), .A1(n841), .B0(n1061), .B1(n804), .Y(n864) );
  OAI22XL U1049 ( .A0(n846), .A1(n843), .B0(n844), .B1(n806), .Y(n863) );
  OAI22XL U1050 ( .A0(n855), .A1(n852), .B0(n853), .B1(n813), .Y(n867) );
  CMPR32X1 U1051 ( .A(n822), .B(n821), .C(n820), .CO(n833), .S(n879) );
  CMPR32X1 U1052 ( .A(n825), .B(n824), .C(n823), .CO(n794), .S(n828) );
  NOR2XL U1053 ( .A(n827), .B(n826), .Y(mult_x_1_n270) );
  NAND2XL U1054 ( .A(n827), .B(n826), .Y(mult_x_1_n271) );
  OAI22X1 U1055 ( .A0(n1150), .A1(n840), .B0(n1148), .B1(n839), .Y(n882) );
  OAI22X1 U1056 ( .A0(n1060), .A1(n842), .B0(n1061), .B1(n841), .Y(n897) );
  CMPR32X1 U1057 ( .A(n851), .B(n850), .C(n849), .CO(n870), .S(n902) );
  OAI22XL U1058 ( .A0(n855), .A1(n854), .B0(n853), .B1(n852), .Y(n900) );
  CMPR32X1 U1059 ( .A(n864), .B(n863), .C(n862), .CO(n849), .S(n912) );
  CMPR32X1 U1060 ( .A(n867), .B(n866), .C(n865), .CO(n881), .S(n911) );
  NOR2XL U1061 ( .A(n872), .B(n871), .Y(mult_x_1_n277) );
  INVXL U1062 ( .A(n1242), .Y(n873) );
  CMPR22X1 U1063 ( .A(n883), .B(n882), .CO(n890), .S(n919) );
  ADDHXL U1064 ( .A(n885), .B(n884), .CO(n918), .S(n914) );
  CMPR32X1 U1065 ( .A(n888), .B(n887), .C(n886), .CO(n917), .S(n921) );
  CMPR32X1 U1066 ( .A(n891), .B(n890), .C(n889), .CO(n903), .S(n924) );
  CMPR32X1 U1067 ( .A(n894), .B(n893), .C(n892), .CO(n934), .S(n920) );
  CMPR32X1 U1068 ( .A(n897), .B(n896), .C(n895), .CO(n889), .S(n933) );
  CMPR32X1 U1069 ( .A(n900), .B(n899), .C(n898), .CO(n913), .S(n932) );
  NOR2XL U1070 ( .A(n905), .B(n904), .Y(mult_x_1_n288) );
  NAND2XL U1071 ( .A(n905), .B(n904), .Y(mult_x_1_n289) );
  INVXL U1072 ( .A(n1244), .Y(n906) );
  NAND2XL U1073 ( .A(n906), .B(n1245), .Y(n907) );
  CMPR32X1 U1074 ( .A(n913), .B(n912), .C(n911), .CO(n901), .S(n946) );
  CMPR32X1 U1075 ( .A(n922), .B(n921), .C(n920), .CO(n938), .S(n943) );
  CMPR32X1 U1076 ( .A(n925), .B(n924), .C(n923), .CO(n909), .S(n944) );
  NOR2XL U1077 ( .A(n927), .B(n926), .Y(mult_x_1_n291) );
  NAND2XL U1078 ( .A(n927), .B(n926), .Y(mult_x_1_n292) );
  OAI21XL U1079 ( .A0(n952), .A1(n1249), .B0(n1250), .Y(n931) );
  NAND2X1 U1080 ( .A(n929), .B(n1248), .Y(n930) );
  XNOR2X2 U1081 ( .A(n931), .B(n930), .Y(PRODUCT[18]) );
  NOR2XL U1082 ( .A(mult_x_1_n302), .B(mult_x_1_n299), .Y(mult_x_1_n297) );
  NAND2XL U1083 ( .A(n951), .B(n950), .Y(mult_x_1_n300) );
  NAND2XL U1084 ( .A(n954), .B(n953), .Y(mult_x_1_n303) );
  NOR2XL U1085 ( .A(n958), .B(mult_x_1_n312), .Y(mult_x_1_n305) );
  INVXL U1086 ( .A(n958), .Y(n960) );
  NAND2XL U1087 ( .A(n960), .B(n959), .Y(mult_x_1_n78) );
  NAND2XL U1088 ( .A(n961), .B(n1254), .Y(n962) );
  XNOR2X1 U1089 ( .A(n1260), .B(n1256), .Y(PRODUCT[14]) );
  CMPR32X1 U1090 ( .A(n965), .B(n964), .C(n963), .CO(n180), .S(n999) );
  CMPR32X1 U1091 ( .A(n968), .B(n967), .C(n966), .CO(n986), .S(n981) );
  CMPR32X1 U1092 ( .A(n971), .B(n970), .C(n969), .CO(n985), .S(n992) );
  CMPR32X1 U1093 ( .A(n974), .B(n973), .C(n972), .CO(n963), .S(n984) );
  CMPR32X1 U1094 ( .A(n977), .B(n976), .C(n975), .CO(n995), .S(n997) );
  CMPR32X1 U1095 ( .A(n980), .B(n979), .C(n978), .CO(n975), .S(n989) );
  CMPR32X1 U1096 ( .A(n989), .B(n988), .C(n987), .CO(n1002), .S(n1001) );
  NAND2XL U1097 ( .A(n57), .B(n1015), .Y(n1011) );
  NOR2XL U1098 ( .A(n1011), .B(n1007), .Y(mult_x_1_n316) );
  INVXL U1099 ( .A(n1013), .Y(n1016) );
  INVXL U1100 ( .A(n1012), .Y(n1004) );
  OAI21XL U1101 ( .A0(n1010), .A1(n1007), .B0(n1008), .Y(mult_x_1_n317) );
  INVXL U1102 ( .A(n1007), .Y(n1009) );
  NAND2XL U1103 ( .A(n1009), .B(n1008), .Y(mult_x_1_n80) );
  XNOR2X1 U1104 ( .A(n1261), .B(n1257), .Y(PRODUCT[13]) );
  OAI21XL U1105 ( .A0(n1017), .A1(n1011), .B0(n1010), .Y(mult_x_1_n320) );
  NAND2XL U1106 ( .A(n57), .B(n1012), .Y(mult_x_1_n81) );
  NAND2XL U1107 ( .A(n1015), .B(n1013), .Y(n1014) );
  XOR2X1 U1108 ( .A(n1017), .B(n1014), .Y(n1276) );
  OAI21XL U1109 ( .A0(n1017), .A1(n993), .B0(n1013), .Y(mult_x_1_n327) );
  NAND2XL U1110 ( .A(n1023), .B(n1022), .Y(n1024) );
  OAI21XL U1111 ( .A0(n1160), .A1(n1156), .B0(n1157), .Y(n1031) );
  INVXL U1112 ( .A(n1027), .Y(n1029) );
  NOR2X1 U1113 ( .A(n1035), .B(n1046), .Y(n1036) );
  OAI21XL U1114 ( .A0(n1041), .A1(n1217), .B0(n1040), .Y(n1042) );
  AOI21XL U1115 ( .A0(n1044), .A1(n1043), .B0(n1042), .Y(n1045) );
  OAI21XL U1116 ( .A0(n1201), .A1(n1048), .B0(n1047), .Y(n1050) );
  XNOR2X1 U1117 ( .A(n1050), .B(n1049), .Y(PRODUCT[36]) );
  XNOR2X1 U1118 ( .A(n1053), .B(n1052), .Y(PRODUCT[37]) );
  CMPR32X1 U1119 ( .A(n1067), .B(n1066), .C(n1065), .CO(n1084), .S(n1056) );
  CMPR32X1 U1120 ( .A(n1070), .B(n1069), .C(n1068), .CO(n1073), .S(n1055) );
  CMPR32X1 U1121 ( .A(n1078), .B(n1077), .C(n1076), .CO(n1120), .S(n1075) );
  OAI22X1 U1122 ( .A0(n1083), .A1(n1082), .B0(n1081), .B1(n1106), .Y(n1115) );
  CMPR32X1 U1123 ( .A(n1086), .B(n1085), .C(n1084), .CO(n1118), .S(n1074) );
  OAI21XL U1124 ( .A0(n1201), .A1(n1096), .B0(n1095), .Y(n1099) );
  CMPR32X1 U1125 ( .A(n1104), .B(n1103), .C(n1102), .CO(n1122), .S(n1119) );
  OAI22X1 U1126 ( .A0(n1112), .A1(n1111), .B0(n1134), .B1(n1131), .Y(n1145) );
  CMPR32X1 U1127 ( .A(n1115), .B(n1114), .C(n1113), .CO(n1126), .S(n1121) );
  CMPR32X1 U1128 ( .A(n1120), .B(n1119), .C(n1118), .CO(n1125), .S(n1087) );
  CMPR32X1 U1129 ( .A(n1123), .B(n1122), .C(n1121), .CO(n1117), .S(n1124) );
  CMPR32X1 U1130 ( .A(n1128), .B(n1127), .C(n1126), .CO(n1136), .S(n1116) );
  OAI21XL U1131 ( .A0(n1138), .A1(n1206), .B0(n1207), .Y(n1194) );
  OAI21XL U1132 ( .A0(n1201), .A1(n1140), .B0(n1139), .Y(n1142) );
  CMPR32X1 U1133 ( .A(n1145), .B(n1144), .C(n1143), .CO(n1153), .S(n1135) );
  XNOR2XL U1134 ( .A(n6), .B(n1146), .Y(n1147) );
  AOI21XL U1135 ( .A0(n1169), .A1(n1168), .B0(n1162), .Y(n1166) );
  NAND2XL U1136 ( .A(n1168), .B(n1167), .Y(n1170) );
  XNOR2XL U1137 ( .A(n1190), .B(n1189), .Y(n1283) );
  OAI21XL U1138 ( .A0(n1201), .A1(n1200), .B0(n1199), .Y(n1202) );
endmodule


module FFT2048_DW02_mult_2_stage_J1_16 ( A, B, TC, CLK, PRODUCT );
  input [15:0] A;
  input [26:0] B;
  output [42:0] PRODUCT;
  input TC, CLK;
  wire   n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, mult_x_1_n335, mult_x_1_n327, mult_x_1_n320,
         mult_x_1_n317, mult_x_1_n316, mult_x_1_n313, mult_x_1_n312,
         mult_x_1_n306, mult_x_1_n305, mult_x_1_n303, mult_x_1_n302,
         mult_x_1_n300, mult_x_1_n299, mult_x_1_n297, mult_x_1_n292,
         mult_x_1_n291, mult_x_1_n289, mult_x_1_n288, mult_x_1_n278,
         mult_x_1_n277, mult_x_1_n271, mult_x_1_n270, mult_x_1_n260,
         mult_x_1_n259, mult_x_1_n253, mult_x_1_n252, mult_x_1_n242,
         mult_x_1_n241, mult_x_1_n233, mult_x_1_n232, mult_x_1_n224,
         mult_x_1_n223, mult_x_1_n221, mult_x_1_n220, mult_x_1_n210,
         mult_x_1_n209, mult_x_1_n203, mult_x_1_n202, mult_x_1_n192,
         mult_x_1_n191, mult_x_1_n185, mult_x_1_n184, mult_x_1_n174,
         mult_x_1_n173, mult_x_1_n163, mult_x_1_n162, mult_x_1_n150,
         mult_x_1_n149, mult_x_1_n135, mult_x_1_n134, mult_x_1_n126,
         mult_x_1_n125, mult_x_1_n115, mult_x_1_n114, mult_x_1_n106,
         mult_x_1_n105, mult_x_1_n81, mult_x_1_n80, mult_x_1_n78, mult_x_1_n54,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276;

  DFFHQXL clk_r_REG60_S1 ( .D(n1291), .CK(CLK), .Q(PRODUCT[11]) );
  DFFHQXL mult_x_1_clk_r_REG40_S1 ( .D(mult_x_1_n173), .CK(CLK), .Q(n1230) );
  DFFHQXL mult_x_1_clk_r_REG36_S1 ( .D(mult_x_1_n191), .CK(CLK), .Q(n1234) );
  DFFHQXL mult_x_1_clk_r_REG42_S1 ( .D(mult_x_1_n162), .CK(CLK), .Q(n1228) );
  DFFHQX4 mult_x_1_clk_r_REG54_S1 ( .D(mult_x_1_n317), .CK(CLK), .Q(n1273) );
  DFFHQX4 mult_x_1_clk_r_REG1_S1 ( .D(mult_x_1_n306), .CK(CLK), .Q(n1272) );
  DFFHQX4 mult_x_1_clk_r_REG55_S1 ( .D(mult_x_1_n316), .CK(CLK), .Q(n1269) );
  DFFHQX1 mult_x_1_clk_r_REG0_S1 ( .D(mult_x_1_n313), .CK(CLK), .Q(n1268) );
  DFFHQX4 mult_x_1_clk_r_REG5_S1 ( .D(mult_x_1_n303), .CK(CLK), .Q(n1264) );
  DFFHQX1 mult_x_1_clk_r_REG6_S1 ( .D(mult_x_1_n302), .CK(CLK), .Q(n1263) );
  DFFHQX4 mult_x_1_clk_r_REG9_S1 ( .D(mult_x_1_n299), .CK(CLK), .Q(n1261) );
  DFFHQX1 mult_x_1_clk_r_REG27_S1 ( .D(mult_x_1_n271), .CK(CLK), .Q(n1253) );
  DFFHQXL clk_r_REG58_S1 ( .D(n1290), .CK(CLK), .Q(PRODUCT[12]) );
  DFFHQX4 mult_x_1_clk_r_REG61_S1 ( .D(mult_x_1_n335), .CK(CLK), .Q(n1276) );
  DFFHQXL mult_x_1_clk_r_REG39_S1 ( .D(mult_x_1_n174), .CK(CLK), .Q(n1231) );
  DFFHQXL mult_x_1_clk_r_REG4_S1 ( .D(mult_x_1_n78), .CK(CLK), .Q(n1266) );
  DFFHQXL clk_r_REG62_S1 ( .D(n1292), .CK(CLK), .Q(PRODUCT[10]) );
  DFFHQXL mult_x_1_clk_r_REG41_S1 ( .D(mult_x_1_n163), .CK(CLK), .Q(n1229) );
  DFFHQXL mult_x_1_clk_r_REG38_S1 ( .D(mult_x_1_n184), .CK(CLK), .Q(n1232) );
  DFFHQXL clk_r_REG63_S1 ( .D(n1293), .CK(CLK), .Q(PRODUCT[9]) );
  DFFHQXL mult_x_1_clk_r_REG35_S1 ( .D(mult_x_1_n192), .CK(CLK), .Q(n1235) );
  DFFHQXL mult_x_1_clk_r_REG43_S1 ( .D(mult_x_1_n150), .CK(CLK), .Q(n1227) );
  DFFHQXL mult_x_1_clk_r_REG20_S1 ( .D(mult_x_1_n223), .CK(CLK), .Q(n1242) );
  DFFHQXL clk_r_REG64_S1 ( .D(n1294), .CK(CLK), .Q(PRODUCT[8]) );
  DFFHQXL clk_r_REG72_S1 ( .D(n1302), .CK(CLK), .Q(PRODUCT[0]) );
  DFFHQXL clk_r_REG65_S1 ( .D(n1295), .CK(CLK), .Q(PRODUCT[7]) );
  DFFHQXL clk_r_REG67_S1 ( .D(n1297), .CK(CLK), .Q(PRODUCT[5]) );
  DFFHQXL clk_r_REG71_S1 ( .D(n1301), .CK(CLK), .Q(PRODUCT[1]) );
  DFFHQXL mult_x_1_clk_r_REG57_S1 ( .D(mult_x_1_n320), .CK(CLK), .Q(n1274) );
  DFFHQXL mult_x_1_clk_r_REG24_S1 ( .D(mult_x_1_n209), .CK(CLK), .Q(n1238) );
  DFFHQXL mult_x_1_clk_r_REG56_S1 ( .D(mult_x_1_n81), .CK(CLK), .Q(n1271) );
  DFFHQX1 mult_x_1_clk_r_REG53_S1 ( .D(mult_x_1_n80), .CK(CLK), .Q(n1270) );
  DFFHQXL mult_x_1_clk_r_REG17_S1 ( .D(mult_x_1_n233), .CK(CLK), .Q(n1245) );
  DFFHQXL mult_x_1_clk_r_REG21_S1 ( .D(mult_x_1_n221), .CK(CLK), .Q(n1241) );
  DFFHQXL mult_x_1_clk_r_REG23_S1 ( .D(mult_x_1_n210), .CK(CLK), .Q(n1239) );
  DFFHQXL mult_x_1_clk_r_REG33_S1 ( .D(mult_x_1_n203), .CK(CLK), .Q(n1237) );
  DFFHQXL mult_x_1_clk_r_REG34_S1 ( .D(mult_x_1_n202), .CK(CLK), .Q(n1236) );
  DFFHQXL mult_x_1_clk_r_REG37_S1 ( .D(mult_x_1_n185), .CK(CLK), .Q(n1233) );
  DFFHQXL mult_x_1_clk_r_REG44_S1 ( .D(mult_x_1_n149), .CK(CLK), .Q(n1226) );
  DFFHQXL mult_x_1_clk_r_REG45_S1 ( .D(mult_x_1_n135), .CK(CLK), .Q(n1225) );
  DFFHQXL mult_x_1_clk_r_REG46_S1 ( .D(mult_x_1_n134), .CK(CLK), .Q(n1224) );
  DFFHQXL mult_x_1_clk_r_REG47_S1 ( .D(mult_x_1_n126), .CK(CLK), .Q(n1223) );
  DFFHQXL mult_x_1_clk_r_REG48_S1 ( .D(mult_x_1_n125), .CK(CLK), .Q(n1222) );
  DFFHQXL mult_x_1_clk_r_REG49_S1 ( .D(mult_x_1_n115), .CK(CLK), .Q(n1221) );
  DFFHQXL mult_x_1_clk_r_REG50_S1 ( .D(mult_x_1_n114), .CK(CLK), .Q(n1220) );
  DFFHQXL mult_x_1_clk_r_REG51_S1 ( .D(mult_x_1_n106), .CK(CLK), .Q(n1219) );
  DFFHQXL mult_x_1_clk_r_REG52_S1 ( .D(mult_x_1_n105), .CK(CLK), .Q(n1218) );
  DFFHQXL mult_x_1_clk_r_REG12_S1 ( .D(mult_x_1_n54), .CK(CLK), .Q(n1217) );
  DFFHQXL mult_x_1_clk_r_REG59_S1 ( .D(mult_x_1_n327), .CK(CLK), .Q(n1275) );
  DFFHQXL clk_r_REG70_S1 ( .D(n1300), .CK(CLK), .Q(PRODUCT[2]) );
  DFFHQXL clk_r_REG69_S1 ( .D(n1299), .CK(CLK), .Q(PRODUCT[3]) );
  DFFHQXL clk_r_REG68_S1 ( .D(n1298), .CK(CLK), .Q(PRODUCT[4]) );
  DFFHQXL clk_r_REG66_S1 ( .D(n1296), .CK(CLK), .Q(PRODUCT[6]) );
  DFFHQXL mult_x_1_clk_r_REG22_S1 ( .D(mult_x_1_n220), .CK(CLK), .Q(n1240) );
  DFFHQX1 mult_x_1_clk_r_REG7_S1 ( .D(mult_x_1_n297), .CK(CLK), .Q(n1260) );
  DFFHQX1 mult_x_1_clk_r_REG29_S1 ( .D(mult_x_1_n278), .CK(CLK), .Q(n1255) );
  DFFHQX1 mult_x_1_clk_r_REG16_S1 ( .D(mult_x_1_n241), .CK(CLK), .Q(n1246) );
  DFFHQXL mult_x_1_clk_r_REG19_S1 ( .D(mult_x_1_n224), .CK(CLK), .Q(n1243) );
  DFFHQX1 mult_x_1_clk_r_REG25_S1 ( .D(mult_x_1_n260), .CK(CLK), .Q(n1251) );
  DFFHQX1 mult_x_1_clk_r_REG26_S1 ( .D(mult_x_1_n259), .CK(CLK), .Q(n1250) );
  DFFHQX1 mult_x_1_clk_r_REG30_S1 ( .D(mult_x_1_n277), .CK(CLK), .Q(n1254) );
  DFFHQX1 mult_x_1_clk_r_REG8_S1 ( .D(mult_x_1_n300), .CK(CLK), .Q(n1262) );
  DFFHQX1 mult_x_1_clk_r_REG31_S1 ( .D(mult_x_1_n289), .CK(CLK), .Q(n1257) );
  DFFHQX1 mult_x_1_clk_r_REG28_S1 ( .D(mult_x_1_n270), .CK(CLK), .Q(n1252) );
  DFFHQX1 mult_x_1_clk_r_REG14_S1 ( .D(mult_x_1_n252), .CK(CLK), .Q(n1248) );
  DFFHQX1 mult_x_1_clk_r_REG18_S1 ( .D(mult_x_1_n232), .CK(CLK), .Q(n1244) );
  DFFHQX1 mult_x_1_clk_r_REG11_S1 ( .D(mult_x_1_n291), .CK(CLK), .Q(n1258) );
  DFFHQX2 mult_x_1_clk_r_REG10_S1 ( .D(mult_x_1_n292), .CK(CLK), .Q(n1259) );
  DFFHQX2 mult_x_1_clk_r_REG32_S1 ( .D(mult_x_1_n288), .CK(CLK), .Q(n1256) );
  DFFHQX1 mult_x_1_clk_r_REG13_S1 ( .D(mult_x_1_n253), .CK(CLK), .Q(n1249) );
  DFFHQX1 mult_x_1_clk_r_REG2_S1 ( .D(mult_x_1_n312), .CK(CLK), .Q(n1267) );
  DFFHQX2 mult_x_1_clk_r_REG3_S1 ( .D(mult_x_1_n305), .CK(CLK), .Q(n1265) );
  DFFHQX1 mult_x_1_clk_r_REG15_S1 ( .D(mult_x_1_n242), .CK(CLK), .Q(n1247) );
  CMPR32X1 U1 ( .A(n1072), .B(n1071), .C(n1070), .CO(n1088), .S(n496) );
  ADDFX2 U2 ( .A(n843), .B(n842), .CI(n841), .CO(n811), .S(n851) );
  CMPR32X1 U3 ( .A(n1030), .B(n1029), .C(n1028), .CO(n990), .S(n1040) );
  ADDFHX1 U4 ( .A(n560), .B(n559), .CI(n558), .CO(n562), .S(n571) );
  NAND2BX1 U5 ( .AN(n421), .B(n1058), .Y(n81) );
  ADDFX2 U6 ( .A(n621), .B(n620), .CI(n619), .CO(n633), .S(n667) );
  ADDFHX1 U7 ( .A(n944), .B(n943), .CI(n942), .CO(n950), .S(n966) );
  ADDFX2 U8 ( .A(n210), .B(n209), .CI(n208), .CO(n284), .S(n251) );
  CMPR32X1 U9 ( .A(n999), .B(n998), .C(n997), .CO(n248), .S(n1033) );
  ADDFX2 U10 ( .A(n554), .B(n553), .CI(n552), .CO(n576), .S(n610) );
  ADDFX2 U11 ( .A(n720), .B(n719), .CI(n718), .CO(n732), .S(n765) );
  ADDFX2 U12 ( .A(n787), .B(n786), .CI(n785), .CO(n800), .S(n842) );
  ADDFX2 U13 ( .A(n662), .B(n661), .CI(n660), .CO(n654), .S(n710) );
  ADDFX2 U14 ( .A(n695), .B(n694), .CI(n693), .CO(n687), .S(n743) );
  ADDFHX1 U15 ( .A(n1026), .B(n1025), .CI(n1024), .CO(n1034), .S(n418) );
  CMPR32X1 U16 ( .A(n1005), .B(n1004), .C(n1003), .CO(n1019), .S(n1026) );
  ADDFX2 U17 ( .A(n401), .B(n400), .CI(n399), .CO(n1016), .S(n410) );
  XNOR2X1 U18 ( .A(n13), .B(n452), .Y(PRODUCT[35]) );
  XNOR2X1 U19 ( .A(n570), .B(n569), .Y(PRODUCT[31]) );
  XNOR2X1 U20 ( .A(n504), .B(n503), .Y(PRODUCT[33]) );
  OAI21X1 U21 ( .A0(n443), .A1(n437), .B0(n436), .Y(n1212) );
  XNOR2X2 U22 ( .A(n605), .B(n604), .Y(PRODUCT[30]) );
  XNOR2X2 U23 ( .A(n673), .B(n672), .Y(PRODUCT[28]) );
  XNOR2X2 U24 ( .A(n640), .B(n639), .Y(PRODUCT[29]) );
  XNOR2X2 U25 ( .A(n850), .B(n849), .Y(PRODUCT[23]) );
  INVX2 U26 ( .A(n133), .Y(n1215) );
  AOI2BB1X2 U27 ( .A0N(n978), .A1N(n117), .B0(n1272), .Y(n986) );
  NAND2BX1 U28 ( .AN(n428), .B(n129), .Y(n566) );
  AND2X1 U29 ( .A(n1106), .B(n1223), .Y(n1067) );
  XOR2X1 U30 ( .A(n986), .B(n985), .Y(PRODUCT[17]) );
  XOR2XL U31 ( .A(A[2]), .B(A[3]), .Y(n142) );
  XNOR2XL U32 ( .A(n1161), .B(B[9]), .Y(n715) );
  XNOR2XL U33 ( .A(n833), .B(B[3]), .Y(n387) );
  XNOR2XL U34 ( .A(n581), .B(B[4]), .Y(n342) );
  XNOR2XL U35 ( .A(A[11]), .B(B[12]), .Y(n756) );
  XNOR2XL U36 ( .A(n833), .B(n826), .Y(n215) );
  XNOR2XL U37 ( .A(n1160), .B(n35), .Y(n535) );
  XNOR2XL U38 ( .A(A[2]), .B(A[1]), .Y(n397) );
  XNOR2XL U39 ( .A(A[12]), .B(A[11]), .Y(n144) );
  BUFX3 U40 ( .A(A[1]), .Y(n581) );
  XNOR2XL U41 ( .A(A[15]), .B(B[21]), .Y(n1096) );
  XNOR2XL U42 ( .A(A[13]), .B(n1160), .Y(n1145) );
  XOR2XL U43 ( .A(n631), .B(n22), .Y(n641) );
  ADDFX2 U44 ( .A(n270), .B(n269), .CI(n268), .CO(n974), .S(n283) );
  XOR2XL U45 ( .A(n1181), .B(n1180), .Y(n1295) );
  XOR2X1 U46 ( .A(n1175), .B(n1174), .Y(n1294) );
  NAND2XL U47 ( .A(n595), .B(n596), .Y(n30) );
  OAI21XL U48 ( .A0(n42), .A1(n741), .B0(n739), .Y(n45) );
  NAND2XL U49 ( .A(n811), .B(n812), .Y(n23) );
  OAI21XL U50 ( .A0(n811), .A1(n812), .B0(n810), .Y(n24) );
  INVX1 U51 ( .A(n1034), .Y(n54) );
  NAND2X1 U52 ( .A(n1040), .B(n1039), .Y(n1042) );
  NAND2X1 U53 ( .A(n418), .B(n417), .Y(n1052) );
  NAND2X1 U54 ( .A(n42), .B(n741), .Y(n44) );
  NAND2XL U55 ( .A(n667), .B(n668), .Y(n88) );
  ADDFHX1 U56 ( .A(n256), .B(n255), .CI(n254), .CO(n257), .S(n991) );
  INVX1 U57 ( .A(n741), .Y(n43) );
  NAND2XL U58 ( .A(n799), .B(n800), .Y(n36) );
  NAND2X1 U59 ( .A(n56), .B(n55), .Y(n268) );
  INVX1 U60 ( .A(n812), .Y(n25) );
  NOR2X1 U61 ( .A(n367), .B(n366), .Y(n1171) );
  INVXL U62 ( .A(n596), .Y(n32) );
  NAND2XL U63 ( .A(n49), .B(n48), .Y(n47) );
  INVX1 U64 ( .A(n535), .Y(n34) );
  INVX1 U65 ( .A(n50), .Y(n49) );
  OAI22X1 U66 ( .A0(n50), .A1(n875), .B0(n873), .B1(n46), .Y(n797) );
  OAI22X1 U67 ( .A0(n819), .A1(n1064), .B0(n17), .B1(n820), .Y(n120) );
  XNOR2X1 U68 ( .A(n462), .B(n1160), .Y(n463) );
  XNOR2X1 U69 ( .A(n1216), .B(n1217), .Y(PRODUCT[40]) );
  XOR2X1 U70 ( .A(n1068), .B(n1067), .Y(PRODUCT[37]) );
  XNOR2X1 U71 ( .A(n462), .B(B[13]), .Y(n265) );
  XNOR2X1 U72 ( .A(A[15]), .B(n818), .Y(n483) );
  XNOR2X1 U73 ( .A(B[20]), .B(A[3]), .Y(n751) );
  BUFX3 U74 ( .A(B[5]), .Y(n821) );
  INVX1 U75 ( .A(n566), .Y(n443) );
  NAND2XL U76 ( .A(n133), .B(n636), .Y(n116) );
  INVX1 U77 ( .A(n866), .Y(n40) );
  NAND2X1 U78 ( .A(n442), .B(n435), .Y(n437) );
  NAND2BXL U79 ( .AN(n931), .B(n426), .Y(n108) );
  INVXL U80 ( .A(n873), .Y(n48) );
  AOI21X1 U81 ( .A0(n599), .A1(n638), .B0(n600), .Y(n601) );
  INVXL U82 ( .A(n425), .Y(n132) );
  AND2X2 U83 ( .A(n738), .B(n1245), .Y(n61) );
  INVX1 U84 ( .A(n581), .Y(n6) );
  INVX1 U85 ( .A(n462), .Y(n5) );
  INVX1 U86 ( .A(n1238), .Y(n638) );
  INVX1 U87 ( .A(n1234), .Y(n568) );
  INVX1 U88 ( .A(n1222), .Y(n1106) );
  INVX1 U89 ( .A(n1226), .Y(n431) );
  NAND2X1 U90 ( .A(n98), .B(n97), .Y(n565) );
  XNOR2X1 U91 ( .A(n1063), .B(n1062), .Y(n1293) );
  OAI2BB1X1 U92 ( .A0N(n900), .A1N(n899), .B0(n118), .Y(n891) );
  NAND2X1 U93 ( .A(n45), .B(n44), .Y(n733) );
  NAND2X1 U94 ( .A(n24), .B(n23), .Y(n801) );
  INVXL U95 ( .A(n1048), .Y(n1027) );
  NAND2X1 U96 ( .A(n58), .B(n1048), .Y(n1045) );
  NAND2BX1 U97 ( .AN(n1035), .B(n54), .Y(n1048) );
  NAND2BXL U98 ( .AN(n595), .B(n32), .Y(n31) );
  NAND2XL U99 ( .A(n632), .B(n633), .Y(n20) );
  NOR2XL U100 ( .A(n977), .B(n976), .Y(mult_x_1_n291) );
  NAND2X1 U101 ( .A(n1035), .B(n1034), .Y(n1046) );
  XNOR2X1 U102 ( .A(n798), .B(n38), .Y(n810) );
  NAND2X1 U103 ( .A(n798), .B(n37), .Y(n29) );
  NAND2X1 U104 ( .A(n1179), .B(n1183), .Y(n365) );
  NAND2X1 U105 ( .A(n1017), .B(n1016), .Y(n52) );
  OR2X2 U106 ( .A(n799), .B(n800), .Y(n37) );
  NAND2X1 U107 ( .A(n367), .B(n366), .Y(n1172) );
  INVXL U108 ( .A(n363), .Y(n78) );
  ADDFHX2 U109 ( .A(n755), .B(n754), .CI(n753), .CO(n766), .S(n799) );
  XNOR2X1 U110 ( .A(n615), .B(n614), .Y(n655) );
  ADDFHX1 U111 ( .A(n797), .B(n796), .CI(n795), .CO(n815), .S(n854) );
  XNOR2X1 U112 ( .A(n833), .B(n1160), .Y(n468) );
  XNOR2X1 U113 ( .A(n823), .B(n1160), .Y(n1074) );
  OAI22X1 U114 ( .A0(n26), .A1(n866), .B0(n751), .B1(n864), .Y(n793) );
  OAI22X1 U115 ( .A0(n685), .A1(n864), .B0(n866), .B1(n41), .Y(n725) );
  OAI22X1 U116 ( .A0(n875), .A1(n721), .B0(n873), .B1(n690), .Y(n729) );
  NAND2BX1 U117 ( .AN(n751), .B(n40), .Y(n39) );
  XNOR2X1 U118 ( .A(B[11]), .B(n1078), .Y(n789) );
  OAI2BB1XL U119 ( .A0N(n528), .A1N(n133), .B0(n443), .Y(n570) );
  NOR2X1 U120 ( .A(n567), .B(n437), .Y(n427) );
  NAND3X1 U121 ( .A(n87), .B(n86), .C(n770), .Y(n85) );
  NAND3X1 U122 ( .A(n77), .B(n74), .C(n73), .Y(n72) );
  AOI21X1 U123 ( .A0(n426), .A1(n131), .B0(n125), .Y(n124) );
  NAND2X1 U124 ( .A(n429), .B(n599), .Y(n129) );
  NAND2XL U125 ( .A(n846), .B(n735), .Y(n87) );
  NAND2X1 U126 ( .A(n132), .B(n846), .Y(n10) );
  INVX1 U127 ( .A(A[3]), .Y(n27) );
  AND2X2 U128 ( .A(n771), .B(n1247), .Y(n60) );
  NAND2X1 U129 ( .A(n807), .B(n1249), .Y(n808) );
  AND2X2 U130 ( .A(n932), .B(n1255), .Y(n59) );
  NAND2X1 U131 ( .A(n531), .B(n1233), .Y(n532) );
  NAND2X1 U132 ( .A(n502), .B(n1231), .Y(n503) );
  NAND2X1 U133 ( .A(n568), .B(n1235), .Y(n569) );
  INVX1 U134 ( .A(A[3]), .Y(n35) );
  INVX1 U135 ( .A(n1228), .Y(n457) );
  NOR2X1 U136 ( .A(n1234), .B(n1232), .Y(n442) );
  XNOR2X1 U137 ( .A(A[6]), .B(A[5]), .Y(n139) );
  XOR2X1 U138 ( .A(A[10]), .B(A[11]), .Y(n136) );
  NAND2XL U139 ( .A(n572), .B(n573), .Y(n97) );
  XOR3X2 U140 ( .A(n573), .B(n571), .C(n572), .Y(n598) );
  XNOR2X1 U141 ( .A(n594), .B(n33), .Y(n606) );
  OAI2BB1X1 U142 ( .A0N(n31), .A1N(n594), .B0(n30), .Y(n572) );
  XNOR3X2 U143 ( .A(n740), .B(n43), .C(n739), .Y(n768) );
  XNOR3X2 U144 ( .A(n25), .B(n810), .C(n811), .Y(n845) );
  NAND2X1 U145 ( .A(n29), .B(n36), .Y(n773) );
  XNOR2X1 U146 ( .A(n595), .B(n596), .Y(n33) );
  NAND2XL U147 ( .A(n952), .B(n951), .Y(mult_x_1_n278) );
  OR2X2 U148 ( .A(n632), .B(n633), .Y(n21) );
  NOR2X1 U149 ( .A(n1040), .B(n1039), .Y(n1041) );
  INVX1 U150 ( .A(n414), .Y(n1056) );
  ADDFHX2 U151 ( .A(n975), .B(n974), .CI(n973), .CO(n976), .S(n983) );
  ADDFHX1 U152 ( .A(n958), .B(n957), .CI(n956), .CO(n951), .S(n969) );
  NOR2X1 U153 ( .A(n991), .B(n990), .Y(mult_x_1_n312) );
  NOR2X1 U154 ( .A(n416), .B(n415), .Y(n414) );
  OR2XL U155 ( .A(n1168), .B(n1167), .Y(n1170) );
  NAND2BXL U156 ( .AN(n731), .B(n111), .Y(n110) );
  INVXL U157 ( .A(n899), .Y(n119) );
  OAI2BB1X1 U158 ( .A0N(n53), .A1N(n1015), .B0(n52), .Y(n1022) );
  OAI2BB1XL U159 ( .A0N(n93), .A1N(n589), .B0(n92), .Y(n583) );
  ADDFHX1 U160 ( .A(n972), .B(n971), .CI(n970), .CO(n968), .S(n977) );
  ADDFHX2 U161 ( .A(n701), .B(n700), .CI(n699), .CO(n675), .S(n706) );
  ADDFHX1 U162 ( .A(n1033), .B(n1032), .CI(n1031), .CO(n1039), .S(n1037) );
  NAND2XL U163 ( .A(n967), .B(n966), .Y(n67) );
  ADDFHX2 U164 ( .A(n950), .B(n949), .CI(n948), .CO(n934), .S(n956) );
  XOR3X2 U165 ( .A(n1016), .B(n1017), .C(n1015), .Y(n1024) );
  OR2X2 U166 ( .A(n889), .B(n890), .Y(n64) );
  ADDFHX1 U167 ( .A(n410), .B(n409), .CI(n408), .CO(n417), .S(n416) );
  NAND2BXL U168 ( .AN(n1177), .B(n1178), .Y(n105) );
  NAND2X1 U169 ( .A(n78), .B(n106), .Y(n1179) );
  INVXL U170 ( .A(n732), .Y(n111) );
  XNOR2X1 U171 ( .A(n889), .B(n890), .Y(n71) );
  OAI22X2 U172 ( .A0(n586), .A1(n866), .B0(n864), .B1(n34), .Y(n553) );
  NAND2XL U173 ( .A(n191), .B(n192), .Y(n55) );
  INVXL U174 ( .A(n190), .Y(n57) );
  ADDFHX2 U175 ( .A(n830), .B(n829), .CI(n828), .CO(n843), .S(n889) );
  ADDFHX1 U176 ( .A(n407), .B(n406), .CI(n405), .CO(n1025), .S(n408) );
  OR2X2 U177 ( .A(n1017), .B(n1016), .Y(n53) );
  INVXL U178 ( .A(n362), .Y(n106) );
  XOR2X1 U179 ( .A(n69), .B(n276), .Y(n273) );
  OR2X2 U180 ( .A(n358), .B(n357), .Y(n356) );
  OAI22XL U181 ( .A0(n551), .A1(n1077), .B0(n1076), .B1(n91), .Y(n591) );
  OAI22X1 U182 ( .A0(n858), .A1(n859), .B0(n1064), .B1(n17), .Y(n905) );
  OAI22X1 U183 ( .A0(n721), .A1(n873), .B0(n875), .B1(n46), .Y(n763) );
  OAI21XL U184 ( .A0(n864), .A1(n41), .B0(n39), .Y(n759) );
  OAI22X1 U185 ( .A0(n242), .A1(n1064), .B0(n859), .B1(n51), .Y(n374) );
  XNOR2X1 U186 ( .A(n1114), .B(n1113), .Y(PRODUCT[38]) );
  XNOR2X1 U187 ( .A(n1156), .B(n1155), .Y(PRODUCT[39]) );
  XNOR2X1 U188 ( .A(n441), .B(n440), .Y(PRODUCT[36]) );
  OR2X2 U189 ( .A(n339), .B(n338), .Y(n337) );
  NOR2BX1 U190 ( .AN(n451), .B(n14), .Y(n13) );
  INVXL U191 ( .A(n1212), .Y(n438) );
  AND2XL U192 ( .A(n1201), .B(n1200), .Y(n1301) );
  OR2XL U193 ( .A(n1199), .B(n1198), .Y(n1201) );
  OAI22XL U194 ( .A0(n1165), .A1(n170), .B0(n1163), .B1(n275), .Y(n276) );
  OAI22XL U195 ( .A0(n380), .A1(n379), .B0(n1077), .B1(n378), .Y(n384) );
  NAND3X2 U196 ( .A(n10), .B(n9), .C(n11), .Y(n133) );
  AND2XL U197 ( .A(n1205), .B(n1207), .Y(n1211) );
  INVXL U198 ( .A(n846), .Y(n736) );
  NAND2X1 U199 ( .A(n142), .B(n397), .Y(n391) );
  NOR2BXL U200 ( .AN(B[0]), .B(n1127), .Y(n386) );
  NAND2X1 U201 ( .A(n135), .B(n341), .Y(n371) );
  NOR2X1 U202 ( .A(n130), .B(n423), .Y(n11) );
  NAND2X1 U203 ( .A(n15), .B(n1241), .Y(n599) );
  NAND2X1 U204 ( .A(n131), .B(n1259), .Y(n211) );
  NAND2BX1 U205 ( .AN(n1240), .B(n16), .Y(n15) );
  AND2X2 U206 ( .A(n431), .B(n1227), .Y(n452) );
  NAND2X1 U207 ( .A(n138), .B(n139), .Y(n791) );
  NAND2X1 U208 ( .A(n136), .B(n137), .Y(n1126) );
  NAND2X1 U209 ( .A(n143), .B(n144), .Y(n1147) );
  NAND2X1 U210 ( .A(n149), .B(n150), .Y(n484) );
  NAND2X1 U211 ( .A(n704), .B(n1243), .Y(n705) );
  NAND2XL U212 ( .A(n954), .B(n1257), .Y(n955) );
  INVXL U213 ( .A(n735), .Y(n769) );
  NAND2X1 U214 ( .A(n429), .B(n636), .Y(n567) );
  INVXL U215 ( .A(n1247), .Y(n75) );
  NOR2X1 U216 ( .A(n1238), .B(n1236), .Y(n429) );
  INVX1 U217 ( .A(n1243), .Y(n16) );
  INVX1 U218 ( .A(n1224), .Y(n1104) );
  INVX1 U219 ( .A(n1258), .Y(n131) );
  INVXL U220 ( .A(n1267), .Y(n995) );
  XNOR2X1 U221 ( .A(A[10]), .B(A[9]), .Y(n137) );
  INVX1 U222 ( .A(n1250), .Y(n848) );
  INVX1 U223 ( .A(A[0]), .Y(n747) );
  OAI21X4 U224 ( .A0(n978), .A1(n113), .B0(n7), .Y(n426) );
  NOR2X4 U225 ( .A(n12), .B(n8), .Y(n7) );
  AND2X2 U226 ( .A(n1260), .B(n1272), .Y(n8) );
  AOI21X4 U227 ( .A0(n1269), .A1(n1276), .B0(n1273), .Y(n978) );
  NOR2X1 U228 ( .A(n1250), .B(n1248), .Y(n735) );
  NAND2X1 U229 ( .A(n96), .B(n426), .Y(n9) );
  XOR2X2 U230 ( .A(n1215), .B(n705), .Y(PRODUCT[27]) );
  OAI21X1 U231 ( .A0(n1261), .A1(n1264), .B0(n1262), .Y(n12) );
  INVX1 U232 ( .A(n567), .Y(n528) );
  NOR3BX1 U233 ( .AN(n450), .B(n567), .C(n1215), .Y(n14) );
  OAI2BB1X1 U234 ( .A0N(n110), .A1N(n730), .B0(n109), .Y(n707) );
  BUFX3 U235 ( .A(B[19]), .Y(n818) );
  XOR2X1 U236 ( .A(n818), .B(n6), .Y(n17) );
  NOR2X1 U237 ( .A(n597), .B(n598), .Y(mult_x_1_n191) );
  NAND2XL U238 ( .A(n590), .B(n18), .Y(n92) );
  INVXL U239 ( .A(n94), .Y(n18) );
  XNOR2X2 U240 ( .A(n590), .B(n94), .Y(n95) );
  AOI2BB1X4 U241 ( .A0N(n587), .A1N(n1098), .B0(n19), .Y(n94) );
  NOR2X1 U242 ( .A(n547), .B(n1127), .Y(n19) );
  OAI2BB1X2 U243 ( .A0N(n21), .A1N(n631), .B0(n20), .Y(n607) );
  XOR2X1 U244 ( .A(n632), .B(n633), .Y(n22) );
  OAI22X1 U245 ( .A0(n28), .A1(n866), .B0(n864), .B1(n26), .Y(n836) );
  XOR2X2 U246 ( .A(n818), .B(n27), .Y(n26) );
  OAI22X1 U247 ( .A0(n121), .A1(n866), .B0(n864), .B1(n28), .Y(n883) );
  XNOR2X1 U248 ( .A(n783), .B(A[3]), .Y(n28) );
  NOR2X1 U249 ( .A(n767), .B(n768), .Y(mult_x_1_n232) );
  NAND2X1 U250 ( .A(n597), .B(n598), .Y(mult_x_1_n192) );
  XNOR2X1 U251 ( .A(n799), .B(n800), .Y(n38) );
  XNOR2X1 U252 ( .A(B[21]), .B(A[3]), .Y(n41) );
  BUFX2 U253 ( .A(n740), .Y(n42) );
  XOR2X1 U254 ( .A(n783), .B(n5), .Y(n46) );
  OAI21XL U255 ( .A0(n831), .A1(n875), .B0(n47), .Y(n840) );
  XNOR2X1 U256 ( .A(n825), .B(n462), .Y(n50) );
  OAI22X1 U257 ( .A0(n377), .A1(n859), .B0(n1064), .B1(n51), .Y(n385) );
  XNOR2X1 U258 ( .A(n788), .B(n581), .Y(n51) );
  OAI21XL U259 ( .A0(n191), .A1(n192), .B0(n190), .Y(n56) );
  XNOR3X2 U260 ( .A(n192), .B(n191), .C(n57), .Y(n253) );
  XOR3X2 U261 ( .A(n285), .B(n284), .C(n283), .Y(n988) );
  XNOR2X1 U262 ( .A(B[14]), .B(A[3]), .Y(n175) );
  XNOR2XL U263 ( .A(A[11]), .B(B[2]), .Y(n225) );
  NAND2X1 U264 ( .A(n133), .B(n704), .Y(n66) );
  XNOR2X1 U265 ( .A(n888), .B(n71), .Y(n898) );
  XNOR2X1 U266 ( .A(n581), .B(B[20]), .Y(n819) );
  INVX1 U267 ( .A(n1265), .Y(n117) );
  BUFX4 U268 ( .A(B[7]), .Y(n826) );
  XNOR2XL U269 ( .A(n833), .B(B[16]), .Y(n757) );
  XNOR2XL U270 ( .A(A[3]), .B(B[16]), .Y(n865) );
  XNOR2XL U271 ( .A(n833), .B(B[23]), .Y(n544) );
  NAND2X1 U272 ( .A(n1265), .B(n1260), .Y(n113) );
  NAND2XL U273 ( .A(n1104), .B(n1225), .Y(n440) );
  NAND2XL U274 ( .A(n427), .B(n1104), .Y(n1066) );
  NAND2XL U275 ( .A(n457), .B(n1229), .Y(n458) );
  INVXL U276 ( .A(n1261), .Y(n979) );
  XNOR2XL U277 ( .A(n462), .B(B[20]), .Y(n690) );
  XNOR2XL U278 ( .A(n833), .B(n783), .Y(n692) );
  XNOR2X1 U279 ( .A(n462), .B(n818), .Y(n721) );
  XNOR2X1 U280 ( .A(n833), .B(n825), .Y(n723) );
  XNOR2X1 U281 ( .A(n823), .B(n788), .Y(n863) );
  XNOR2XL U282 ( .A(n833), .B(B[12]), .Y(n880) );
  XNOR2XL U283 ( .A(n833), .B(B[11]), .Y(n267) );
  XNOR2XL U284 ( .A(n833), .B(n788), .Y(n147) );
  OAI21XL U285 ( .A0(n103), .A1(n161), .B0(n160), .Y(n100) );
  XNOR2XL U286 ( .A(n462), .B(B[9]), .Y(n204) );
  XNOR2XL U287 ( .A(n1078), .B(B[3]), .Y(n218) );
  OAI22XL U288 ( .A0(n1135), .A1(n165), .B0(n1148), .B1(n164), .Y(n222) );
  OAI22XL U289 ( .A0(n859), .A1(n224), .B0(n163), .B1(n1064), .Y(n223) );
  NAND2BXL U290 ( .AN(B[0]), .B(A[13]), .Y(n164) );
  XNOR2X1 U291 ( .A(n462), .B(B[21]), .Y(n657) );
  XNOR2XL U292 ( .A(n833), .B(n818), .Y(n659) );
  XNOR2XL U293 ( .A(n1078), .B(B[16]), .Y(n623) );
  XNOR2X1 U294 ( .A(A[3]), .B(B[24]), .Y(n617) );
  XNOR2XL U295 ( .A(n462), .B(B[25]), .Y(n542) );
  XNOR2X1 U296 ( .A(n1118), .B(n825), .Y(n543) );
  XNOR2X1 U297 ( .A(n823), .B(B[21]), .Y(n545) );
  XNOR2XL U298 ( .A(n1078), .B(n818), .Y(n546) );
  XNOR2XL U299 ( .A(n823), .B(B[25]), .Y(n485) );
  XNOR2X1 U300 ( .A(n823), .B(B[24]), .Y(n472) );
  XNOR2X1 U301 ( .A(n1118), .B(B[20]), .Y(n470) );
  XNOR2XL U302 ( .A(n833), .B(B[25]), .Y(n473) );
  XNOR2XL U303 ( .A(n1078), .B(B[20]), .Y(n506) );
  XNOR2XL U304 ( .A(B[6]), .B(n581), .Y(n308) );
  NAND2XL U305 ( .A(n1112), .B(n1221), .Y(n1113) );
  INVXL U306 ( .A(n1220), .Y(n1112) );
  OAI22XL U307 ( .A0(n1135), .A1(n867), .B0(n1148), .B1(n827), .Y(n882) );
  OAI22XL U308 ( .A0(n1135), .A1(n176), .B0(n1148), .B1(n264), .Y(n277) );
  XNOR2XL U309 ( .A(n1118), .B(B[16]), .Y(n577) );
  ADDFX2 U310 ( .A(n627), .B(n626), .CI(n625), .CO(n619), .S(n678) );
  OAI2BB1XL U311 ( .A0N(n747), .A1N(n859), .B0(n582), .Y(n625) );
  OAI22XL U312 ( .A0(n1165), .A1(n613), .B0(n1163), .B1(n580), .Y(n626) );
  OAI22XL U313 ( .A0(n616), .A1(n1076), .B0(n1077), .B1(n91), .Y(n627) );
  XNOR2XL U314 ( .A(n1118), .B(B[22]), .Y(n1080) );
  XNOR2X1 U315 ( .A(n1118), .B(B[21]), .Y(n482) );
  XNOR2XL U316 ( .A(n1078), .B(B[23]), .Y(n486) );
  XNOR2X1 U317 ( .A(n1078), .B(B[24]), .Y(n1079) );
  XNOR2XL U318 ( .A(n823), .B(B[22]), .Y(n510) );
  XNOR2XL U319 ( .A(n1078), .B(B[22]), .Y(n471) );
  NAND2XL U320 ( .A(n1207), .B(n1219), .Y(n1155) );
  NAND2XL U321 ( .A(n427), .B(n1205), .Y(n1154) );
  XNOR2XL U322 ( .A(n1118), .B(B[25]), .Y(n1134) );
  XNOR2X1 U323 ( .A(n1118), .B(B[24]), .Y(n1119) );
  NOR2BXL U324 ( .AN(B[0]), .B(n341), .Y(n355) );
  OAI22XL U325 ( .A0(n866), .A1(n345), .B0(n397), .B1(n344), .Y(n353) );
  OAI22XL U326 ( .A0(n859), .A1(n343), .B0(n342), .B1(n1064), .Y(n354) );
  OAI22XL U327 ( .A0(n371), .A1(n327), .B0(n873), .B1(n326), .Y(n351) );
  OAI22XL U328 ( .A0(n866), .A1(n344), .B0(n864), .B1(n325), .Y(n352) );
  NOR2X1 U329 ( .A(n1258), .B(n1256), .Y(n928) );
  INVXL U330 ( .A(n1239), .Y(n600) );
  NAND2XL U331 ( .A(n636), .B(n638), .Y(n602) );
  NAND2XL U332 ( .A(n426), .B(n803), .Y(n126) );
  AOI21XL U333 ( .A0(n846), .A1(n848), .B0(n804), .Y(n805) );
  INVXL U334 ( .A(n1251), .Y(n804) );
  AOI21XL U335 ( .A0(n566), .A1(n568), .B0(n529), .Y(n128) );
  XNOR2XL U336 ( .A(A[3]), .B(B[9]), .Y(n396) );
  XNOR2XL U337 ( .A(n833), .B(n821), .Y(n392) );
  NAND2BXL U338 ( .AN(B[0]), .B(n823), .Y(n290) );
  XOR2X1 U339 ( .A(n996), .B(n978), .Y(PRODUCT[15]) );
  XNOR2X1 U340 ( .A(n1274), .B(n1270), .Y(PRODUCT[14]) );
  XOR2X1 U341 ( .A(n127), .B(n1266), .Y(PRODUCT[16]) );
  AOI2BB1X2 U342 ( .A0N(n978), .A1N(n1267), .B0(n989), .Y(n127) );
  AND2X2 U343 ( .A(n123), .B(n894), .Y(n122) );
  XOR2X2 U344 ( .A(n85), .B(n60), .Y(PRODUCT[25]) );
  NAND2X1 U345 ( .A(n66), .B(n1243), .Y(n673) );
  XNOR2X1 U346 ( .A(A[13]), .B(n788), .Y(n752) );
  XNOR2XL U347 ( .A(n823), .B(B[11]), .Y(n862) );
  XNOR2XL U348 ( .A(n823), .B(B[8]), .Y(n173) );
  XNOR2XL U349 ( .A(n462), .B(B[11]), .Y(n148) );
  NAND2BXL U350 ( .AN(B[0]), .B(n1161), .Y(n151) );
  XNOR2X1 U351 ( .A(A[3]), .B(B[13]), .Y(n178) );
  XNOR2XL U352 ( .A(n833), .B(B[9]), .Y(n182) );
  XOR2X1 U353 ( .A(B[14]), .B(n6), .Y(n152) );
  XNOR2XL U354 ( .A(n1118), .B(B[2]), .Y(n158) );
  XNOR2X1 U355 ( .A(A[3]), .B(n788), .Y(n227) );
  XNOR2XL U356 ( .A(n462), .B(B[8]), .Y(n228) );
  XNOR2XL U357 ( .A(n823), .B(B[4]), .Y(n241) );
  NOR2BXL U358 ( .AN(B[0]), .B(n1148), .Y(n247) );
  OAI22XL U359 ( .A0(n1098), .A1(n394), .B0(n1127), .B1(n225), .Y(n245) );
  XNOR2XL U360 ( .A(n833), .B(B[22]), .Y(n549) );
  NAND2BXL U361 ( .AN(n590), .B(n94), .Y(n93) );
  XNOR2XL U362 ( .A(n823), .B(B[20]), .Y(n551) );
  XNOR2XL U363 ( .A(n1118), .B(n818), .Y(n474) );
  XNOR2XL U364 ( .A(n823), .B(B[3]), .Y(n372) );
  NAND2BXL U365 ( .AN(B[0]), .B(A[11]), .Y(n243) );
  XNOR2XL U366 ( .A(n462), .B(B[4]), .Y(n287) );
  NAND2BXL U367 ( .AN(B[0]), .B(n833), .Y(n288) );
  XOR2X1 U368 ( .A(n826), .B(n6), .Y(n82) );
  NOR2XL U369 ( .A(n1151), .B(n1220), .Y(n1205) );
  INVXL U370 ( .A(n1218), .Y(n1207) );
  OAI22XL U371 ( .A0(n1135), .A1(n686), .B0(n1148), .B1(n653), .Y(n693) );
  OAI22X1 U372 ( .A0(n1076), .A1(n684), .B0(n1077), .B1(n651), .Y(n695) );
  OAI22XL U373 ( .A0(n1135), .A1(n717), .B0(n1148), .B1(n686), .Y(n724) );
  ADDFX2 U374 ( .A(n729), .B(n728), .CI(n727), .CO(n744), .S(n775) );
  OAI22X1 U375 ( .A0(n1098), .A1(n722), .B0(n1127), .B1(n691), .Y(n728) );
  OAI22XL U376 ( .A0(n881), .A1(n790), .B0(n879), .B1(n757), .Y(n795) );
  OAI22XL U377 ( .A0(n1135), .A1(n827), .B0(n1148), .B1(n784), .Y(n835) );
  OAI22XL U378 ( .A0(n881), .A1(n878), .B0(n879), .B1(n834), .Y(n885) );
  ADDFX2 U379 ( .A(n913), .B(n912), .CI(n911), .CO(n925), .S(n949) );
  OAI22XL U380 ( .A0(n881), .A1(n880), .B0(n879), .B1(n878), .Y(n920) );
  OAI22XL U381 ( .A0(n875), .A1(n874), .B0(n873), .B1(n872), .Y(n922) );
  OAI22XL U382 ( .A0(n1135), .A1(n264), .B0(n1148), .B1(n868), .Y(n908) );
  OAI22X1 U383 ( .A0(n866), .A1(n263), .B0(n864), .B1(n865), .Y(n909) );
  OAI22XL U384 ( .A0(n881), .A1(n147), .B0(n879), .B1(n267), .Y(n259) );
  OAI22X1 U385 ( .A0(n174), .A1(n1077), .B0(n380), .B1(n159), .Y(n103) );
  OAI22XL U386 ( .A0(n1165), .A1(n157), .B0(n1163), .B1(n156), .Y(n161) );
  CMPR32X1 U387 ( .A(n207), .B(n206), .C(n205), .CO(n214), .S(n232) );
  CMPR32X1 U388 ( .A(n221), .B(n220), .C(n219), .CO(n212), .S(n249) );
  OAI22XL U389 ( .A0(n881), .A1(n215), .B0(n879), .B1(n183), .Y(n220) );
  OAI22X1 U390 ( .A0(n875), .A1(n588), .B0(n873), .B1(n548), .Y(n590) );
  ADDFX2 U391 ( .A(n593), .B(n592), .CI(n591), .CO(n611), .S(n644) );
  OAI22X1 U392 ( .A0(n1165), .A1(n580), .B0(n1163), .B1(n550), .Y(n592) );
  OAI22XL U393 ( .A0(n881), .A1(n578), .B0(n879), .B1(n549), .Y(n593) );
  OAI22XL U394 ( .A0(n820), .A1(n649), .B0(n612), .B1(n1064), .Y(n648) );
  OAI22XL U395 ( .A0(n1135), .A1(n653), .B0(n1148), .B1(n618), .Y(n660) );
  OAI22XL U396 ( .A0(n1076), .A1(n651), .B0(n1077), .B1(n616), .Y(n662) );
  ADDFX2 U397 ( .A(n665), .B(n664), .CI(n663), .CO(n679), .S(n709) );
  OAI22XL U398 ( .A0(n1126), .A1(n658), .B0(n1127), .B1(n623), .Y(n664) );
  OAI22XL U399 ( .A0(n875), .A1(n657), .B0(n873), .B1(n622), .Y(n665) );
  XNOR2XL U400 ( .A(n823), .B(B[23]), .Y(n505) );
  OAI22XL U401 ( .A0(n1076), .A1(n545), .B0(n1077), .B1(n510), .Y(n536) );
  OAI22XL U402 ( .A0(n1165), .A1(n534), .B0(n1163), .B1(n508), .Y(n538) );
  OAI22XL U403 ( .A0(n1098), .A1(n546), .B0(n1127), .B1(n506), .Y(n541) );
  OAI22XL U404 ( .A0(n881), .A1(n544), .B0(n879), .B1(n507), .Y(n540) );
  XNOR2X1 U405 ( .A(n1078), .B(B[21]), .Y(n475) );
  OAI2BB1XL U406 ( .A0N(n873), .A1N(n875), .B0(n464), .Y(n514) );
  INVXL U407 ( .A(n463), .Y(n464) );
  OAI2BB1XL U408 ( .A0N(n879), .A1N(n791), .B0(n469), .Y(n487) );
  INVXL U409 ( .A(n468), .Y(n469) );
  OAI22XL U410 ( .A0(n1076), .A1(n472), .B0(n1077), .B1(n485), .Y(n490) );
  OAI22XL U411 ( .A0(n1135), .A1(n470), .B0(n1148), .B1(n482), .Y(n492) );
  CMPR32X1 U412 ( .A(n404), .B(n403), .C(n402), .CO(n409), .S(n411) );
  OAI22XL U413 ( .A0(n391), .A1(n289), .B0(n397), .B1(n390), .Y(n404) );
  XNOR2XL U414 ( .A(A[3]), .B(B[4]), .Y(n316) );
  OAI22XL U415 ( .A0(n875), .A1(n5), .B0(n873), .B1(n318), .Y(n328) );
  XNOR2XL U416 ( .A(A[3]), .B(B[3]), .Y(n325) );
  NOR2BXL U417 ( .AN(B[0]), .B(n879), .Y(n321) );
  OAI22X1 U418 ( .A0(n859), .A1(n317), .B0(n308), .B1(n1064), .Y(n320) );
  OAI22XL U419 ( .A0(n875), .A1(n326), .B0(n873), .B1(n309), .Y(n319) );
  INVXL U420 ( .A(n1209), .Y(n1210) );
  AOI21XL U421 ( .A0(n1208), .A1(n1207), .B0(n1206), .Y(n1209) );
  INVXL U422 ( .A(n1219), .Y(n1206) );
  OAI2BB1XL U423 ( .A0N(n1127), .A1N(n1126), .B0(n1125), .Y(n1136) );
  OAI22XL U424 ( .A0(n1165), .A1(n1123), .B0(n1163), .B1(n1133), .Y(n1137) );
  INVXL U425 ( .A(n1124), .Y(n1125) );
  INVXL U426 ( .A(n1138), .Y(n1120) );
  OAI22XL U427 ( .A0(n1135), .A1(n1095), .B0(n1148), .B1(n1119), .Y(n1122) );
  OAI22XL U428 ( .A0(n1165), .A1(n1096), .B0(n1163), .B1(n1123), .Y(n1121) );
  OAI22XL U429 ( .A0(n1098), .A1(n1079), .B0(n1127), .B1(n1097), .Y(n1101) );
  OAI22XL U430 ( .A0(n1135), .A1(n1080), .B0(n1148), .B1(n1095), .Y(n1100) );
  CMPR32X1 U431 ( .A(n871), .B(n870), .C(n869), .CO(n890), .S(n924) );
  AND2X1 U432 ( .A(n69), .B(n276), .Y(n940) );
  INVX1 U433 ( .A(n668), .Y(n90) );
  OAI22XL U434 ( .A0(n1147), .A1(n579), .B0(n1148), .B1(n577), .Y(n621) );
  OR2X2 U435 ( .A(n1060), .B(n1172), .Y(n83) );
  NAND2XL U436 ( .A(A[1]), .B(n747), .Y(n820) );
  OAI21XL U437 ( .A0(n365), .A1(n1176), .B0(n364), .Y(n1059) );
  NAND2X1 U438 ( .A(n105), .B(n1179), .Y(n364) );
  AOI21XL U439 ( .A0(n1192), .A1(n337), .B0(n340), .Y(n1189) );
  INVXL U440 ( .A(n1191), .Y(n340) );
  NOR2XL U441 ( .A(n349), .B(n348), .Y(n1186) );
  NAND2XL U442 ( .A(n349), .B(n348), .Y(n1187) );
  OAI22XL U443 ( .A0(n1165), .A1(n1164), .B0(n1163), .B1(n1162), .Y(n1166) );
  OAI2BB1XL U444 ( .A0N(n1148), .A1N(n1147), .B0(n1146), .Y(n1157) );
  OAI22XL U445 ( .A0(n1165), .A1(n1144), .B0(n1163), .B1(n1164), .Y(n1158) );
  INVXL U446 ( .A(n1145), .Y(n1146) );
  OAI22XL U447 ( .A0(n859), .A1(B[0]), .B0(n330), .B1(n1064), .Y(n1199) );
  NAND2XL U448 ( .A(n331), .B(n820), .Y(n1198) );
  NAND2BXL U449 ( .AN(B[0]), .B(n581), .Y(n331) );
  NAND2XL U450 ( .A(n1199), .B(n1198), .Y(n1200) );
  INVXL U451 ( .A(n1176), .Y(n1184) );
  NOR2X1 U452 ( .A(n769), .B(n1246), .Y(n76) );
  INVXL U453 ( .A(n1225), .Y(n1107) );
  NAND2X1 U454 ( .A(n424), .B(n735), .Y(n425) );
  OAI21XL U455 ( .A0(n1251), .A1(n1248), .B0(n1249), .Y(n737) );
  NOR2X1 U456 ( .A(n1244), .B(n1246), .Y(n424) );
  INVXL U457 ( .A(n1151), .Y(n1109) );
  AOI21XL U458 ( .A0(n1212), .A1(n1104), .B0(n1107), .Y(n1065) );
  INVXL U459 ( .A(n1231), .Y(n446) );
  INVX1 U460 ( .A(n1259), .Y(n125) );
  NAND2BXL U461 ( .AN(n895), .B(n426), .Y(n123) );
  NAND3XL U462 ( .A(n803), .B(n426), .C(n735), .Y(n86) );
  INVXL U463 ( .A(n737), .Y(n770) );
  INVXL U464 ( .A(n1246), .Y(n771) );
  INVXL U465 ( .A(n1242), .Y(n704) );
  NAND3XL U466 ( .A(n803), .B(n426), .C(n76), .Y(n73) );
  AOI21XL U467 ( .A0(n846), .A1(n76), .B0(n75), .Y(n74) );
  NAND2BXL U468 ( .AN(n770), .B(n771), .Y(n77) );
  INVXL U469 ( .A(n1118), .Y(n165) );
  XNOR2XL U470 ( .A(n1078), .B(B[0]), .Y(n395) );
  XNOR2XL U471 ( .A(n1078), .B(B[1]), .Y(n394) );
  XNOR2XL U472 ( .A(n581), .B(B[11]), .Y(n242) );
  INVXL U473 ( .A(n1229), .Y(n445) );
  AOI21XL U474 ( .A0(n1107), .A1(n1106), .B0(n1105), .Y(n1152) );
  INVXL U475 ( .A(n1223), .Y(n1105) );
  NAND2XL U476 ( .A(n1104), .B(n1106), .Y(n1151) );
  NOR2X1 U477 ( .A(n425), .B(n847), .Y(n96) );
  AOI21XL U478 ( .A0(n1212), .A1(n1109), .B0(n1108), .Y(n1110) );
  INVXL U479 ( .A(n1152), .Y(n1108) );
  NAND2XL U480 ( .A(n427), .B(n1109), .Y(n1111) );
  INVXL U481 ( .A(n1236), .Y(n603) );
  NAND2X1 U482 ( .A(n108), .B(n930), .Y(n107) );
  NAND2X1 U483 ( .A(n736), .B(n126), .Y(n850) );
  XNOR2X2 U484 ( .A(n809), .B(n808), .Y(PRODUCT[24]) );
  INVXL U485 ( .A(n1248), .Y(n807) );
  XOR2X1 U486 ( .A(n72), .B(n61), .Y(PRODUCT[26]) );
  INVXL U487 ( .A(n1244), .Y(n738) );
  NAND2X1 U488 ( .A(n116), .B(n637), .Y(n640) );
  INVXL U489 ( .A(n599), .Y(n637) );
  INVXL U490 ( .A(n1232), .Y(n531) );
  XNOR2XL U491 ( .A(n833), .B(B[15]), .Y(n790) );
  XNOR2XL U492 ( .A(n462), .B(B[16]), .Y(n831) );
  XNOR2XL U493 ( .A(n833), .B(B[14]), .Y(n834) );
  XNOR2XL U494 ( .A(n581), .B(B[16]), .Y(n169) );
  XNOR2XL U495 ( .A(n833), .B(B[13]), .Y(n878) );
  XNOR2XL U496 ( .A(n1161), .B(n821), .Y(n860) );
  XNOR2XL U497 ( .A(n1161), .B(B[4]), .Y(n861) );
  XNOR2XL U498 ( .A(n823), .B(B[9]), .Y(n262) );
  XNOR2XL U499 ( .A(n1078), .B(B[4]), .Y(n181) );
  XNOR2X1 U500 ( .A(n462), .B(n788), .Y(n162) );
  XNOR2XL U501 ( .A(n833), .B(B[8]), .Y(n183) );
  OAI22XL U502 ( .A0(n866), .A1(n396), .B0(n397), .B1(n227), .Y(n1007) );
  XNOR2XL U503 ( .A(n1161), .B(B[11]), .Y(n650) );
  XNOR2XL U504 ( .A(B[23]), .B(A[3]), .Y(n652) );
  XNOR2X1 U505 ( .A(n833), .B(B[21]), .Y(n578) );
  XNOR2XL U506 ( .A(n1118), .B(B[14]), .Y(n618) );
  XNOR2XL U507 ( .A(n833), .B(B[20]), .Y(n624) );
  XNOR2XL U508 ( .A(A[15]), .B(B[16]), .Y(n508) );
  INVXL U509 ( .A(n823), .Y(n465) );
  NAND2BXL U510 ( .AN(B[0]), .B(n462), .Y(n318) );
  XNOR2XL U511 ( .A(n581), .B(B[5]), .Y(n317) );
  AOI21XL U512 ( .A0(n1212), .A1(n1205), .B0(n1208), .Y(n1153) );
  AOI21XL U513 ( .A0(n431), .A1(n445), .B0(n430), .Y(n432) );
  INVXL U514 ( .A(n1227), .Y(n430) );
  INVXL U515 ( .A(A[15]), .Y(n460) );
  XNOR2XL U516 ( .A(A[15]), .B(B[22]), .Y(n1123) );
  XNOR2XL U517 ( .A(n1118), .B(B[23]), .Y(n1095) );
  XNOR2XL U518 ( .A(n1078), .B(B[25]), .Y(n1097) );
  CMPR32X1 U519 ( .A(n698), .B(n697), .C(n696), .CO(n711), .S(n742) );
  OAI22XL U520 ( .A0(n1098), .A1(n691), .B0(n1127), .B1(n658), .Y(n697) );
  OAI22XL U521 ( .A0(n875), .A1(n690), .B0(n873), .B1(n657), .Y(n698) );
  ADDFX2 U522 ( .A(n763), .B(n762), .CI(n761), .CO(n777), .S(n813) );
  OAI22X1 U523 ( .A0(n1098), .A1(n756), .B0(n1127), .B1(n722), .Y(n762) );
  OAI22XL U524 ( .A0(n1135), .A1(n752), .B0(n1148), .B1(n717), .Y(n758) );
  OAI22XL U525 ( .A0(n1135), .A1(n784), .B0(n1148), .B1(n752), .Y(n792) );
  CMPR32X1 U526 ( .A(n840), .B(n839), .C(n838), .CO(n856), .S(n901) );
  OAI22XL U527 ( .A0(n791), .A1(n834), .B0(n879), .B1(n790), .Y(n838) );
  OAI22XL U528 ( .A0(n1098), .A1(n832), .B0(n1127), .B1(n789), .Y(n839) );
  OAI22X1 U529 ( .A0(n274), .A1(n1064), .B0(n859), .B1(n169), .Y(n69) );
  ADDFX2 U530 ( .A(n919), .B(n918), .CI(n917), .CO(n911), .S(n960) );
  OAI22XL U531 ( .A0(n1135), .A1(n868), .B0(n1148), .B1(n867), .Y(n917) );
  OAI22X1 U532 ( .A0(n121), .A1(n864), .B0(n866), .B1(n865), .Y(n918) );
  OAI22XL U533 ( .A0(n881), .A1(n267), .B0(n879), .B1(n880), .Y(n914) );
  OAI22XL U534 ( .A0(n875), .A1(n265), .B0(n873), .B1(n874), .Y(n916) );
  OAI22XL U535 ( .A0(n1135), .A1(n177), .B0(n1148), .B1(n176), .Y(n184) );
  OAI22XL U536 ( .A0(n866), .A1(n178), .B0(n864), .B1(n175), .Y(n185) );
  OAI22XL U537 ( .A0(n875), .A1(n148), .B0(n341), .B1(n145), .Y(n189) );
  OAI21XL U538 ( .A0(n102), .A1(n101), .B0(n100), .Y(n166) );
  INVXL U539 ( .A(n161), .Y(n101) );
  INVXL U540 ( .A(n103), .Y(n102) );
  CMPR32X1 U541 ( .A(n195), .B(n194), .C(n193), .CO(n192), .S(n231) );
  OAI22XL U542 ( .A0(n881), .A1(n183), .B0(n879), .B1(n182), .Y(n193) );
  OAI22XL U543 ( .A0(n1098), .A1(n181), .B0(n1127), .B1(n180), .Y(n194) );
  OAI22XL U544 ( .A0(n866), .A1(n179), .B0(n864), .B1(n178), .Y(n195) );
  NOR2BXL U545 ( .AN(B[0]), .B(n1163), .Y(n201) );
  OAI22XL U546 ( .A0(n1135), .A1(n216), .B0(n1148), .B1(n158), .Y(n199) );
  OAI22X1 U547 ( .A0(n866), .A1(n227), .B0(n864), .B1(n203), .Y(n239) );
  OAI22XL U548 ( .A0(n1135), .A1(n217), .B0(n1148), .B1(n216), .Y(n236) );
  OAI22XL U549 ( .A0(n1098), .A1(n225), .B0(n1127), .B1(n218), .Y(n235) );
  OAI22XL U550 ( .A0(n1076), .A1(n372), .B0(n1077), .B1(n241), .Y(n1014) );
  OAI22XL U551 ( .A0(n791), .A1(n624), .B0(n879), .B1(n578), .Y(n615) );
  OAI22XL U552 ( .A0(n866), .A1(n617), .B0(n864), .B1(n586), .Y(n630) );
  OAI2BB1XL U553 ( .A0N(n864), .A1N(n866), .B0(n535), .Y(n552) );
  OAI22XL U554 ( .A0(n881), .A1(n549), .B0(n879), .B1(n544), .Y(n555) );
  INVXL U555 ( .A(n488), .Y(n476) );
  OAI22XL U556 ( .A0(n1098), .A1(n506), .B0(n1127), .B1(n475), .Y(n511) );
  OAI22XL U557 ( .A0(n881), .A1(n507), .B0(n879), .B1(n473), .Y(n513) );
  CMPR32X1 U558 ( .A(n383), .B(n382), .C(n381), .CO(n405), .S(n413) );
  OAI22XL U559 ( .A0(n1076), .A1(n286), .B0(n1077), .B1(n379), .Y(n382) );
  OAI22XL U560 ( .A0(n371), .A1(n388), .B0(n873), .B1(n370), .Y(n1005) );
  XNOR2XL U561 ( .A(n581), .B(B[3]), .Y(n343) );
  NOR2BXL U562 ( .AN(B[0]), .B(n1077), .Y(n295) );
  OAI22XL U563 ( .A0(n881), .A1(n297), .B0(n879), .B1(n292), .Y(n293) );
  OAI22X1 U564 ( .A0(n82), .A1(n859), .B0(n291), .B1(n1064), .Y(n294) );
  INVXL U565 ( .A(n833), .Y(n466) );
  OAI22XL U566 ( .A0(n881), .A1(n298), .B0(n879), .B1(n297), .Y(n311) );
  OAI22XL U567 ( .A0(n875), .A1(n309), .B0(n873), .B1(n299), .Y(n310) );
  OAI22XL U568 ( .A0(n866), .A1(n35), .B0(n864), .B1(n336), .Y(n338) );
  NAND2BXL U569 ( .AN(B[0]), .B(A[3]), .Y(n336) );
  OAI22XL U570 ( .A0(n859), .A1(n330), .B0(n334), .B1(n1064), .Y(n333) );
  NOR2BXL U571 ( .AN(B[0]), .B(n397), .Y(n332) );
  OAI2BB1XL U572 ( .A0N(n1077), .A1N(n1076), .B0(n1075), .Y(n1092) );
  OAI22XL U573 ( .A0(n1165), .A1(n1073), .B0(n1163), .B1(n1096), .Y(n1094) );
  INVXL U574 ( .A(n1074), .Y(n1075) );
  XOR2XL U575 ( .A(n104), .B(n103), .Y(n213) );
  XOR2XL U576 ( .A(n160), .B(n161), .Y(n104) );
  OAI22XL U577 ( .A0(n1135), .A1(n482), .B0(n1148), .B1(n1080), .Y(n1083) );
  OAI22XL U578 ( .A0(n484), .A1(n483), .B0(n1163), .B1(n1073), .Y(n1082) );
  INVXL U579 ( .A(n1093), .Y(n1081) );
  OAI22XL U580 ( .A0(n1098), .A1(n486), .B0(n1127), .B1(n1079), .Y(n1086) );
  OAI22XL U581 ( .A0(n1076), .A1(n510), .B0(n1077), .B1(n505), .Y(n519) );
  OAI22XL U582 ( .A0(n1098), .A1(n475), .B0(n1127), .B1(n471), .Y(n481) );
  OAI22XL U583 ( .A0(n484), .A1(n461), .B0(n1163), .B1(n467), .Y(n480) );
  ADDFX2 U584 ( .A(n324), .B(n65), .CI(n322), .CO(n362), .S(n361) );
  OAI22XL U585 ( .A0(n866), .A1(n325), .B0(n397), .B1(n316), .Y(n324) );
  NAND2XL U586 ( .A(n427), .B(n1211), .Y(n1214) );
  NAND2XL U587 ( .A(n339), .B(n338), .Y(n1191) );
  NOR2XL U588 ( .A(n333), .B(n332), .Y(n1194) );
  NAND2XL U589 ( .A(n333), .B(n332), .Y(n1195) );
  OAI22XL U590 ( .A0(n1165), .A1(n1133), .B0(n1163), .B1(n1144), .Y(n1143) );
  INVXL U591 ( .A(n1159), .Y(n1142) );
  OAI22XL U592 ( .A0(n1135), .A1(n1119), .B0(n1148), .B1(n1134), .Y(n1132) );
  OAI21XL U593 ( .A0(n572), .A1(n573), .B0(n571), .Y(n98) );
  NAND2XL U594 ( .A(n731), .B(n732), .Y(n109) );
  NAND2XL U595 ( .A(n889), .B(n890), .Y(n70) );
  OAI21XL U596 ( .A0(n899), .A1(n900), .B0(n898), .Y(n118) );
  XNOR3X2 U597 ( .A(n900), .B(n898), .C(n119), .Y(n927) );
  OAI2BB1X1 U598 ( .A0N(n68), .A1N(n965), .B0(n67), .Y(n957) );
  OR2X2 U599 ( .A(n967), .B(n966), .Y(n68) );
  OAI2BB1X1 U600 ( .A0N(n285), .A1N(n284), .B0(n99), .Y(n982) );
  OAI21XL U601 ( .A0(n284), .A1(n285), .B0(n283), .Y(n99) );
  NOR2X1 U602 ( .A(n258), .B(n257), .Y(n992) );
  NAND2XL U603 ( .A(n257), .B(n258), .Y(n993) );
  NAND2BXL U604 ( .AN(n667), .B(n90), .Y(n89) );
  CLKINVX3 U605 ( .A(mult_x_1_n335), .Y(n1050) );
  AOI21X1 U606 ( .A0(n58), .A1(n1049), .B0(n1038), .Y(n1044) );
  NAND2X1 U607 ( .A(n80), .B(n1059), .Y(n79) );
  NOR2X1 U608 ( .A(n1171), .B(n1060), .Y(n80) );
  NAND2X1 U609 ( .A(n362), .B(n363), .Y(n1178) );
  NAND2XL U610 ( .A(n802), .B(n801), .Y(mult_x_1_n242) );
  NAND2XL U611 ( .A(n1088), .B(n1087), .Y(mult_x_1_n150) );
  INVXL U612 ( .A(n1060), .Y(n84) );
  NAND2XL U613 ( .A(n1183), .B(n1182), .Y(n1185) );
  XOR2XL U614 ( .A(n1190), .B(n1189), .Y(n1298) );
  NAND2XL U615 ( .A(n1188), .B(n1187), .Y(n1190) );
  INVXL U616 ( .A(n1186), .Y(n1188) );
  XNOR2XL U617 ( .A(n1193), .B(n1192), .Y(n1299) );
  NAND2XL U618 ( .A(n337), .B(n1191), .Y(n1193) );
  XOR2XL U619 ( .A(n1197), .B(n1200), .Y(n1300) );
  NAND2XL U620 ( .A(n1196), .B(n1195), .Y(n1197) );
  INVXL U621 ( .A(n1194), .Y(n1196) );
  NAND2XL U622 ( .A(n969), .B(n968), .Y(mult_x_1_n289) );
  NAND2XL U623 ( .A(n1170), .B(n1169), .Y(mult_x_1_n54) );
  NAND2XL U624 ( .A(n1168), .B(n1167), .Y(n1169) );
  INVXL U625 ( .A(n1166), .Y(n1167) );
  NOR2XL U626 ( .A(n1150), .B(n1149), .Y(mult_x_1_n105) );
  NAND2XL U627 ( .A(n1150), .B(n1149), .Y(mult_x_1_n106) );
  NOR2XL U628 ( .A(n1140), .B(n1139), .Y(mult_x_1_n114) );
  NAND2XL U629 ( .A(n1140), .B(n1139), .Y(mult_x_1_n115) );
  NOR2XL U630 ( .A(n1129), .B(n1128), .Y(mult_x_1_n125) );
  NAND2XL U631 ( .A(n1129), .B(n1128), .Y(mult_x_1_n126) );
  NOR2XL U632 ( .A(n1103), .B(n1102), .Y(mult_x_1_n134) );
  NAND2XL U633 ( .A(n1103), .B(n1102), .Y(mult_x_1_n135) );
  NOR2XL U634 ( .A(n1088), .B(n1087), .Y(mult_x_1_n149) );
  NOR2XL U635 ( .A(mult_x_1_n302), .B(mult_x_1_n299), .Y(mult_x_1_n297) );
  NOR2X1 U636 ( .A(n988), .B(n987), .Y(mult_x_1_n302) );
  OAI21XL U637 ( .A0(n992), .A1(mult_x_1_n313), .B0(n993), .Y(mult_x_1_n306)
         );
  OAI21XL U638 ( .A0(n1050), .A1(n1045), .B0(n1044), .Y(mult_x_1_n320) );
  NAND2XL U639 ( .A(n356), .B(n1202), .Y(n1204) );
  NAND2XL U640 ( .A(n1179), .B(n1178), .Y(n1180) );
  AOI21XL U641 ( .A0(n1184), .A1(n1183), .B0(n1177), .Y(n1181) );
  NOR2BXL U642 ( .AN(B[0]), .B(n1064), .Y(n1302) );
  BUFX3 U643 ( .A(A[5]), .Y(n462) );
  OR2X2 U644 ( .A(n1037), .B(n1036), .Y(n58) );
  OR2X2 U645 ( .A(n418), .B(n417), .Y(n62) );
  AND2X2 U646 ( .A(n83), .B(n1061), .Y(n63) );
  NOR2X1 U647 ( .A(n369), .B(n368), .Y(n1060) );
  NAND2X1 U648 ( .A(n928), .B(n422), .Y(n847) );
  INVX1 U649 ( .A(n847), .Y(n803) );
  BUFX3 U650 ( .A(A[7]), .Y(n833) );
  CMPR22X1 U651 ( .A(n307), .B(n306), .CO(n300), .S(n315) );
  OAI22X1 U652 ( .A0(n82), .A1(n1064), .B0(n308), .B1(n859), .Y(n307) );
  OAI22X1 U653 ( .A0(n1165), .A1(n683), .B0(n1163), .B1(n650), .Y(n680) );
  OAI22X1 U654 ( .A0(n1165), .A1(n749), .B0(n1163), .B1(n715), .Y(n745) );
  OAI22X1 U655 ( .A0(n1165), .A1(n822), .B0(n1163), .B1(n781), .Y(n816) );
  OAI22X1 U656 ( .A0(n1165), .A1(n861), .B0(n1163), .B1(n860), .Y(n904) );
  OAI22X1 U657 ( .A0(n881), .A1(n473), .B0(n879), .B1(n468), .Y(n488) );
  BUFX3 U658 ( .A(A[9]), .Y(n823) );
  OAI22X1 U659 ( .A0(n875), .A1(n542), .B0(n873), .B1(n463), .Y(n515) );
  BUFX1 U660 ( .A(n323), .Y(n65) );
  ADDHXL U661 ( .A(n223), .B(n222), .CO(n219), .S(n999) );
  OAI22X1 U662 ( .A0(n1165), .A1(n781), .B0(n1163), .B1(n749), .Y(n778) );
  OAI22X1 U663 ( .A0(n1165), .A1(n715), .B0(n1163), .B1(n683), .Y(n712) );
  OAI22X1 U664 ( .A0(n881), .A1(n387), .B0(n879), .B1(n393), .Y(n401) );
  NAND2X1 U665 ( .A(n896), .B(n1253), .Y(n897) );
  XOR2X1 U666 ( .A(n124), .B(n955), .Y(PRODUCT[20]) );
  XOR2X1 U667 ( .A(n120), .B(n857), .Y(n913) );
  AND2X2 U668 ( .A(n120), .B(n857), .Y(n870) );
  INVX1 U669 ( .A(n426), .Y(n953) );
  XNOR2X1 U670 ( .A(B[15]), .B(n1161), .Y(n534) );
  XNOR2X1 U671 ( .A(n581), .B(B[15]), .Y(n153) );
  XOR3X2 U672 ( .A(n966), .B(n967), .C(n965), .Y(n970) );
  OAI2BB1X1 U673 ( .A0N(n64), .A1N(n888), .B0(n70), .Y(n852) );
  NAND2X2 U674 ( .A(n79), .B(n63), .Y(n1058) );
  NAND2X2 U675 ( .A(n420), .B(n81), .Y(mult_x_1_n335) );
  OAI2BB1X1 U676 ( .A0N(n89), .A1N(n666), .B0(n88), .Y(n642) );
  XNOR3X2 U677 ( .A(n667), .B(n90), .C(n666), .Y(n674) );
  XNOR2X1 U678 ( .A(n818), .B(n823), .Y(n91) );
  XOR2X1 U679 ( .A(n589), .B(n95), .Y(n645) );
  NAND2X2 U680 ( .A(n114), .B(n115), .Y(n846) );
  XOR2X2 U681 ( .A(n107), .B(n59), .Y(PRODUCT[21]) );
  XOR2X1 U682 ( .A(n730), .B(n112), .Y(n739) );
  XOR2X1 U683 ( .A(n731), .B(n732), .Y(n112) );
  NOR2BX1 U684 ( .AN(n1253), .B(n134), .Y(n114) );
  NAND2X1 U685 ( .A(n929), .B(n422), .Y(n115) );
  CMPR22X1 U686 ( .A(n172), .B(n171), .CO(n272), .S(n168) );
  OAI22X1 U687 ( .A0(n859), .A1(n152), .B0(n153), .B1(n1064), .Y(n155) );
  XOR2X1 U688 ( .A(n825), .B(n35), .Y(n121) );
  XOR2X2 U689 ( .A(n122), .B(n897), .Y(PRODUCT[22]) );
  OAI21X1 U690 ( .A0(n530), .A1(n1215), .B0(n128), .Y(n533) );
  AND2X2 U691 ( .A(n737), .B(n424), .Y(n130) );
  OAI21X1 U692 ( .A0(n1215), .A1(n602), .B0(n601), .Y(n605) );
  NOR2X1 U693 ( .A(n1252), .B(n1255), .Y(n134) );
  NOR2X1 U694 ( .A(n1252), .B(n1254), .Y(n422) );
  OAI21X1 U695 ( .A0(n1256), .A1(n1259), .B0(n1257), .Y(n929) );
  OAI21XL U696 ( .A0(n1244), .A1(n1247), .B0(n1245), .Y(n423) );
  OAI22X1 U697 ( .A0(n1076), .A1(n862), .B0(n1077), .B1(n824), .Y(n884) );
  AOI21XL U698 ( .A0(n929), .A1(n932), .B0(n893), .Y(n894) );
  XNOR2XL U699 ( .A(A[13]), .B(B[11]), .Y(n717) );
  XNOR2XL U700 ( .A(n1185), .B(n1184), .Y(n1296) );
  XOR2XL U701 ( .A(A[4]), .B(A[5]), .Y(n135) );
  XNOR2X1 U702 ( .A(A[4]), .B(A[3]), .Y(n341) );
  BUFX3 U703 ( .A(n371), .Y(n875) );
  XNOR2X1 U704 ( .A(n462), .B(B[12]), .Y(n145) );
  BUFX3 U705 ( .A(n1126), .Y(n1098) );
  BUFX3 U706 ( .A(A[11]), .Y(n1078) );
  INVXL U707 ( .A(n1078), .Y(n244) );
  XNOR2X1 U708 ( .A(A[11]), .B(n821), .Y(n180) );
  BUFX3 U709 ( .A(n137), .Y(n1127) );
  XNOR2X1 U710 ( .A(A[11]), .B(B[6]), .Y(n146) );
  OAI22XL U711 ( .A0(n1098), .A1(n180), .B0(n1127), .B1(n146), .Y(n188) );
  XOR2XL U712 ( .A(A[6]), .B(A[7]), .Y(n138) );
  BUFX3 U713 ( .A(n791), .Y(n881) );
  BUFX3 U714 ( .A(n139), .Y(n879) );
  BUFX3 U715 ( .A(B[10]), .Y(n788) );
  OAI22XL U716 ( .A0(n881), .A1(n182), .B0(n879), .B1(n147), .Y(n187) );
  XOR2XL U717 ( .A(A[8]), .B(A[9]), .Y(n140) );
  XNOR2XL U718 ( .A(A[8]), .B(A[7]), .Y(n141) );
  NAND2X1 U719 ( .A(n140), .B(n141), .Y(n380) );
  BUFX3 U720 ( .A(n380), .Y(n1076) );
  BUFX3 U721 ( .A(n141), .Y(n1077) );
  OAI22XL U722 ( .A0(n1076), .A1(n173), .B0(n1077), .B1(n262), .Y(n279) );
  BUFX3 U723 ( .A(n391), .Y(n866) );
  BUFX3 U724 ( .A(n397), .Y(n864) );
  XNOR2X1 U725 ( .A(A[3]), .B(B[15]), .Y(n263) );
  OAI22X1 U726 ( .A0(n866), .A1(n175), .B0(n864), .B1(n263), .Y(n278) );
  XOR2XL U727 ( .A(A[12]), .B(A[13]), .Y(n143) );
  BUFX3 U728 ( .A(n1147), .Y(n1135) );
  BUFX1 U729 ( .A(A[13]), .Y(n1118) );
  XNOR2X1 U730 ( .A(A[13]), .B(B[4]), .Y(n176) );
  BUFX3 U731 ( .A(n144), .Y(n1148) );
  XNOR2X1 U732 ( .A(A[13]), .B(n821), .Y(n264) );
  BUFX3 U733 ( .A(n341), .Y(n873) );
  OAI22XL U734 ( .A0(n371), .A1(n145), .B0(n873), .B1(n265), .Y(n261) );
  XNOR2X1 U735 ( .A(A[11]), .B(n826), .Y(n266) );
  OAI22XL U736 ( .A0(n1098), .A1(n146), .B0(n1127), .B1(n266), .Y(n260) );
  OAI22XL U737 ( .A0(n875), .A1(n162), .B0(n873), .B1(n148), .Y(n198) );
  BUFX3 U738 ( .A(n820), .Y(n859) );
  BUFX3 U739 ( .A(n747), .Y(n1064) );
  XOR2XL U740 ( .A(A[14]), .B(A[15]), .Y(n149) );
  XNOR2XL U741 ( .A(A[14]), .B(A[13]), .Y(n150) );
  BUFX3 U742 ( .A(n484), .Y(n1165) );
  BUFX3 U743 ( .A(n150), .Y(n1163) );
  CLKINVX3 U744 ( .A(n460), .Y(n1161) );
  OAI22X1 U745 ( .A0(n1165), .A1(n460), .B0(n1163), .B1(n151), .Y(n154) );
  XNOR2X1 U746 ( .A(n581), .B(B[13]), .Y(n163) );
  OAI22X1 U747 ( .A0(n859), .A1(n163), .B0(n152), .B1(n1064), .Y(n200) );
  XNOR2XL U748 ( .A(n1118), .B(B[1]), .Y(n216) );
  OAI22X1 U749 ( .A0(n859), .A1(n153), .B0(n169), .B1(n1064), .Y(n172) );
  XNOR2XL U750 ( .A(n1161), .B(B[1]), .Y(n156) );
  XNOR2X1 U751 ( .A(n1161), .B(B[2]), .Y(n170) );
  OAI22X1 U752 ( .A0(n1165), .A1(n156), .B0(n1163), .B1(n170), .Y(n171) );
  CMPR22X1 U753 ( .A(n155), .B(n154), .CO(n167), .S(n197) );
  XNOR2XL U754 ( .A(n823), .B(B[6]), .Y(n159) );
  XNOR2X1 U755 ( .A(n823), .B(n826), .Y(n174) );
  XNOR2XL U756 ( .A(n1161), .B(B[0]), .Y(n157) );
  XNOR2X1 U757 ( .A(n1118), .B(B[3]), .Y(n177) );
  OAI22X1 U758 ( .A0(n1135), .A1(n158), .B0(n1148), .B1(n177), .Y(n160) );
  XNOR2X1 U759 ( .A(n823), .B(n821), .Y(n202) );
  OAI22XL U760 ( .A0(n380), .A1(n202), .B0(n1077), .B1(n159), .Y(n207) );
  OAI22XL U761 ( .A0(n1098), .A1(n218), .B0(n1127), .B1(n181), .Y(n206) );
  XNOR2X1 U762 ( .A(A[3]), .B(B[11]), .Y(n203) );
  XNOR2X1 U763 ( .A(A[3]), .B(B[12]), .Y(n179) );
  OAI22XL U764 ( .A0(n866), .A1(n203), .B0(n397), .B1(n179), .Y(n205) );
  OAI22XL U765 ( .A0(n875), .A1(n204), .B0(n873), .B1(n162), .Y(n221) );
  XNOR2X1 U766 ( .A(n581), .B(B[12]), .Y(n224) );
  CMPR32X1 U767 ( .A(n168), .B(n167), .C(n166), .CO(n270), .S(n209) );
  BUFX3 U768 ( .A(B[17]), .Y(n825) );
  XNOR2X1 U769 ( .A(n581), .B(n825), .Y(n274) );
  XNOR2X1 U770 ( .A(n1161), .B(B[3]), .Y(n275) );
  OAI22XL U771 ( .A0(n380), .A1(n174), .B0(n1077), .B1(n173), .Y(n186) );
  CMPR32X1 U772 ( .A(n186), .B(n185), .C(n184), .CO(n271), .S(n191) );
  CMPR32X1 U773 ( .A(n189), .B(n188), .C(n187), .CO(n282), .S(n190) );
  CMPR32X1 U774 ( .A(n198), .B(n197), .C(n196), .CO(n210), .S(n230) );
  ADDFHX1 U775 ( .A(n201), .B(n200), .CI(n199), .CO(n196), .S(n234) );
  OAI22XL U776 ( .A0(n1076), .A1(n241), .B0(n1077), .B1(n202), .Y(n240) );
  OAI22XL U777 ( .A0(n875), .A1(n228), .B0(n873), .B1(n204), .Y(n238) );
  XOR2X2 U778 ( .A(n953), .B(n211), .Y(PRODUCT[19]) );
  CMPR32X1 U779 ( .A(n214), .B(n213), .C(n212), .CO(n208), .S(n256) );
  XNOR2XL U780 ( .A(n833), .B(B[6]), .Y(n226) );
  OAI22XL U781 ( .A0(n881), .A1(n226), .B0(n879), .B1(n215), .Y(n237) );
  XNOR2XL U782 ( .A(n1118), .B(B[0]), .Y(n217) );
  OAI22X1 U783 ( .A0(n859), .A1(n242), .B0(n224), .B1(n1064), .Y(n246) );
  OAI22XL U784 ( .A0(n881), .A1(n392), .B0(n879), .B1(n226), .Y(n1008) );
  XNOR2X1 U785 ( .A(n462), .B(n826), .Y(n370) );
  OAI22XL U786 ( .A0(n875), .A1(n370), .B0(n341), .B1(n228), .Y(n1006) );
  ADDFHX1 U787 ( .A(n231), .B(n230), .CI(n229), .CO(n252), .S(n254) );
  CMPR32X1 U788 ( .A(n234), .B(n233), .C(n232), .CO(n229), .S(n1030) );
  CMPR32X1 U789 ( .A(n237), .B(n236), .C(n235), .CO(n250), .S(n1011) );
  ADDFHX1 U790 ( .A(n240), .B(n239), .CI(n238), .CO(n233), .S(n1010) );
  OAI22X1 U791 ( .A0(n1098), .A1(n244), .B0(n1127), .B1(n243), .Y(n373) );
  ADDFHX1 U792 ( .A(n247), .B(n246), .CI(n245), .CO(n998), .S(n1012) );
  CMPR32X1 U793 ( .A(n250), .B(n249), .C(n248), .CO(n255), .S(n1028) );
  NAND2XL U794 ( .A(n991), .B(n990), .Y(mult_x_1_n313) );
  CMPR32X1 U795 ( .A(n253), .B(n252), .C(n251), .CO(n987), .S(n258) );
  CMPR32X1 U796 ( .A(n261), .B(n260), .C(n259), .CO(n947), .S(n280) );
  OAI22XL U797 ( .A0(n1076), .A1(n262), .B0(n1077), .B1(n863), .Y(n910) );
  XNOR2X1 U798 ( .A(A[13]), .B(B[6]), .Y(n868) );
  XNOR2X1 U799 ( .A(n462), .B(B[14]), .Y(n874) );
  XNOR2X1 U800 ( .A(A[11]), .B(B[8]), .Y(n877) );
  OAI22XL U801 ( .A0(n1098), .A1(n266), .B0(n1127), .B1(n877), .Y(n915) );
  CMPR32X1 U802 ( .A(n273), .B(n272), .C(n271), .CO(n964), .S(n269) );
  BUFX3 U803 ( .A(B[18]), .Y(n783) );
  XNOR2X1 U804 ( .A(n581), .B(n783), .Y(n858) );
  OAI22X1 U805 ( .A0(n859), .A1(n274), .B0(n858), .B1(n1064), .Y(n907) );
  OAI22X1 U806 ( .A0(n1165), .A1(n275), .B0(n1163), .B1(n861), .Y(n906) );
  CMPR32X1 U807 ( .A(n279), .B(n278), .C(n277), .CO(n939), .S(n281) );
  CMPR32X1 U808 ( .A(n282), .B(n281), .C(n280), .CO(n962), .S(n285) );
  NOR2X1 U809 ( .A(n983), .B(n982), .Y(mult_x_1_n299) );
  XNOR2XL U810 ( .A(n833), .B(B[2]), .Y(n292) );
  OAI22XL U811 ( .A0(n881), .A1(n292), .B0(n879), .B1(n387), .Y(n383) );
  XNOR2XL U812 ( .A(n823), .B(B[0]), .Y(n286) );
  XNOR2XL U813 ( .A(n823), .B(B[1]), .Y(n379) );
  XNOR2X1 U814 ( .A(n462), .B(n821), .Y(n389) );
  OAI22XL U815 ( .A0(n875), .A1(n287), .B0(n341), .B1(n389), .Y(n381) );
  XNOR2X1 U816 ( .A(A[3]), .B(n821), .Y(n296) );
  XNOR2X1 U817 ( .A(A[3]), .B(B[6]), .Y(n289) );
  OAI22XL U818 ( .A0(n391), .A1(n296), .B0(n864), .B1(n289), .Y(n302) );
  XNOR2X1 U819 ( .A(n462), .B(B[3]), .Y(n299) );
  OAI22XL U820 ( .A0(n371), .A1(n299), .B0(n873), .B1(n287), .Y(n301) );
  OAI22X1 U821 ( .A0(n881), .A1(n466), .B0(n879), .B1(n288), .Y(n306) );
  XNOR2X1 U822 ( .A(A[3]), .B(n826), .Y(n390) );
  XNOR2X1 U823 ( .A(n581), .B(B[8]), .Y(n291) );
  XNOR2X1 U824 ( .A(n581), .B(B[9]), .Y(n377) );
  OAI22X1 U825 ( .A0(n859), .A1(n291), .B0(n377), .B1(n1064), .Y(n376) );
  OAI22X1 U826 ( .A0(n1076), .A1(n465), .B0(n1077), .B1(n290), .Y(n375) );
  XNOR2XL U827 ( .A(n833), .B(B[1]), .Y(n297) );
  CMPR32X1 U828 ( .A(n295), .B(n294), .C(n293), .CO(n402), .S(n305) );
  OAI22XL U829 ( .A0(n391), .A1(n316), .B0(n397), .B1(n296), .Y(n312) );
  XNOR2XL U830 ( .A(n833), .B(B[0]), .Y(n298) );
  XNOR2XL U831 ( .A(n462), .B(B[2]), .Y(n309) );
  CMPR32X1 U832 ( .A(n302), .B(n301), .C(n300), .CO(n412), .S(n303) );
  CMPR32X1 U833 ( .A(n305), .B(n304), .C(n303), .CO(n368), .S(n367) );
  XNOR2XL U834 ( .A(n462), .B(B[1]), .Y(n326) );
  CMPR32X1 U835 ( .A(n312), .B(n311), .C(n310), .CO(n304), .S(n313) );
  CMPR32X1 U836 ( .A(n315), .B(n314), .C(n313), .CO(n366), .S(n363) );
  OAI22XL U837 ( .A0(n859), .A1(n342), .B0(n317), .B1(n1064), .Y(n329) );
  CMPR32X1 U838 ( .A(n321), .B(n320), .C(n319), .CO(n314), .S(n322) );
  XNOR2XL U839 ( .A(A[3]), .B(B[2]), .Y(n344) );
  XNOR2XL U840 ( .A(n462), .B(B[0]), .Y(n327) );
  ADDHXL U841 ( .A(n329), .B(n328), .CO(n323), .S(n350) );
  OR2X2 U842 ( .A(n361), .B(n360), .Y(n1183) );
  XNOR2XL U843 ( .A(n581), .B(B[1]), .Y(n330) );
  XNOR2XL U844 ( .A(n581), .B(B[2]), .Y(n334) );
  OAI21XL U845 ( .A0(n1194), .A1(n1200), .B0(n1195), .Y(n1192) );
  OAI22X1 U846 ( .A0(n859), .A1(n334), .B0(n343), .B1(n1064), .Y(n347) );
  XNOR2XL U847 ( .A(A[3]), .B(B[0]), .Y(n335) );
  XNOR2XL U848 ( .A(A[3]), .B(B[1]), .Y(n345) );
  OAI22X1 U849 ( .A0(n866), .A1(n335), .B0(n397), .B1(n345), .Y(n346) );
  CMPR22X1 U850 ( .A(n347), .B(n346), .CO(n348), .S(n339) );
  OAI21XL U851 ( .A0(n1189), .A1(n1186), .B0(n1187), .Y(n1203) );
  CMPR32X1 U852 ( .A(n352), .B(n351), .C(n350), .CO(n360), .S(n358) );
  CMPR32X1 U853 ( .A(n355), .B(n354), .C(n353), .CO(n357), .S(n349) );
  NAND2XL U854 ( .A(n358), .B(n357), .Y(n1202) );
  INVXL U855 ( .A(n1202), .Y(n359) );
  AOI21XL U856 ( .A0(n1203), .A1(n356), .B0(n359), .Y(n1176) );
  NAND2XL U857 ( .A(n361), .B(n360), .Y(n1182) );
  INVXL U858 ( .A(n1182), .Y(n1177) );
  NAND2XL U859 ( .A(n369), .B(n368), .Y(n1061) );
  XNOR2X1 U860 ( .A(n462), .B(B[6]), .Y(n388) );
  XNOR2XL U861 ( .A(n823), .B(B[2]), .Y(n378) );
  OAI22X1 U862 ( .A0(n1076), .A1(n378), .B0(n1077), .B1(n372), .Y(n1004) );
  CMPR22X1 U863 ( .A(n374), .B(n373), .CO(n1013), .S(n1003) );
  CMPR22X1 U864 ( .A(n376), .B(n375), .CO(n407), .S(n403) );
  ADDFHX1 U865 ( .A(n386), .B(n385), .CI(n384), .CO(n1017), .S(n406) );
  XNOR2X1 U866 ( .A(n833), .B(B[4]), .Y(n393) );
  OAI22X1 U867 ( .A0(n875), .A1(n389), .B0(n873), .B1(n388), .Y(n400) );
  XNOR2X1 U868 ( .A(A[3]), .B(B[8]), .Y(n398) );
  OAI22XL U869 ( .A0(n391), .A1(n390), .B0(n397), .B1(n398), .Y(n399) );
  OAI22XL U870 ( .A0(n881), .A1(n393), .B0(n879), .B1(n392), .Y(n1002) );
  OAI22XL U871 ( .A0(n1098), .A1(n395), .B0(n1127), .B1(n394), .Y(n1001) );
  OAI22XL U872 ( .A0(n866), .A1(n398), .B0(n397), .B1(n396), .Y(n1000) );
  CMPR32X1 U873 ( .A(n413), .B(n412), .C(n411), .CO(n415), .S(n369) );
  NAND2XL U874 ( .A(n62), .B(n1056), .Y(n421) );
  NAND2XL U875 ( .A(n416), .B(n415), .Y(n1055) );
  INVXL U876 ( .A(n1055), .Y(n1051) );
  INVXL U877 ( .A(n1052), .Y(n419) );
  AOI21X1 U878 ( .A0(n62), .A1(n1051), .B0(n419), .Y(n420) );
  NOR2XL U879 ( .A(n1242), .B(n1240), .Y(n636) );
  NAND2XL U880 ( .A(n457), .B(n431), .Y(n433) );
  NOR2XL U881 ( .A(n1230), .B(n433), .Y(n435) );
  INVXL U882 ( .A(n427), .Y(n439) );
  OAI21XL U883 ( .A0(n1236), .A1(n1239), .B0(n1237), .Y(n428) );
  OAI21XL U884 ( .A0(n1232), .A1(n1235), .B0(n1233), .Y(n444) );
  OAI21XL U885 ( .A0(n433), .A1(n1231), .B0(n432), .Y(n434) );
  AOI21XL U886 ( .A0(n444), .A1(n435), .B0(n434), .Y(n436) );
  OAI21XL U887 ( .A0(n1215), .A1(n439), .B0(n438), .Y(n441) );
  INVXL U888 ( .A(n442), .Y(n498) );
  INVXL U889 ( .A(n1230), .Y(n502) );
  NAND2XL U890 ( .A(n502), .B(n457), .Y(n448) );
  NOR2XL U891 ( .A(n498), .B(n448), .Y(n450) );
  INVXL U892 ( .A(n444), .Y(n499) );
  AOI21XL U893 ( .A0(n446), .A1(n457), .B0(n445), .Y(n447) );
  OAI21XL U894 ( .A0(n499), .A1(n448), .B0(n447), .Y(n449) );
  AOI21XL U895 ( .A0(n566), .A1(n450), .B0(n449), .Y(n451) );
  NOR2XL U896 ( .A(n498), .B(n1230), .Y(n454) );
  NAND2XL U897 ( .A(n528), .B(n454), .Y(n456) );
  OAI21XL U898 ( .A0(n499), .A1(n1230), .B0(n1231), .Y(n453) );
  AOI21XL U899 ( .A0(n566), .A1(n454), .B0(n453), .Y(n455) );
  OAI21XL U900 ( .A0(n1215), .A1(n456), .B0(n455), .Y(n459) );
  XNOR2X1 U901 ( .A(n459), .B(n458), .Y(PRODUCT[34]) );
  XNOR2X1 U902 ( .A(A[15]), .B(n825), .Y(n461) );
  XNOR2X1 U903 ( .A(A[15]), .B(n783), .Y(n467) );
  OAI22XL U904 ( .A0(n484), .A1(n508), .B0(n1163), .B1(n461), .Y(n516) );
  BUFX3 U905 ( .A(B[26]), .Y(n1160) );
  OAI22XL U906 ( .A0(n1147), .A1(n474), .B0(n1148), .B1(n470), .Y(n478) );
  OAI22XL U907 ( .A0(n1076), .A1(n505), .B0(n1077), .B1(n472), .Y(n477) );
  OAI22XL U908 ( .A0(n484), .A1(n467), .B0(n1163), .B1(n483), .Y(n489) );
  OAI22XL U909 ( .A0(n1098), .A1(n471), .B0(n1127), .B1(n486), .Y(n491) );
  XNOR2X1 U910 ( .A(n833), .B(B[24]), .Y(n507) );
  XNOR2X1 U911 ( .A(n1118), .B(n783), .Y(n509) );
  OAI22XL U912 ( .A0(n1147), .A1(n509), .B0(n1148), .B1(n474), .Y(n512) );
  CMPR32X1 U913 ( .A(n478), .B(n477), .C(n476), .CO(n495), .S(n521) );
  CMPR32X1 U914 ( .A(n481), .B(n480), .C(n479), .CO(n525), .S(n520) );
  XNOR2X1 U915 ( .A(A[15]), .B(B[20]), .Y(n1073) );
  OAI22X1 U916 ( .A0(n1076), .A1(n485), .B0(n1077), .B1(n1074), .Y(n1093) );
  CMPR32X1 U917 ( .A(n489), .B(n488), .C(n487), .CO(n1085), .S(n494) );
  CMPR32X1 U918 ( .A(n492), .B(n491), .C(n490), .CO(n1084), .S(n493) );
  CMPR32X1 U919 ( .A(n495), .B(n494), .C(n493), .CO(n1070), .S(n524) );
  NOR2XL U920 ( .A(n497), .B(n496), .Y(mult_x_1_n162) );
  NAND2XL U921 ( .A(n497), .B(n496), .Y(mult_x_1_n163) );
  NAND2XL U922 ( .A(n528), .B(n442), .Y(n501) );
  AOI21XL U923 ( .A0(n566), .A1(n442), .B0(n444), .Y(n500) );
  OAI21XL U924 ( .A0(n1215), .A1(n501), .B0(n500), .Y(n504) );
  INVXL U925 ( .A(n515), .Y(n539) );
  OAI22XL U926 ( .A0(n1135), .A1(n543), .B0(n1148), .B1(n509), .Y(n537) );
  CMPR32X1 U927 ( .A(n513), .B(n512), .C(n511), .CO(n522), .S(n560) );
  CMPR32X1 U928 ( .A(n516), .B(n515), .C(n514), .CO(n479), .S(n559) );
  ADDFHX1 U929 ( .A(n519), .B(n518), .CI(n517), .CO(n563), .S(n558) );
  CMPR32X1 U930 ( .A(n522), .B(n521), .C(n520), .CO(n523), .S(n561) );
  CMPR32X1 U931 ( .A(n525), .B(n524), .C(n523), .CO(n497), .S(n526) );
  NOR2XL U932 ( .A(n527), .B(n526), .Y(mult_x_1_n173) );
  NAND2XL U933 ( .A(n527), .B(n526), .Y(mult_x_1_n174) );
  NAND2XL U934 ( .A(n528), .B(n568), .Y(n530) );
  INVXL U935 ( .A(n1235), .Y(n529) );
  XNOR2X2 U936 ( .A(n533), .B(n532), .Y(PRODUCT[32]) );
  XNOR2X1 U937 ( .A(n1161), .B(B[14]), .Y(n550) );
  OAI22XL U938 ( .A0(n1165), .A1(n550), .B0(n1163), .B1(n534), .Y(n554) );
  XNOR2X1 U939 ( .A(A[3]), .B(B[25]), .Y(n586) );
  CMPR32X1 U940 ( .A(n538), .B(n537), .C(n536), .CO(n517), .S(n575) );
  CMPR32X1 U941 ( .A(n541), .B(n540), .C(n539), .CO(n518), .S(n574) );
  XNOR2X1 U942 ( .A(n462), .B(B[24]), .Y(n548) );
  OAI22XL U943 ( .A0(n875), .A1(n548), .B0(n873), .B1(n542), .Y(n557) );
  OAI22XL U944 ( .A0(n1147), .A1(n577), .B0(n1148), .B1(n543), .Y(n556) );
  OAI22XL U945 ( .A0(n1076), .A1(n551), .B0(n1077), .B1(n545), .Y(n585) );
  XNOR2X1 U946 ( .A(n1078), .B(n783), .Y(n547) );
  OAI22XL U947 ( .A0(n1098), .A1(n547), .B0(n1127), .B1(n546), .Y(n584) );
  XNOR2X1 U948 ( .A(n1078), .B(n825), .Y(n587) );
  XNOR2X1 U949 ( .A(n462), .B(B[23]), .Y(n588) );
  INVXL U950 ( .A(n553), .Y(n589) );
  XNOR2X1 U951 ( .A(n1161), .B(B[13]), .Y(n580) );
  CMPR32X1 U952 ( .A(n557), .B(n556), .C(n555), .CO(n596), .S(n609) );
  CMPR32X1 U953 ( .A(n563), .B(n562), .C(n561), .CO(n527), .S(n564) );
  NOR2XL U954 ( .A(n565), .B(n564), .Y(mult_x_1_n184) );
  NAND2XL U955 ( .A(n565), .B(n564), .Y(mult_x_1_n185) );
  CMPR32X1 U956 ( .A(n576), .B(n575), .C(n574), .CO(n573), .S(n608) );
  XNOR2X1 U957 ( .A(n1118), .B(B[15]), .Y(n579) );
  OAI22XL U958 ( .A0(n1135), .A1(n618), .B0(n1148), .B1(n579), .Y(n614) );
  OR2X1 U959 ( .A(n615), .B(n614), .Y(n620) );
  XNOR2X1 U960 ( .A(n823), .B(n783), .Y(n616) );
  XNOR2X1 U961 ( .A(n1161), .B(B[12]), .Y(n613) );
  XNOR2X1 U962 ( .A(n581), .B(n1160), .Y(n612) );
  INVXL U963 ( .A(n612), .Y(n582) );
  CMPR32X1 U964 ( .A(n585), .B(n584), .C(n583), .CO(n595), .S(n632) );
  OAI22X1 U965 ( .A0(n1126), .A1(n623), .B0(n1127), .B1(n587), .Y(n629) );
  XNOR2X1 U966 ( .A(n462), .B(B[22]), .Y(n622) );
  OAI22XL U967 ( .A0(n875), .A1(n622), .B0(n873), .B1(n588), .Y(n628) );
  NAND2X1 U968 ( .A(n603), .B(n1237), .Y(n604) );
  CMPR32X1 U969 ( .A(n608), .B(n607), .C(n606), .CO(n597), .S(n635) );
  CMPR32X1 U970 ( .A(n611), .B(n610), .C(n609), .CO(n594), .S(n643) );
  XNOR2X1 U971 ( .A(n581), .B(B[25]), .Y(n649) );
  OAI22XL U972 ( .A0(n1165), .A1(n650), .B0(n1163), .B1(n613), .Y(n647) );
  XNOR2X1 U973 ( .A(n823), .B(n825), .Y(n651) );
  OAI22X1 U974 ( .A0(n866), .A1(n652), .B0(n864), .B1(n617), .Y(n661) );
  XNOR2X1 U975 ( .A(A[13]), .B(B[13]), .Y(n653) );
  XNOR2X1 U976 ( .A(n1078), .B(B[15]), .Y(n658) );
  OAI22XL U977 ( .A0(n881), .A1(n659), .B0(n879), .B1(n624), .Y(n663) );
  ADDFHX1 U978 ( .A(n630), .B(n629), .CI(n628), .CO(n646), .S(n677) );
  NOR2XL U979 ( .A(n635), .B(n634), .Y(mult_x_1_n202) );
  NAND2XL U980 ( .A(n635), .B(n634), .Y(mult_x_1_n203) );
  NAND2X1 U981 ( .A(n638), .B(n1239), .Y(n639) );
  CMPR32X1 U982 ( .A(n643), .B(n642), .C(n641), .CO(n634), .S(n670) );
  CMPR32X1 U983 ( .A(n646), .B(n645), .C(n644), .CO(n631), .S(n676) );
  ADDHXL U984 ( .A(n648), .B(n647), .CO(n656), .S(n689) );
  XNOR2X1 U985 ( .A(n581), .B(B[24]), .Y(n682) );
  OAI22X1 U986 ( .A0(n859), .A1(n682), .B0(n649), .B1(n1064), .Y(n681) );
  XNOR2X1 U987 ( .A(n1161), .B(n788), .Y(n683) );
  XNOR2X1 U988 ( .A(n823), .B(B[16]), .Y(n684) );
  XNOR2X1 U989 ( .A(A[3]), .B(B[22]), .Y(n685) );
  OAI22X1 U990 ( .A0(n866), .A1(n685), .B0(n864), .B1(n652), .Y(n694) );
  XNOR2X1 U991 ( .A(A[13]), .B(B[12]), .Y(n686) );
  ADDFHX1 U992 ( .A(n656), .B(n655), .CI(n654), .CO(n668), .S(n700) );
  XNOR2X1 U993 ( .A(A[11]), .B(B[14]), .Y(n691) );
  OAI22XL U994 ( .A0(n881), .A1(n692), .B0(n879), .B1(n659), .Y(n696) );
  NOR2XL U995 ( .A(n670), .B(n669), .Y(mult_x_1_n209) );
  NAND2XL U996 ( .A(n670), .B(n669), .Y(mult_x_1_n210) );
  INVXL U997 ( .A(n1240), .Y(n671) );
  NAND2X1 U998 ( .A(n671), .B(n1241), .Y(n672) );
  CMPR32X1 U999 ( .A(n676), .B(n675), .C(n674), .CO(n669), .S(n703) );
  CMPR32X1 U1000 ( .A(n679), .B(n678), .C(n677), .CO(n666), .S(n708) );
  CMPR22X1 U1001 ( .A(n681), .B(n680), .CO(n688), .S(n720) );
  XNOR2X1 U1002 ( .A(n581), .B(B[23]), .Y(n714) );
  OAI22X1 U1003 ( .A0(n859), .A1(n714), .B0(n682), .B1(n1064), .Y(n713) );
  XNOR2X1 U1004 ( .A(n823), .B(B[15]), .Y(n716) );
  OAI22XL U1005 ( .A0(n1076), .A1(n716), .B0(n1077), .B1(n684), .Y(n726) );
  ADDFHX1 U1006 ( .A(n689), .B(n688), .CI(n687), .CO(n701), .S(n731) );
  XNOR2X1 U1007 ( .A(A[11]), .B(B[13]), .Y(n722) );
  OAI22XL U1008 ( .A0(n791), .A1(n723), .B0(n879), .B1(n692), .Y(n727) );
  NOR2XL U1009 ( .A(n703), .B(n702), .Y(mult_x_1_n220) );
  NAND2XL U1010 ( .A(n703), .B(n702), .Y(mult_x_1_n221) );
  CMPR32X1 U1011 ( .A(n708), .B(n707), .C(n706), .CO(n702), .S(n734) );
  CMPR32X1 U1012 ( .A(n711), .B(n710), .C(n709), .CO(n699), .S(n741) );
  CMPR22X1 U1013 ( .A(n713), .B(n712), .CO(n719), .S(n755) );
  XNOR2X1 U1014 ( .A(n581), .B(B[22]), .Y(n748) );
  OAI22X1 U1015 ( .A0(n859), .A1(n748), .B0(n714), .B1(n1064), .Y(n746) );
  XNOR2X1 U1016 ( .A(n1161), .B(B[8]), .Y(n749) );
  XNOR2X1 U1017 ( .A(n823), .B(B[14]), .Y(n750) );
  OAI22XL U1018 ( .A0(n1076), .A1(n750), .B0(n1077), .B1(n716), .Y(n760) );
  OAI22XL U1019 ( .A0(n791), .A1(n757), .B0(n879), .B1(n723), .Y(n761) );
  CMPR32X1 U1020 ( .A(n726), .B(n725), .C(n724), .CO(n718), .S(n776) );
  NOR2XL U1021 ( .A(n734), .B(n733), .Y(mult_x_1_n223) );
  NAND2XL U1022 ( .A(n734), .B(n733), .Y(mult_x_1_n224) );
  CMPR32X1 U1023 ( .A(n744), .B(n743), .C(n742), .CO(n730), .S(n774) );
  CMPR22X1 U1024 ( .A(n746), .B(n745), .CO(n754), .S(n787) );
  XNOR2X1 U1025 ( .A(n581), .B(B[21]), .Y(n780) );
  OAI22X1 U1026 ( .A0(n859), .A1(n780), .B0(n748), .B1(n747), .Y(n779) );
  XNOR2X1 U1027 ( .A(n1161), .B(n826), .Y(n781) );
  XNOR2X1 U1028 ( .A(n823), .B(B[13]), .Y(n782) );
  OAI22XL U1029 ( .A0(n1076), .A1(n782), .B0(n1077), .B1(n750), .Y(n794) );
  XNOR2X1 U1030 ( .A(A[13]), .B(B[9]), .Y(n784) );
  OAI22X1 U1031 ( .A0(n1098), .A1(n789), .B0(n1127), .B1(n756), .Y(n796) );
  CMPR32X1 U1032 ( .A(n760), .B(n759), .C(n758), .CO(n753), .S(n814) );
  ADDFHX1 U1033 ( .A(n766), .B(n765), .CI(n764), .CO(n740), .S(n772) );
  NAND2XL U1034 ( .A(n768), .B(n767), .Y(mult_x_1_n233) );
  CMPR32X1 U1035 ( .A(n774), .B(n773), .C(n772), .CO(n767), .S(n802) );
  CMPR32X1 U1036 ( .A(n777), .B(n776), .C(n775), .CO(n764), .S(n812) );
  CMPR22X1 U1037 ( .A(n779), .B(n778), .CO(n786), .S(n830) );
  OAI22X1 U1038 ( .A0(n820), .A1(n819), .B0(n780), .B1(n1064), .Y(n817) );
  XNOR2X1 U1039 ( .A(n1161), .B(B[6]), .Y(n822) );
  XNOR2X1 U1040 ( .A(n823), .B(B[12]), .Y(n824) );
  OAI22XL U1041 ( .A0(n1076), .A1(n824), .B0(n1077), .B1(n782), .Y(n837) );
  XNOR2X1 U1042 ( .A(A[13]), .B(B[8]), .Y(n827) );
  XNOR2X1 U1043 ( .A(A[11]), .B(n788), .Y(n832) );
  CMPR32X1 U1044 ( .A(n794), .B(n793), .C(n792), .CO(n785), .S(n855) );
  NOR2XL U1045 ( .A(n802), .B(n801), .Y(mult_x_1_n241) );
  NAND2XL U1046 ( .A(n803), .B(n848), .Y(n806) );
  OAI21XL U1047 ( .A0(n953), .A1(n806), .B0(n805), .Y(n809) );
  CMPR32X1 U1048 ( .A(n815), .B(n814), .C(n813), .CO(n798), .S(n853) );
  CMPR22X1 U1049 ( .A(n817), .B(n816), .CO(n829), .S(n871) );
  OAI22X1 U1050 ( .A0(n1165), .A1(n860), .B0(n1163), .B1(n822), .Y(n857) );
  XNOR2X1 U1051 ( .A(A[13]), .B(n826), .Y(n867) );
  XNOR2X1 U1052 ( .A(n462), .B(B[15]), .Y(n872) );
  OAI22XL U1053 ( .A0(n875), .A1(n872), .B0(n873), .B1(n831), .Y(n887) );
  XNOR2X1 U1054 ( .A(A[11]), .B(B[9]), .Y(n876) );
  OAI22XL U1055 ( .A0(n1098), .A1(n876), .B0(n1127), .B1(n832), .Y(n886) );
  CMPR32X1 U1056 ( .A(n837), .B(n836), .C(n835), .CO(n828), .S(n902) );
  NOR2XL U1057 ( .A(n845), .B(n844), .Y(mult_x_1_n252) );
  NAND2XL U1058 ( .A(n845), .B(n844), .Y(mult_x_1_n253) );
  NAND2X1 U1059 ( .A(n848), .B(n1251), .Y(n849) );
  CMPR32X1 U1060 ( .A(n853), .B(n852), .C(n851), .CO(n844), .S(n892) );
  CMPR32X1 U1061 ( .A(n856), .B(n855), .C(n854), .CO(n841), .S(n900) );
  OAI22XL U1062 ( .A0(n1076), .A1(n863), .B0(n1077), .B1(n862), .Y(n919) );
  OAI22XL U1063 ( .A0(n1098), .A1(n877), .B0(n1127), .B1(n876), .Y(n921) );
  ADDFHX1 U1064 ( .A(n884), .B(n883), .CI(n882), .CO(n869), .S(n937) );
  CMPR32X1 U1065 ( .A(n887), .B(n886), .C(n885), .CO(n903), .S(n936) );
  NOR2XL U1066 ( .A(n892), .B(n891), .Y(mult_x_1_n259) );
  NAND2XL U1067 ( .A(n892), .B(n891), .Y(mult_x_1_n260) );
  INVX1 U1068 ( .A(n1254), .Y(n932) );
  NAND2XL U1069 ( .A(n928), .B(n932), .Y(n895) );
  INVXL U1070 ( .A(n1255), .Y(n893) );
  INVXL U1071 ( .A(n1252), .Y(n896) );
  CMPR32X1 U1072 ( .A(n903), .B(n902), .C(n901), .CO(n888), .S(n935) );
  CMPR22X1 U1073 ( .A(n905), .B(n904), .CO(n912), .S(n944) );
  CMPR22X1 U1074 ( .A(n907), .B(n906), .CO(n943), .S(n941) );
  CMPR32X1 U1075 ( .A(n910), .B(n909), .C(n908), .CO(n942), .S(n946) );
  CMPR32X1 U1076 ( .A(n916), .B(n915), .C(n914), .CO(n961), .S(n945) );
  CMPR32X1 U1077 ( .A(n922), .B(n921), .C(n920), .CO(n938), .S(n959) );
  CMPR32X1 U1078 ( .A(n925), .B(n924), .C(n923), .CO(n899), .S(n933) );
  NOR2XL U1079 ( .A(n927), .B(n926), .Y(mult_x_1_n270) );
  NAND2XL U1080 ( .A(n927), .B(n926), .Y(mult_x_1_n271) );
  INVXL U1081 ( .A(n928), .Y(n931) );
  INVXL U1082 ( .A(n929), .Y(n930) );
  CMPR32X1 U1083 ( .A(n935), .B(n934), .C(n933), .CO(n926), .S(n952) );
  CMPR32X1 U1084 ( .A(n938), .B(n937), .C(n936), .CO(n923), .S(n958) );
  CMPR32X1 U1085 ( .A(n941), .B(n940), .C(n939), .CO(n967), .S(n963) );
  CMPR32X1 U1086 ( .A(n947), .B(n946), .C(n945), .CO(n965), .S(n975) );
  NOR2XL U1087 ( .A(n952), .B(n951), .Y(mult_x_1_n277) );
  INVXL U1088 ( .A(n1256), .Y(n954) );
  CMPR32X1 U1089 ( .A(n961), .B(n960), .C(n959), .CO(n948), .S(n972) );
  CMPR32X1 U1090 ( .A(n964), .B(n963), .C(n962), .CO(n971), .S(n973) );
  NOR2XL U1091 ( .A(n969), .B(n968), .Y(mult_x_1_n288) );
  NAND2XL U1092 ( .A(n977), .B(n976), .Y(mult_x_1_n292) );
  OAI21XL U1093 ( .A0(n986), .A1(n1263), .B0(n1264), .Y(n981) );
  NAND2X1 U1094 ( .A(n979), .B(n1262), .Y(n980) );
  XNOR2X2 U1095 ( .A(n981), .B(n980), .Y(PRODUCT[18]) );
  NAND2XL U1096 ( .A(n983), .B(n982), .Y(mult_x_1_n300) );
  INVXL U1097 ( .A(n1263), .Y(n984) );
  NAND2X1 U1098 ( .A(n984), .B(n1264), .Y(n985) );
  NAND2XL U1099 ( .A(n988), .B(n987), .Y(mult_x_1_n303) );
  INVXL U1100 ( .A(n1268), .Y(n989) );
  NOR2XL U1101 ( .A(n992), .B(mult_x_1_n312), .Y(mult_x_1_n305) );
  INVXL U1102 ( .A(n992), .Y(n994) );
  NAND2XL U1103 ( .A(n994), .B(n993), .Y(mult_x_1_n78) );
  NAND2XL U1104 ( .A(n995), .B(n1268), .Y(n996) );
  CMPR32X1 U1105 ( .A(n1002), .B(n1001), .C(n1000), .CO(n1020), .S(n1015) );
  CMPR32X1 U1106 ( .A(n1008), .B(n1007), .C(n1006), .CO(n997), .S(n1018) );
  CMPR32X1 U1107 ( .A(n1011), .B(n1010), .C(n1009), .CO(n1029), .S(n1031) );
  CMPR32X1 U1108 ( .A(n1014), .B(n1013), .C(n1012), .CO(n1009), .S(n1023) );
  CMPR32X1 U1109 ( .A(n1020), .B(n1019), .C(n1018), .CO(n1032), .S(n1021) );
  CMPR32X1 U1110 ( .A(n1023), .B(n1022), .C(n1021), .CO(n1036), .S(n1035) );
  NOR2XL U1111 ( .A(n1045), .B(n1041), .Y(mult_x_1_n316) );
  INVXL U1112 ( .A(n1046), .Y(n1049) );
  NAND2XL U1113 ( .A(n1037), .B(n1036), .Y(n1069) );
  INVXL U1114 ( .A(n1069), .Y(n1038) );
  OAI21XL U1115 ( .A0(n1044), .A1(n1041), .B0(n1042), .Y(mult_x_1_n317) );
  INVXL U1116 ( .A(n1041), .Y(n1043) );
  NAND2XL U1117 ( .A(n1043), .B(n1042), .Y(mult_x_1_n80) );
  XNOR2X1 U1118 ( .A(n1275), .B(n1271), .Y(PRODUCT[13]) );
  NAND2XL U1119 ( .A(n1048), .B(n1046), .Y(n1047) );
  XOR2X1 U1120 ( .A(n1050), .B(n1047), .Y(n1290) );
  OAI21XL U1121 ( .A0(n1050), .A1(n1027), .B0(n1046), .Y(mult_x_1_n327) );
  AOI21XL U1122 ( .A0(n1058), .A1(n1056), .B0(n1051), .Y(n1054) );
  NAND2XL U1123 ( .A(n62), .B(n1052), .Y(n1053) );
  XOR2X1 U1124 ( .A(n1054), .B(n1053), .Y(n1291) );
  NAND2XL U1125 ( .A(n1056), .B(n1055), .Y(n1057) );
  XNOR2X1 U1126 ( .A(n1058), .B(n1057), .Y(n1292) );
  INVXL U1127 ( .A(n1059), .Y(n1175) );
  OAI21XL U1128 ( .A0(n1175), .A1(n1171), .B0(n1172), .Y(n1063) );
  NAND2XL U1129 ( .A(n84), .B(n1061), .Y(n1062) );
  OAI21XL U1130 ( .A0(n1215), .A1(n1066), .B0(n1065), .Y(n1068) );
  NAND2XL U1131 ( .A(n58), .B(n1069), .Y(mult_x_1_n81) );
  CMPR32X1 U1132 ( .A(n1083), .B(n1082), .C(n1081), .CO(n1099), .S(n1072) );
  CMPR32X1 U1133 ( .A(n1086), .B(n1085), .C(n1084), .CO(n1089), .S(n1071) );
  CMPR32X1 U1134 ( .A(n1091), .B(n1090), .C(n1089), .CO(n1103), .S(n1087) );
  CMPR32X1 U1135 ( .A(n1094), .B(n1093), .C(n1092), .CO(n1117), .S(n1091) );
  XNOR2X1 U1136 ( .A(A[11]), .B(n1160), .Y(n1124) );
  OAI22X1 U1137 ( .A0(n1098), .A1(n1097), .B0(n1127), .B1(n1124), .Y(n1138) );
  CMPR32X1 U1138 ( .A(n1101), .B(n1100), .C(n1099), .CO(n1115), .S(n1090) );
  OAI21XL U1139 ( .A0(n1215), .A1(n1111), .B0(n1110), .Y(n1114) );
  CMPR32X1 U1140 ( .A(n1117), .B(n1116), .C(n1115), .CO(n1129), .S(n1102) );
  CMPR32X1 U1141 ( .A(n1122), .B(n1121), .C(n1120), .CO(n1131), .S(n1116) );
  XNOR2X1 U1142 ( .A(A[15]), .B(B[23]), .Y(n1133) );
  CMPR32X1 U1143 ( .A(n1132), .B(n1131), .C(n1130), .CO(n1140), .S(n1128) );
  XNOR2X1 U1144 ( .A(A[15]), .B(B[24]), .Y(n1144) );
  OAI22X1 U1145 ( .A0(n1135), .A1(n1134), .B0(n1148), .B1(n1145), .Y(n1159) );
  CMPR32X1 U1146 ( .A(n1138), .B(n1137), .C(n1136), .CO(n1141), .S(n1130) );
  CMPR32X1 U1147 ( .A(n1143), .B(n1142), .C(n1141), .CO(n1150), .S(n1139) );
  XNOR2X1 U1148 ( .A(A[15]), .B(B[25]), .Y(n1164) );
  OAI21XL U1149 ( .A0(n1152), .A1(n1220), .B0(n1221), .Y(n1208) );
  OAI21XL U1150 ( .A0(n1215), .A1(n1154), .B0(n1153), .Y(n1156) );
  CMPR32X1 U1151 ( .A(n1159), .B(n1158), .C(n1157), .CO(n1168), .S(n1149) );
  XNOR2XL U1152 ( .A(n1161), .B(n1160), .Y(n1162) );
  INVXL U1153 ( .A(n1171), .Y(n1173) );
  NAND2XL U1154 ( .A(n1173), .B(n1172), .Y(n1174) );
  XNOR2XL U1155 ( .A(n1204), .B(n1203), .Y(n1297) );
  AOI21XL U1156 ( .A0(n1212), .A1(n1211), .B0(n1210), .Y(n1213) );
  OAI21XL U1157 ( .A0(n1215), .A1(n1214), .B0(n1213), .Y(n1216) );
endmodule


module FFT2048_DW02_mult_2_stage_J1_15 ( A, B, TC, CLK, PRODUCT );
  input [15:0] A;
  input [26:0] B;
  output [42:0] PRODUCT;
  input TC, CLK;
  wire   n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, mult_x_1_n327, mult_x_1_n320, mult_x_1_n315,
         mult_x_1_n313, mult_x_1_n312, mult_x_1_n306, mult_x_1_n305,
         mult_x_1_n303, mult_x_1_n302, mult_x_1_n300, mult_x_1_n299,
         mult_x_1_n297, mult_x_1_n292, mult_x_1_n291, mult_x_1_n289,
         mult_x_1_n288, mult_x_1_n278, mult_x_1_n277, mult_x_1_n271,
         mult_x_1_n270, mult_x_1_n260, mult_x_1_n259, mult_x_1_n253,
         mult_x_1_n252, mult_x_1_n242, mult_x_1_n241, mult_x_1_n233,
         mult_x_1_n232, mult_x_1_n224, mult_x_1_n223, mult_x_1_n221,
         mult_x_1_n220, mult_x_1_n210, mult_x_1_n209, mult_x_1_n203,
         mult_x_1_n202, mult_x_1_n192, mult_x_1_n191, mult_x_1_n185,
         mult_x_1_n184, mult_x_1_n174, mult_x_1_n173, mult_x_1_n163,
         mult_x_1_n162, mult_x_1_n150, mult_x_1_n149, mult_x_1_n135,
         mult_x_1_n134, mult_x_1_n126, mult_x_1_n125, mult_x_1_n115,
         mult_x_1_n114, mult_x_1_n106, mult_x_1_n105, mult_x_1_n81,
         mult_x_1_n80, mult_x_1_n78, mult_x_1_n54, n5, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257;

  DFFHQXL mult_x_1_clk_r_REG40_S1 ( .D(mult_x_1_n173), .CK(CLK), .Q(n1213) );
  DFFHQX1 mult_x_1_clk_r_REG6_S1 ( .D(mult_x_1_n302), .CK(CLK), .Q(n1246) );
  DFFHQXL mult_x_1_clk_r_REG24_S1 ( .D(mult_x_1_n209), .CK(CLK), .Q(n1221) );
  DFFHQXL mult_x_1_clk_r_REG36_S1 ( .D(mult_x_1_n191), .CK(CLK), .Q(n1217) );
  DFFHQX4 mult_x_1_clk_r_REG54_S1 ( .D(mult_x_1_n315), .CK(CLK), .Q(n1255) );
  DFFHQX4 mult_x_1_clk_r_REG5_S1 ( .D(mult_x_1_n303), .CK(CLK), .Q(n1247) );
  DFFHQX4 mult_x_1_clk_r_REG10_S1 ( .D(mult_x_1_n292), .CK(CLK), .Q(n1242) );
  DFFHQX4 mult_x_1_clk_r_REG32_S1 ( .D(mult_x_1_n288), .CK(CLK), .Q(n1239) );
  DFFHQX4 mult_x_1_clk_r_REG29_S1 ( .D(mult_x_1_n278), .CK(CLK), .Q(n1238) );
  DFFHQX4 mult_x_1_clk_r_REG28_S1 ( .D(mult_x_1_n270), .CK(CLK), .Q(n1235) );
  DFFHQX4 mult_x_1_clk_r_REG14_S1 ( .D(mult_x_1_n252), .CK(CLK), .Q(n1231) );
  DFFHQX4 mult_x_1_clk_r_REG16_S1 ( .D(mult_x_1_n241), .CK(CLK), .Q(n1229) );
  DFFHQX4 mult_x_1_clk_r_REG18_S1 ( .D(mult_x_1_n232), .CK(CLK), .Q(n1227) );
  DFFHQXL clk_r_REG57_S1 ( .D(n1272), .CK(CLK), .Q(PRODUCT[12]) );
  DFFHQXL mult_x_1_clk_r_REG20_S1 ( .D(mult_x_1_n223), .CK(CLK), .Q(n1225) );
  DFFHQXL mult_x_1_clk_r_REG37_S1 ( .D(mult_x_1_n185), .CK(CLK), .Q(n1216) );
  DFFHQX4 mult_x_1_clk_r_REG13_S1 ( .D(mult_x_1_n253), .CK(CLK), .Q(n1232) );
  DFFHQX4 mult_x_1_clk_r_REG27_S1 ( .D(mult_x_1_n271), .CK(CLK), .Q(n1236) );
  DFFHQXL mult_x_1_clk_r_REG22_S1 ( .D(mult_x_1_n220), .CK(CLK), .Q(n1223) );
  DFFHQXL mult_x_1_clk_r_REG35_S1 ( .D(mult_x_1_n192), .CK(CLK), .Q(n1218) );
  DFFHQXL clk_r_REG59_S1 ( .D(n1273), .CK(CLK), .Q(PRODUCT[11]) );
  DFFHQXL clk_r_REG60_S1 ( .D(n1274), .CK(CLK), .Q(PRODUCT[10]) );
  DFFHQXL mult_x_1_clk_r_REG42_S1 ( .D(mult_x_1_n162), .CK(CLK), .Q(n1211) );
  DFFHQXL mult_x_1_clk_r_REG38_S1 ( .D(mult_x_1_n184), .CK(CLK), .Q(n1215) );
  DFFHQXL mult_x_1_clk_r_REG41_S1 ( .D(mult_x_1_n163), .CK(CLK), .Q(n1212) );
  DFFHQXL clk_r_REG70_S1 ( .D(n1284), .CK(CLK), .Q(PRODUCT[0]) );
  DFFHQXL mult_x_1_clk_r_REG21_S1 ( .D(mult_x_1_n221), .CK(CLK), .Q(n1224) );
  DFFHQXL mult_x_1_clk_r_REG12_S1 ( .D(mult_x_1_n54), .CK(CLK), .Q(n1200) );
  DFFHQX4 mult_x_1_clk_r_REG31_S1 ( .D(mult_x_1_n289), .CK(CLK), .Q(n1240) );
  DFFHQX4 mult_x_1_clk_r_REG1_S1 ( .D(mult_x_1_n306), .CK(CLK), .Q(n1254) );
  DFFHQXL mult_x_1_clk_r_REG39_S1 ( .D(mult_x_1_n174), .CK(CLK), .Q(n1214) );
  DFFHQXL clk_r_REG61_S1 ( .D(n1275), .CK(CLK), .Q(PRODUCT[9]) );
  DFFHQXL clk_r_REG62_S1 ( .D(n1276), .CK(CLK), .Q(PRODUCT[8]) );
  DFFHQXL clk_r_REG63_S1 ( .D(n1277), .CK(CLK), .Q(PRODUCT[7]) );
  DFFHQXL clk_r_REG64_S1 ( .D(n1278), .CK(CLK), .Q(PRODUCT[6]) );
  DFFHQXL clk_r_REG65_S1 ( .D(n1279), .CK(CLK), .Q(PRODUCT[5]) );
  DFFHQXL clk_r_REG66_S1 ( .D(n1280), .CK(CLK), .Q(PRODUCT[4]) );
  DFFHQXL clk_r_REG67_S1 ( .D(n1281), .CK(CLK), .Q(PRODUCT[3]) );
  DFFHQXL clk_r_REG68_S1 ( .D(n1282), .CK(CLK), .Q(PRODUCT[2]) );
  DFFHQXL clk_r_REG69_S1 ( .D(n1283), .CK(CLK), .Q(PRODUCT[1]) );
  DFFHQX2 mult_x_1_clk_r_REG2_S1 ( .D(mult_x_1_n312), .CK(CLK), .Q(n1250) );
  DFFHQXL mult_x_1_clk_r_REG55_S1 ( .D(mult_x_1_n81), .CK(CLK), .Q(n1253) );
  DFFHQXL mult_x_1_clk_r_REG4_S1 ( .D(mult_x_1_n78), .CK(CLK), .Q(n1249) );
  DFFHQXL mult_x_1_clk_r_REG23_S1 ( .D(mult_x_1_n210), .CK(CLK), .Q(n1222) );
  DFFHQXL mult_x_1_clk_r_REG33_S1 ( .D(mult_x_1_n203), .CK(CLK), .Q(n1220) );
  DFFHQXL mult_x_1_clk_r_REG43_S1 ( .D(mult_x_1_n150), .CK(CLK), .Q(n1210) );
  DFFHQXL mult_x_1_clk_r_REG44_S1 ( .D(mult_x_1_n149), .CK(CLK), .Q(n1209) );
  DFFHQXL mult_x_1_clk_r_REG45_S1 ( .D(mult_x_1_n135), .CK(CLK), .Q(n1208) );
  DFFHQXL mult_x_1_clk_r_REG46_S1 ( .D(mult_x_1_n134), .CK(CLK), .Q(n1207) );
  DFFHQXL mult_x_1_clk_r_REG47_S1 ( .D(mult_x_1_n126), .CK(CLK), .Q(n1206) );
  DFFHQXL mult_x_1_clk_r_REG48_S1 ( .D(mult_x_1_n125), .CK(CLK), .Q(n1205) );
  DFFHQXL mult_x_1_clk_r_REG49_S1 ( .D(mult_x_1_n115), .CK(CLK), .Q(n1204) );
  DFFHQXL mult_x_1_clk_r_REG50_S1 ( .D(mult_x_1_n114), .CK(CLK), .Q(n1203) );
  DFFHQXL mult_x_1_clk_r_REG51_S1 ( .D(mult_x_1_n106), .CK(CLK), .Q(n1202) );
  DFFHQXL mult_x_1_clk_r_REG52_S1 ( .D(mult_x_1_n105), .CK(CLK), .Q(n1201) );
  DFFHQXL mult_x_1_clk_r_REG34_S1 ( .D(mult_x_1_n202), .CK(CLK), .Q(n1219) );
  DFFHQX1 mult_x_1_clk_r_REG56_S1 ( .D(mult_x_1_n320), .CK(CLK), .Q(n1256) );
  DFFHQX1 mult_x_1_clk_r_REG0_S1 ( .D(mult_x_1_n313), .CK(CLK), .Q(n1251) );
  DFFHQXL mult_x_1_clk_r_REG58_S1 ( .D(mult_x_1_n327), .CK(CLK), .Q(n1257) );
  DFFHQX1 mult_x_1_clk_r_REG11_S1 ( .D(mult_x_1_n291), .CK(CLK), .Q(n1241) );
  DFFHQXL mult_x_1_clk_r_REG53_S1 ( .D(mult_x_1_n80), .CK(CLK), .Q(n1252) );
  DFFHQX2 mult_x_1_clk_r_REG30_S1 ( .D(mult_x_1_n277), .CK(CLK), .Q(n1237) );
  DFFHQX1 mult_x_1_clk_r_REG25_S1 ( .D(mult_x_1_n260), .CK(CLK), .Q(n1234) );
  DFFHQX1 mult_x_1_clk_r_REG9_S1 ( .D(mult_x_1_n299), .CK(CLK), .Q(n1244) );
  DFFHQX2 mult_x_1_clk_r_REG26_S1 ( .D(mult_x_1_n259), .CK(CLK), .Q(n1233) );
  DFFHQX2 mult_x_1_clk_r_REG7_S1 ( .D(mult_x_1_n297), .CK(CLK), .Q(n1243) );
  DFFHQX2 mult_x_1_clk_r_REG3_S1 ( .D(mult_x_1_n305), .CK(CLK), .Q(n1248) );
  DFFHQX1 mult_x_1_clk_r_REG17_S1 ( .D(mult_x_1_n233), .CK(CLK), .Q(n1228) );
  DFFHQX1 mult_x_1_clk_r_REG15_S1 ( .D(mult_x_1_n242), .CK(CLK), .Q(n1230) );
  DFFHQX1 mult_x_1_clk_r_REG19_S1 ( .D(mult_x_1_n224), .CK(CLK), .Q(n1226) );
  DFFHQX1 mult_x_1_clk_r_REG8_S1 ( .D(mult_x_1_n300), .CK(CLK), .Q(n1245) );
  ADDFHX1 U1 ( .A(n527), .B(n526), .CI(n525), .CO(n512), .S(n557) );
  ADDFHX1 U2 ( .A(n480), .B(n479), .CI(n478), .CO(n454), .S(n485) );
  ADDFHX1 U3 ( .A(n447), .B(n446), .CI(n445), .CO(n422), .S(n453) );
  ADDFHX1 U4 ( .A(n810), .B(n809), .CI(n808), .CO(n793), .S(n815) );
  ADDFHX1 U5 ( .A(n813), .B(n812), .CI(n811), .CO(n814), .S(n818) );
  ADDFHX1 U6 ( .A(n804), .B(n803), .CI(n802), .CO(n809), .S(n811) );
  ADDFX2 U7 ( .A(n771), .B(n770), .CI(n769), .CO(n745), .S(n775) );
  ADDFHX1 U8 ( .A(n376), .B(n375), .CI(n374), .CO(n351), .S(n386) );
  ADDFX2 U9 ( .A(n831), .B(n830), .CI(n829), .CO(n821), .S(n851) );
  ADDFHX1 U10 ( .A(n759), .B(n758), .CI(n757), .CO(n771), .S(n791) );
  CMPR32X1 U11 ( .A(n786), .B(n785), .C(n784), .CO(n792), .S(n803) );
  ADDFHX1 U12 ( .A(n586), .B(n585), .CI(n584), .CO(n602), .S(n634) );
  ADDFX2 U13 ( .A(n583), .B(n582), .CI(n581), .CO(n574), .S(n635) );
  CMPR32X1 U14 ( .A(n474), .B(n473), .C(n472), .CO(n466), .S(n529) );
  OAI22X1 U15 ( .A0(n577), .A1(n962), .B0(n37), .B1(n960), .Y(n586) );
  ADDFX2 U16 ( .A(n647), .B(n646), .CI(n645), .CO(n658), .S(n693) );
  OAI22X1 U17 ( .A0(n966), .A1(n365), .B0(n964), .B1(n315), .Y(n333) );
  XNOR2X2 U18 ( .A(B[22]), .B(n908), .Y(n464) );
  XOR2X1 U19 ( .A(B[18]), .B(n10), .Y(n675) );
  BUFX3 U20 ( .A(A[7]), .Y(n866) );
  BUFX3 U21 ( .A(A[3]), .Y(n908) );
  BUFX3 U22 ( .A(A[1]), .Y(n905) );
  XOR2X1 U23 ( .A(n64), .B(n349), .Y(PRODUCT[31]) );
  OAI21X1 U24 ( .A0(n225), .A1(n219), .B0(n32), .Y(n1195) );
  XOR2X2 U25 ( .A(n313), .B(n81), .Y(PRODUCT[32]) );
  OAI21XL U26 ( .A0(n1198), .A1(n347), .B0(n225), .Y(n64) );
  OAI21X1 U27 ( .A0(n95), .A1(n311), .B0(n310), .Y(n313) );
  OAI21XL U28 ( .A0(n95), .A1(n241), .B0(n240), .Y(n244) );
  XNOR2X2 U29 ( .A(n71), .B(n385), .Y(PRODUCT[30]) );
  XOR2X1 U30 ( .A(n61), .B(n743), .Y(PRODUCT[20]) );
  OAI21X1 U31 ( .A0(n1198), .A1(n383), .B0(n382), .Y(n71) );
  XNOR2X2 U32 ( .A(n702), .B(n701), .Y(PRODUCT[21]) );
  XOR2X2 U33 ( .A(n57), .B(n666), .Y(PRODUCT[22]) );
  NOR2BX1 U34 ( .AN(n663), .B(n58), .Y(n57) );
  OAI21X2 U35 ( .A0(n700), .A1(n73), .B0(n699), .Y(n702) );
  NOR2XL U36 ( .A(n1221), .B(n1219), .Y(n215) );
  NAND2X1 U37 ( .A(n35), .B(n1224), .Y(n380) );
  AOI21X2 U38 ( .A0(n215), .A1(n380), .B0(n214), .Y(n225) );
  OAI21X2 U39 ( .A0(n1242), .A1(n1239), .B0(n1240), .Y(n698) );
  AOI21XL U40 ( .A0(n628), .A1(n593), .B0(n592), .Y(n68) );
  AND2X1 U41 ( .A(n348), .B(n1218), .Y(n349) );
  AOI21XL U42 ( .A0(n828), .A1(n826), .B0(n819), .Y(n820) );
  XNOR2XL U43 ( .A(n1148), .B(B[9]), .Y(n493) );
  XNOR2XL U44 ( .A(n905), .B(n1147), .Y(n392) );
  XNOR2XL U45 ( .A(n1199), .B(n1200), .Y(PRODUCT[40]) );
  XNOR2XL U46 ( .A(n866), .B(n856), .Y(n135) );
  XNOR2XL U47 ( .A(n866), .B(n1147), .Y(n249) );
  XNOR2XL U48 ( .A(A[9]), .B(B[21]), .Y(n325) );
  XNOR2XL U49 ( .A(A[15]), .B(B[21]), .Y(n1080) );
  ADDFX2 U50 ( .A(n179), .B(n178), .CI(n177), .CO(n833), .S(n996) );
  OAI22X1 U51 ( .A0(n956), .A1(n287), .B0(n43), .B1(n958), .Y(n321) );
  ADDFX2 U52 ( .A(n334), .B(n333), .CI(n332), .CO(n355), .S(n390) );
  AOI21XL U53 ( .A0(n1031), .A1(n49), .B0(n48), .Y(n1021) );
  XOR2XL U54 ( .A(n1041), .B(n1040), .Y(n1276) );
  INVX1 U55 ( .A(n1062), .Y(n13) );
  INVX1 U56 ( .A(n1102), .Y(n12) );
  BUFX3 U57 ( .A(A[5]), .Y(n895) );
  BUFX1 U58 ( .A(A[9]), .Y(n858) );
  OR2X2 U59 ( .A(n554), .B(n555), .Y(n5) );
  XOR2XL U60 ( .A(n1053), .B(n1052), .Y(PRODUCT[36]) );
  NAND2X1 U61 ( .A(n692), .B(n25), .Y(n24) );
  NAND2X1 U62 ( .A(n211), .B(n210), .Y(n824) );
  OR2X2 U63 ( .A(n693), .B(n694), .Y(n25) );
  OAI2BB1XL U64 ( .A0N(n206), .A1N(n205), .B0(n112), .Y(n799) );
  NAND2BXL U65 ( .AN(n329), .B(n42), .Y(n41) );
  XNOR2X1 U66 ( .A(n1102), .B(B[17]), .Y(n324) );
  XNOR2X1 U67 ( .A(n866), .B(B[22]), .Y(n329) );
  OAI22XL U68 ( .A0(n957), .A1(n958), .B0(n956), .B1(n91), .Y(n972) );
  AOI21XL U69 ( .A0(n34), .A1(n226), .B0(n33), .Y(n32) );
  XOR2X2 U70 ( .A(n56), .B(n55), .Y(PRODUCT[18]) );
  INVX1 U71 ( .A(n895), .Y(n9) );
  NAND2X1 U72 ( .A(n593), .B(n1234), .Y(n629) );
  NAND2X1 U73 ( .A(n1190), .B(n1202), .Y(n1132) );
  OR2X2 U74 ( .A(n1246), .B(n53), .Y(n54) );
  INVX1 U75 ( .A(n517), .Y(n11) );
  NAND2X1 U76 ( .A(n235), .B(n1210), .Y(n236) );
  INVXL U77 ( .A(n1247), .Y(n53) );
  INVX1 U78 ( .A(n905), .Y(n8) );
  BUFX3 U79 ( .A(A[11]), .Y(n1062) );
  INVX1 U80 ( .A(n1201), .Y(n1190) );
  BUFX3 U81 ( .A(A[13]), .Y(n1102) );
  XNOR2X1 U82 ( .A(A[12]), .B(A[11]), .Y(n128) );
  INVX1 U83 ( .A(n1239), .Y(n742) );
  INVX1 U84 ( .A(n1227), .Y(n522) );
  INVX1 U85 ( .A(n1235), .Y(n665) );
  XNOR2X1 U86 ( .A(n1036), .B(n1035), .Y(n1275) );
  INVX1 U87 ( .A(n1031), .Y(n1041) );
  NAND2X1 U88 ( .A(n24), .B(n23), .Y(n668) );
  INVX1 U89 ( .A(n825), .Y(n823) );
  INVX1 U90 ( .A(n211), .Y(n22) );
  XNOR2X1 U91 ( .A(n1167), .B(n1166), .Y(n1278) );
  NOR2X1 U92 ( .A(n822), .B(n821), .Y(mult_x_1_n312) );
  INVX1 U93 ( .A(n985), .Y(n1028) );
  OR2X2 U94 ( .A(n511), .B(n510), .Y(n20) );
  NAND2X1 U95 ( .A(n851), .B(n850), .Y(n1044) );
  ADDFHX2 U96 ( .A(n807), .B(n806), .CI(n805), .CO(n817), .S(n211) );
  NAND2X1 U97 ( .A(n939), .B(n938), .Y(n1033) );
  NAND2X1 U98 ( .A(n934), .B(n933), .Y(n1160) );
  ADDFHX1 U99 ( .A(n708), .B(n707), .CI(n706), .CO(n692), .S(n746) );
  NAND2X1 U100 ( .A(n932), .B(n931), .Y(n1164) );
  XNOR2X1 U101 ( .A(n1102), .B(n1147), .Y(n1138) );
  XNOR2X1 U102 ( .A(n1062), .B(n1147), .Y(n1108) );
  XNOR2X1 U103 ( .A(n858), .B(n1147), .Y(n1058) );
  BUFX3 U104 ( .A(B[26]), .Y(n1147) );
  XOR2X1 U105 ( .A(n223), .B(n222), .Y(PRODUCT[37]) );
  NAND2X1 U106 ( .A(n67), .B(n11), .Y(n66) );
  AOI21X1 U107 ( .A0(n380), .A1(n418), .B0(n381), .Y(n382) );
  INVX1 U108 ( .A(n380), .Y(n416) );
  NOR2BX2 U109 ( .AN(n63), .B(n104), .Y(n18) );
  INVX1 U110 ( .A(n697), .Y(n700) );
  AND2X2 U111 ( .A(n312), .B(n1216), .Y(n81) );
  INVX1 U112 ( .A(n908), .Y(n114) );
  AOI21X1 U113 ( .A0(n828), .A1(n1248), .B0(n1254), .Y(n816) );
  INVX1 U114 ( .A(n1217), .Y(n348) );
  INVX1 U115 ( .A(n1221), .Y(n418) );
  INVX1 U116 ( .A(n1209), .Y(n235) );
  INVX1 U117 ( .A(n1242), .Y(n62) );
  INVX1 U118 ( .A(n1205), .Y(n1093) );
  INVX1 U119 ( .A(n905), .Y(n10) );
  NAND2XL U120 ( .A(n668), .B(n669), .Y(n101) );
  XOR2X1 U121 ( .A(n103), .B(n667), .Y(n696) );
  XNOR2X1 U122 ( .A(n1030), .B(n1029), .Y(n1274) );
  INVX1 U123 ( .A(n1021), .Y(n1030) );
  NAND2XL U124 ( .A(n513), .B(n512), .Y(mult_x_1_n224) );
  XOR2X1 U125 ( .A(n1163), .B(n1162), .Y(n1277) );
  ADDFHX1 U126 ( .A(n599), .B(n598), .CI(n597), .CO(n590), .S(n626) );
  NAND2X1 U127 ( .A(n22), .B(n21), .Y(n825) );
  NOR2X1 U128 ( .A(n815), .B(n814), .Y(mult_x_1_n299) );
  NOR2X1 U129 ( .A(n818), .B(n817), .Y(mult_x_1_n302) );
  INVXL U130 ( .A(n1022), .Y(n1027) );
  INVXL U131 ( .A(n387), .Y(n116) );
  OAI2BB1X1 U132 ( .A0N(n509), .A1N(n20), .B0(n92), .Y(n486) );
  INVXL U133 ( .A(n388), .Y(n117) );
  NOR2X1 U134 ( .A(n851), .B(n850), .Y(n1045) );
  OAI21XL U135 ( .A0(n39), .A1(n40), .B0(n38), .Y(n772) );
  XNOR3X2 U136 ( .A(n554), .B(n31), .C(n553), .Y(n561) );
  NAND2XL U137 ( .A(n693), .B(n694), .Y(n23) );
  INVX1 U138 ( .A(n210), .Y(n21) );
  NAND2BXL U139 ( .AN(n1158), .B(n1165), .Y(n51) );
  ADDFHX2 U140 ( .A(n658), .B(n657), .CI(n656), .CO(n632), .S(n667) );
  INVXL U141 ( .A(n776), .Y(n39) );
  INVXL U142 ( .A(n1014), .Y(n76) );
  INVX1 U143 ( .A(n1015), .Y(n75) );
  INVXL U144 ( .A(n986), .Y(n100) );
  OAI2BB1XL U145 ( .A0N(n652), .A1N(n29), .B0(n26), .Y(n645) );
  OR2XL U146 ( .A(n1155), .B(n1154), .Y(n1157) );
  ADDFHX2 U147 ( .A(n1010), .B(n1009), .CI(n1008), .CO(n1012), .S(n989) );
  ADDFHX1 U148 ( .A(n995), .B(n994), .CI(n993), .CO(n850), .S(n1015) );
  ADDFHX1 U149 ( .A(n370), .B(n369), .CI(n368), .CO(n362), .S(n425) );
  NAND2X1 U150 ( .A(n937), .B(n936), .Y(n1038) );
  NOR2X1 U151 ( .A(n937), .B(n936), .Y(n1037) );
  NAND2XL U152 ( .A(n27), .B(n651), .Y(n26) );
  OAI2BB1XL U153 ( .A0N(n956), .A1N(n580), .B0(n250), .Y(n267) );
  NAND2XL U154 ( .A(n975), .B(n974), .Y(n78) );
  OR2XL U155 ( .A(n974), .B(n975), .Y(n79) );
  ADDFHX1 U156 ( .A(n688), .B(n687), .CI(n686), .CO(n680), .S(n748) );
  INVXL U157 ( .A(n182), .Y(n110) );
  INVXL U158 ( .A(n249), .Y(n250) );
  ADDFHX1 U159 ( .A(n972), .B(n971), .CI(n970), .CO(n1000), .S(n981) );
  OAI22XL U160 ( .A0(n77), .A1(n1042), .B0(n947), .B1(n881), .Y(n877) );
  OAI22XL U161 ( .A0(n1114), .A1(n720), .B0(n1141), .B1(n679), .Y(n731) );
  NAND2XL U162 ( .A(n47), .B(n45), .Y(n44) );
  OR2X2 U163 ( .A(n912), .B(n911), .Y(n910) );
  XNOR2X1 U164 ( .A(n1133), .B(n1132), .Y(PRODUCT[39]) );
  AND2XL U165 ( .A(n1183), .B(n1182), .Y(n1283) );
  XNOR2X1 U166 ( .A(n1101), .B(n1100), .Y(PRODUCT[38]) );
  OR2XL U167 ( .A(n1181), .B(n1180), .Y(n1183) );
  AOI2BB1X2 U168 ( .A0N(n559), .A1N(n73), .B0(n66), .Y(n65) );
  OAI22XL U169 ( .A0(n1060), .A1(n949), .B0(n1061), .B1(n948), .Y(n953) );
  NAND2X2 U170 ( .A(n19), .B(n18), .Y(n17) );
  AND2XL U171 ( .A(n1188), .B(n1190), .Y(n1194) );
  INVXL U172 ( .A(n628), .Y(n516) );
  INVXL U173 ( .A(n947), .Y(n45) );
  INVXL U174 ( .A(n958), .Y(n42) );
  CLKINVX3 U175 ( .A(n60), .Y(n16) );
  NAND2BX1 U176 ( .AN(n96), .B(n628), .Y(n19) );
  NAND2BX2 U177 ( .AN(n105), .B(n69), .Y(n628) );
  NOR2BXL U178 ( .AN(B[0]), .B(n1081), .Y(n955) );
  XOR2X2 U179 ( .A(n816), .B(n54), .Y(PRODUCT[17]) );
  AND2X2 U180 ( .A(n1091), .B(n1208), .Y(n1052) );
  NAND2X1 U181 ( .A(n129), .B(n130), .Y(n898) );
  NAND2X1 U182 ( .A(n120), .B(n1111), .Y(n1110) );
  NAND2X1 U183 ( .A(n665), .B(n1236), .Y(n666) );
  NAND2X1 U184 ( .A(n384), .B(n1220), .Y(n385) );
  AND2X2 U185 ( .A(n59), .B(n1230), .Y(n560) );
  NAND2X1 U186 ( .A(n127), .B(n128), .Y(n1140) );
  NAND2X1 U187 ( .A(n379), .B(n215), .Y(n347) );
  NAND2X1 U188 ( .A(n594), .B(n1232), .Y(n595) );
  INVXL U189 ( .A(n514), .Y(n558) );
  NAND2X1 U190 ( .A(n522), .B(n1228), .Y(n523) );
  AND2X2 U191 ( .A(n1093), .B(n1206), .Y(n222) );
  NAND2X1 U192 ( .A(n242), .B(n1212), .Y(n243) );
  INVXL U193 ( .A(n1226), .Y(n36) );
  INVX1 U194 ( .A(n1233), .Y(n593) );
  INVXL U195 ( .A(n1229), .Y(n59) );
  INVX1 U196 ( .A(n1211), .Y(n242) );
  INVXL U197 ( .A(n1241), .Y(n72) );
  CLKINVX3 U198 ( .A(n866), .Y(n14) );
  INVX1 U199 ( .A(n1207), .Y(n1091) );
  INVX1 U200 ( .A(n1237), .Y(n662) );
  XNOR2X1 U201 ( .A(A[14]), .B(A[13]), .Y(n125) );
  NOR2X1 U202 ( .A(n1217), .B(n1215), .Y(n224) );
  NAND2X2 U203 ( .A(n514), .B(n212), .Y(n96) );
  OAI21X4 U204 ( .A0(n1198), .A1(n1225), .B0(n1226), .Y(n452) );
  NOR2X4 U205 ( .A(n17), .B(n15), .Y(n1198) );
  NOR3X4 U206 ( .A(n16), .B(n96), .C(n515), .Y(n15) );
  OAI21X1 U207 ( .A0(n1234), .A1(n1231), .B0(n1232), .Y(n517) );
  XOR2X1 U208 ( .A(B[15]), .B(n10), .Y(n197) );
  XOR3X2 U209 ( .A(n694), .B(n693), .C(n692), .Y(n703) );
  NOR2X1 U210 ( .A(n659), .B(n660), .Y(mult_x_1_n259) );
  OR2X2 U211 ( .A(n652), .B(n29), .Y(n27) );
  XOR2X1 U212 ( .A(n652), .B(n28), .Y(n707) );
  XOR2X1 U213 ( .A(n651), .B(n29), .Y(n28) );
  OAI22X1 U214 ( .A0(n608), .A1(n964), .B0(n966), .B1(n643), .Y(n29) );
  NOR2X1 U215 ( .A(n1227), .B(n1229), .Y(n212) );
  NOR2X2 U216 ( .A(n1233), .B(n1231), .Y(n514) );
  NAND2XL U217 ( .A(n557), .B(n556), .Y(mult_x_1_n233) );
  OAI2BB1X2 U218 ( .A0N(n5), .A1N(n553), .B0(n30), .Y(n526) );
  NAND2X1 U219 ( .A(n554), .B(n555), .Y(n30) );
  INVX1 U220 ( .A(n555), .Y(n31) );
  OAI21XL U221 ( .A0(n218), .A1(n1214), .B0(n217), .Y(n33) );
  NAND2X1 U222 ( .A(n34), .B(n224), .Y(n219) );
  NOR2X1 U223 ( .A(n218), .B(n1213), .Y(n34) );
  NAND2BX1 U224 ( .AN(n1223), .B(n36), .Y(n35) );
  OAI22X1 U225 ( .A0(n500), .A1(n960), .B0(n37), .B1(n962), .Y(n552) );
  XNOR2X1 U226 ( .A(B[18]), .B(n895), .Y(n37) );
  OAI21XL U227 ( .A0(n776), .A1(n777), .B0(n775), .Y(n38) );
  XNOR3X2 U228 ( .A(n40), .B(n775), .C(n776), .Y(n794) );
  INVX1 U229 ( .A(n777), .Y(n40) );
  XNOR2X1 U230 ( .A(B[20]), .B(n1062), .Y(n286) );
  OAI21XL U231 ( .A0(n956), .A1(n43), .B0(n41), .Y(n335) );
  XOR2X2 U232 ( .A(B[23]), .B(n14), .Y(n43) );
  OAI21XL U233 ( .A0(n1042), .A1(n881), .B0(n44), .Y(n889) );
  OAI21XL U234 ( .A0(n914), .A1(n947), .B0(n46), .Y(n900) );
  NAND2XL U235 ( .A(n47), .B(A[0]), .Y(n46) );
  XNOR2X1 U236 ( .A(B[5]), .B(n8), .Y(n47) );
  INVXL U237 ( .A(n935), .Y(n1161) );
  OAI21XL U238 ( .A0(n1032), .A1(n1038), .B0(n1033), .Y(n48) );
  NOR2X1 U239 ( .A(n1037), .B(n1032), .Y(n49) );
  NOR2X1 U240 ( .A(n939), .B(n938), .Y(n1032) );
  NAND3X1 U241 ( .A(n52), .B(n50), .C(n1160), .Y(n1031) );
  OR2X2 U242 ( .A(n935), .B(n51), .Y(n50) );
  OR2X2 U243 ( .A(n935), .B(n1164), .Y(n52) );
  AND2X2 U244 ( .A(n795), .B(n1245), .Y(n55) );
  OAI21XL U245 ( .A0(n816), .A1(n1246), .B0(n1247), .Y(n56) );
  INVX1 U246 ( .A(n1255), .Y(n828) );
  NAND2X1 U247 ( .A(n517), .B(n212), .Y(n63) );
  NOR2X1 U248 ( .A(n73), .B(n664), .Y(n58) );
  CLKINVX3 U249 ( .A(n60), .Y(n73) );
  NAND4X4 U250 ( .A(n86), .B(n87), .C(n1245), .D(n85), .Y(n60) );
  AND2X2 U251 ( .A(n59), .B(n514), .Y(n519) );
  AOI21X1 U252 ( .A0(n60), .A1(n72), .B0(n62), .Y(n61) );
  XNOR2X1 U253 ( .A(n774), .B(n60), .Y(PRODUCT[19]) );
  NOR2X1 U254 ( .A(n1237), .B(n1235), .Y(n106) );
  XNOR2X4 U255 ( .A(n65), .B(n560), .Y(PRODUCT[25]) );
  NAND2BX1 U256 ( .AN(n558), .B(n628), .Y(n67) );
  NAND2X1 U257 ( .A(n697), .B(n106), .Y(n515) );
  NOR2X2 U258 ( .A(n1239), .B(n1241), .Y(n697) );
  INVX1 U259 ( .A(n515), .Y(n627) );
  OAI21X1 U260 ( .A0(n73), .A1(n70), .B0(n68), .Y(n596) );
  NAND2X1 U261 ( .A(n698), .B(n106), .Y(n69) );
  NAND2XL U262 ( .A(n627), .B(n593), .Y(n70) );
  OAI21XL U263 ( .A0(n515), .A1(n73), .B0(n516), .Y(n630) );
  OAI21XL U264 ( .A0(n521), .A1(n73), .B0(n520), .Y(n524) );
  AOI21X1 U265 ( .A0(n1019), .A1(n1090), .B0(n74), .Y(n1046) );
  INVX1 U266 ( .A(n1089), .Y(n74) );
  NAND2X1 U267 ( .A(n1014), .B(n1015), .Y(n1089) );
  NAND2X1 U268 ( .A(n76), .B(n75), .Y(n1090) );
  XOR2X1 U269 ( .A(B[12]), .B(n8), .Y(n143) );
  OAI22X1 U270 ( .A0(n964), .A1(n643), .B0(n678), .B1(n966), .Y(n687) );
  XNOR2X1 U271 ( .A(B[17]), .B(n908), .Y(n643) );
  XOR2X1 U272 ( .A(n1020), .B(n1017), .Y(n1272) );
  OAI22X1 U273 ( .A0(n77), .A1(n947), .B0(n1042), .B1(n860), .Y(n863) );
  XOR2X1 U274 ( .A(n856), .B(n8), .Y(n77) );
  OAI2BB1X1 U275 ( .A0N(n79), .A1N(n973), .B0(n78), .Y(n980) );
  XOR2X1 U276 ( .A(n973), .B(n80), .Y(n982) );
  XOR2X1 U277 ( .A(n975), .B(n974), .Y(n80) );
  OR2X2 U278 ( .A(n989), .B(n988), .Y(n1024) );
  ADDFX2 U279 ( .A(n497), .B(n498), .CI(n499), .CO(n511), .S(n554) );
  OAI22X1 U280 ( .A0(n537), .A1(n495), .B0(n964), .B1(n464), .Y(n504) );
  XNOR2XL U281 ( .A(B[23]), .B(n908), .Y(n94) );
  XNOR2XL U282 ( .A(n866), .B(B[17]), .Y(n502) );
  XNOR2XL U283 ( .A(A[10]), .B(A[9]), .Y(n1111) );
  BUFX3 U284 ( .A(n1198), .Y(n95) );
  XNOR2XL U285 ( .A(n1102), .B(B[13]), .Y(n432) );
  XNOR2XL U286 ( .A(n1062), .B(B[15]), .Y(n437) );
  XNOR2XL U287 ( .A(n895), .B(B[21]), .Y(n436) );
  XNOR2XL U288 ( .A(n866), .B(B[19]), .Y(n438) );
  XNOR2XL U289 ( .A(n895), .B(B[16]), .Y(n613) );
  XNOR2X1 U290 ( .A(n866), .B(B[14]), .Y(n615) );
  NAND2BXL U291 ( .AN(B[0]), .B(n1062), .Y(n176) );
  XOR2X1 U292 ( .A(B[25]), .B(n9), .Y(n323) );
  XOR2XL U293 ( .A(B[25]), .B(n97), .Y(n265) );
  XNOR2XL U294 ( .A(n1102), .B(B[20]), .Y(n251) );
  XNOR2XL U295 ( .A(n895), .B(B[5]), .Y(n961) );
  XNOR2XL U296 ( .A(n866), .B(B[3]), .Y(n957) );
  NOR2XL U297 ( .A(n1128), .B(n1203), .Y(n1188) );
  INVX1 U298 ( .A(A[15]), .Y(n98) );
  XNOR2XL U299 ( .A(n1062), .B(B[23]), .Y(n266) );
  XNOR2X1 U300 ( .A(n1102), .B(B[22]), .Y(n1064) );
  XOR2XL U301 ( .A(B[25]), .B(n13), .Y(n1082) );
  XNOR2XL U302 ( .A(n1102), .B(B[23]), .Y(n1079) );
  XNOR2XL U303 ( .A(A[15]), .B(B[20]), .Y(n1057) );
  XNOR2XL U304 ( .A(n1062), .B(B[4]), .Y(n147) );
  XNOR2XL U305 ( .A(n908), .B(B[12]), .Y(n146) );
  XOR2XL U306 ( .A(n856), .B(n97), .Y(n113) );
  XNOR2XL U307 ( .A(n1102), .B(B[3]), .Y(n187) );
  NOR2BXL U308 ( .AN(B[0]), .B(n1141), .Y(n179) );
  OAI22XL U309 ( .A0(n1083), .A1(n836), .B0(n1081), .B1(n144), .Y(n177) );
  OAI22X1 U310 ( .A0(n107), .A1(n947), .B0(n1042), .B1(n143), .Y(n178) );
  XNOR2XL U311 ( .A(n866), .B(B[8]), .Y(n148) );
  NAND2BXL U312 ( .AN(B[0]), .B(n1102), .Y(n134) );
  XNOR2X1 U313 ( .A(n1062), .B(B[22]), .Y(n252) );
  XNOR2XL U314 ( .A(n905), .B(B[4]), .Y(n914) );
  XOR2XL U315 ( .A(B[25]), .B(n98), .Y(n1151) );
  XNOR2XL U316 ( .A(A[15]), .B(B[24]), .Y(n1137) );
  XNOR2XL U317 ( .A(A[15]), .B(B[23]), .Y(n1112) );
  XOR2XL U318 ( .A(B[25]), .B(n12), .Y(n1113) );
  XNOR2XL U319 ( .A(n1102), .B(B[24]), .Y(n1103) );
  NAND2BX1 U320 ( .AN(n181), .B(n110), .Y(n109) );
  ADDFX2 U321 ( .A(n893), .B(n84), .CI(n891), .CO(n933), .S(n932) );
  OAI22XL U322 ( .A0(n966), .A1(n894), .B0(n964), .B1(n886), .Y(n893) );
  OAI22XL U323 ( .A0(n898), .A1(n897), .B0(n960), .B1(n896), .Y(n923) );
  OAI22XL U324 ( .A0(n966), .A1(n916), .B0(n964), .B1(n894), .Y(n924) );
  AOI21XL U325 ( .A0(n1186), .A1(n1185), .B0(n930), .Y(n1158) );
  INVXL U326 ( .A(n1184), .Y(n930) );
  INVXL U327 ( .A(n226), .Y(n279) );
  INVXL U328 ( .A(n1218), .Y(n309) );
  INVXL U329 ( .A(n1195), .Y(n1050) );
  NAND2XL U330 ( .A(n483), .B(n1226), .Y(n484) );
  XNOR2X2 U331 ( .A(n524), .B(n523), .Y(PRODUCT[26]) );
  INVXL U332 ( .A(n1219), .Y(n384) );
  XNOR2X1 U333 ( .A(n630), .B(n629), .Y(PRODUCT[23]) );
  OAI21X1 U334 ( .A0(n95), .A1(n281), .B0(n280), .Y(n284) );
  XNOR2XL U335 ( .A(n1148), .B(B[11]), .Y(n430) );
  XOR2X1 U336 ( .A(B[18]), .B(n97), .Y(n396) );
  INVXL U337 ( .A(A[9]), .Y(n97) );
  XNOR2XL U338 ( .A(n1102), .B(B[14]), .Y(n398) );
  XNOR2X1 U339 ( .A(B[20]), .B(n866), .Y(n404) );
  XNOR2XL U340 ( .A(n1062), .B(B[12]), .Y(n545) );
  XNOR2XL U341 ( .A(n866), .B(B[16]), .Y(n546) );
  XNOR2XL U342 ( .A(n1062), .B(B[9]), .Y(n649) );
  XNOR2X1 U343 ( .A(n895), .B(B[15]), .Y(n648) );
  XNOR2XL U344 ( .A(n866), .B(B[13]), .Y(n650) );
  XNOR2XL U345 ( .A(n858), .B(B[11]), .Y(n642) );
  XNOR2XL U346 ( .A(n1102), .B(n856), .Y(n644) );
  XNOR2XL U347 ( .A(n1062), .B(B[8]), .Y(n684) );
  XNOR2XL U348 ( .A(n866), .B(B[12]), .Y(n685) );
  XNOR2XL U349 ( .A(n1102), .B(B[6]), .Y(n679) );
  XNOR2XL U350 ( .A(n1148), .B(B[14]), .Y(n330) );
  XNOR2XL U351 ( .A(n866), .B(B[21]), .Y(n357) );
  XOR2X1 U352 ( .A(B[25]), .B(n114), .Y(n365) );
  XNOR2XL U353 ( .A(n908), .B(B[24]), .Y(n397) );
  XOR2X1 U354 ( .A(B[22]), .B(n9), .Y(n402) );
  XNOR2XL U355 ( .A(n1102), .B(B[16]), .Y(n356) );
  XNOR2XL U356 ( .A(n866), .B(B[11]), .Y(n729) );
  XNOR2XL U357 ( .A(n1102), .B(B[5]), .Y(n720) );
  XNOR2XL U358 ( .A(n1062), .B(B[5]), .Y(n189) );
  XNOR2XL U359 ( .A(n895), .B(B[12]), .Y(n726) );
  XNOR2XL U360 ( .A(n866), .B(B[9]), .Y(n190) );
  XNOR2XL U361 ( .A(n866), .B(B[10]), .Y(n730) );
  XNOR2XL U362 ( .A(n858), .B(B[8]), .Y(n717) );
  XNOR2XL U363 ( .A(n1102), .B(B[4]), .Y(n721) );
  XNOR2XL U364 ( .A(n895), .B(B[11]), .Y(n188) );
  XNOR2X1 U365 ( .A(n1148), .B(B[15]), .Y(n314) );
  XOR2XL U366 ( .A(B[18]), .B(n12), .Y(n289) );
  XNOR2XL U367 ( .A(n1102), .B(B[19]), .Y(n255) );
  NAND2BXL U368 ( .AN(B[0]), .B(n895), .Y(n887) );
  XNOR2XL U369 ( .A(n895), .B(B[4]), .Y(n854) );
  NAND2XL U370 ( .A(n1099), .B(n1204), .Y(n1100) );
  INVXL U371 ( .A(n1203), .Y(n1099) );
  CMPR32X1 U372 ( .A(n407), .B(n406), .C(n405), .CO(n399), .S(n457) );
  OAI2BB1XL U373 ( .A0N(n1042), .A1N(n947), .B0(n361), .Y(n405) );
  OAI22XL U374 ( .A0(n1060), .A1(n396), .B0(n1061), .B1(n359), .Y(n407) );
  OAI22XL U375 ( .A0(n1152), .A1(n393), .B0(n1150), .B1(n360), .Y(n406) );
  XNOR2XL U376 ( .A(n1062), .B(B[24]), .Y(n1063) );
  OAI22XL U377 ( .A0(n1114), .A1(n465), .B0(n1141), .B1(n432), .Y(n472) );
  OAI22XL U378 ( .A0(n1060), .A1(n463), .B0(n1061), .B1(n431), .Y(n474) );
  OAI22XL U379 ( .A0(n958), .A1(n471), .B0(n956), .B1(n438), .Y(n475) );
  OAI22XL U380 ( .A0(n962), .A1(n469), .B0(n960), .B1(n436), .Y(n477) );
  ADDFX2 U381 ( .A(n505), .B(n504), .CI(n503), .CO(n497), .S(n565) );
  OAI22XL U382 ( .A0(n1114), .A1(n496), .B0(n1141), .B1(n465), .Y(n503) );
  CMPR32X1 U383 ( .A(n508), .B(n507), .C(n506), .CO(n530), .S(n564) );
  OAI22XL U384 ( .A0(n1083), .A1(n501), .B0(n1081), .B1(n470), .Y(n507) );
  OAI22XL U385 ( .A0(n1114), .A1(n538), .B0(n1141), .B1(n496), .Y(n547) );
  OAI22XL U386 ( .A0(n1114), .A1(n573), .B0(n1141), .B1(n538), .Y(n581) );
  CMPR32X1 U387 ( .A(n621), .B(n620), .C(n619), .CO(n636), .S(n670) );
  OAI22XL U388 ( .A0(n580), .A1(n615), .B0(n956), .B1(n579), .Y(n619) );
  OAI22XL U389 ( .A0(n1083), .A1(n614), .B0(n1081), .B1(n578), .Y(n620) );
  ADDFX2 U390 ( .A(n682), .B(n681), .CI(n680), .CO(n694), .S(n738) );
  OAI22XL U391 ( .A0(n1083), .A1(n837), .B0(n1081), .B1(n836), .Y(n968) );
  OAI22X1 U392 ( .A0(n835), .A1(n956), .B0(n958), .B1(n91), .Y(n969) );
  OAI22XL U393 ( .A0(n966), .A1(n963), .B0(n964), .B1(n838), .Y(n967) );
  OAI22XL U394 ( .A0(n1060), .A1(n840), .B0(n1061), .B1(n175), .Y(n998) );
  XNOR2XL U395 ( .A(n1062), .B(B[21]), .Y(n256) );
  OAI22XL U396 ( .A0(n1114), .A1(n251), .B0(n1141), .B1(n263), .Y(n272) );
  OAI22XL U397 ( .A0(n1060), .A1(n253), .B0(n1061), .B1(n265), .Y(n270) );
  OAI2BB1XL U398 ( .A0N(n960), .A1N(n962), .B0(n247), .Y(n294) );
  OAI22XL U399 ( .A0(n1152), .A1(n288), .B0(n1150), .B1(n245), .Y(n296) );
  INVXL U400 ( .A(n246), .Y(n247) );
  INVXL U401 ( .A(n1192), .Y(n1193) );
  AOI21XL U402 ( .A0(n1191), .A1(n1190), .B0(n1189), .Y(n1192) );
  INVXL U403 ( .A(n1202), .Y(n1189) );
  NAND2XL U404 ( .A(n213), .B(n1188), .Y(n1131) );
  OAI2BB1XL U405 ( .A0N(n1111), .A1N(n1110), .B0(n1109), .Y(n1115) );
  OAI22XL U406 ( .A0(n1152), .A1(n1107), .B0(n1150), .B1(n1112), .Y(n1116) );
  INVXL U407 ( .A(n1108), .Y(n1109) );
  OAI22XL U408 ( .A0(n1152), .A1(n1080), .B0(n1150), .B1(n1107), .Y(n1105) );
  OAI22XL U409 ( .A0(n1114), .A1(n1079), .B0(n1141), .B1(n1103), .Y(n1106) );
  INVXL U410 ( .A(n1117), .Y(n1104) );
  OAI22XL U411 ( .A0(n1114), .A1(n263), .B0(n1141), .B1(n1064), .Y(n1067) );
  OAI22XL U412 ( .A0(n1152), .A1(n264), .B0(n1150), .B1(n1057), .Y(n1066) );
  INVXL U413 ( .A(n1077), .Y(n1065) );
  ADDFX2 U414 ( .A(n468), .B(n83), .CI(n466), .CO(n480), .S(n510) );
  INVX1 U415 ( .A(n82), .Y(n83) );
  INVXL U416 ( .A(n467), .Y(n82) );
  CMPR32X1 U417 ( .A(n165), .B(n164), .C(n163), .CO(n206), .S(n166) );
  OAI22XL U418 ( .A0(n1114), .A1(n153), .B0(n1141), .B1(n187), .Y(n201) );
  OAI22XL U419 ( .A0(n1152), .A1(n126), .B0(n1150), .B1(n198), .Y(n202) );
  OAI22XL U420 ( .A0(n1083), .A1(n144), .B0(n1081), .B1(n137), .Y(n169) );
  OAI22XL U421 ( .A0(n1114), .A1(n136), .B0(n1141), .B1(n154), .Y(n170) );
  CMPR32X1 U422 ( .A(n140), .B(n139), .C(n138), .CO(n204), .S(n181) );
  NOR2BXL U423 ( .AN(B[0]), .B(n960), .Y(n927) );
  OAI22XL U424 ( .A0(n966), .A1(n917), .B0(n964), .B1(n916), .Y(n925) );
  OAI22XL U425 ( .A0(n947), .A1(n915), .B0(n914), .B1(n1042), .Y(n926) );
  CMPR32X1 U426 ( .A(n875), .B(n874), .C(n873), .CO(n938), .S(n937) );
  OAI22XL U427 ( .A0(n1152), .A1(n1151), .B0(n1150), .B1(n1149), .Y(n1153) );
  NOR2BX1 U428 ( .AN(n987), .B(n100), .Y(n1022) );
  OAI2BB1XL U429 ( .A0N(n1141), .A1N(n1140), .B0(n1139), .Y(n1144) );
  OAI22XL U430 ( .A0(n1152), .A1(n1137), .B0(n1150), .B1(n1151), .Y(n1145) );
  INVXL U431 ( .A(n1138), .Y(n1139) );
  OAI22XL U432 ( .A0(n947), .A1(B[0]), .B0(n901), .B1(n1042), .Y(n1181) );
  NAND2XL U433 ( .A(n902), .B(n947), .Y(n1180) );
  NAND2BXL U434 ( .AN(B[0]), .B(n905), .Y(n902) );
  NAND2XL U435 ( .A(n1181), .B(n1180), .Y(n1182) );
  NOR2XL U436 ( .A(n921), .B(n920), .Y(n1168) );
  NAND2XL U437 ( .A(n921), .B(n920), .Y(n1169) );
  AOI21XL U438 ( .A0(n1174), .A1(n910), .B0(n913), .Y(n1171) );
  INVXL U439 ( .A(n1173), .Y(n913) );
  NAND2XL U440 ( .A(n929), .B(n928), .Y(n1184) );
  INVXL U441 ( .A(n1158), .Y(n1166) );
  INVXL U442 ( .A(n213), .Y(n1051) );
  INVXL U443 ( .A(n1208), .Y(n1094) );
  INVXL U444 ( .A(n1128), .Y(n1096) );
  INVXL U445 ( .A(n1222), .Y(n381) );
  NAND2XL U446 ( .A(n379), .B(n418), .Y(n383) );
  AOI21XL U447 ( .A0(n698), .A1(n662), .B0(n661), .Y(n663) );
  INVXL U448 ( .A(n1238), .Y(n661) );
  INVXL U449 ( .A(n1234), .Y(n592) );
  INVXL U450 ( .A(n1214), .Y(n228) );
  INVX1 U451 ( .A(n1250), .Y(n826) );
  XNOR2XL U452 ( .A(n1148), .B(B[6]), .Y(n606) );
  XNOR2XL U453 ( .A(n1148), .B(B[5]), .Y(n640) );
  XNOR2XL U454 ( .A(n1148), .B(B[4]), .Y(n676) );
  XNOR2XL U455 ( .A(n1148), .B(B[3]), .Y(n714) );
  XNOR2XL U456 ( .A(n905), .B(B[16]), .Y(n712) );
  NAND2BXL U457 ( .AN(B[0]), .B(n858), .Y(n859) );
  INVXL U458 ( .A(n1212), .Y(n227) );
  AOI21XL U459 ( .A0(n1094), .A1(n1093), .B0(n1092), .Y(n1129) );
  INVXL U460 ( .A(n1206), .Y(n1092) );
  NOR2XL U461 ( .A(n1225), .B(n1223), .Y(n379) );
  AOI21XL U462 ( .A0(n1195), .A1(n1096), .B0(n1095), .Y(n1097) );
  INVXL U463 ( .A(n1129), .Y(n1095) );
  NAND2XL U464 ( .A(n213), .B(n1096), .Y(n1098) );
  NAND2XL U465 ( .A(n1091), .B(n1093), .Y(n1128) );
  NAND2XL U466 ( .A(n72), .B(n1242), .Y(n774) );
  XNOR2X2 U467 ( .A(n596), .B(n595), .Y(PRODUCT[24]) );
  INVXL U468 ( .A(n1231), .Y(n594) );
  INVXL U469 ( .A(n1215), .Y(n312) );
  INVXL U470 ( .A(n392), .Y(n361) );
  XNOR2XL U471 ( .A(n1148), .B(B[12]), .Y(n393) );
  XNOR2XL U472 ( .A(n1102), .B(B[12]), .Y(n465) );
  XNOR2XL U473 ( .A(n1062), .B(B[14]), .Y(n470) );
  XNOR2XL U474 ( .A(n1102), .B(B[11]), .Y(n496) );
  XNOR2XL U475 ( .A(n905), .B(B[21]), .Y(n569) );
  XNOR2XL U476 ( .A(n1148), .B(n856), .Y(n570) );
  XNOR2XL U477 ( .A(n1148), .B(B[8]), .Y(n532) );
  XNOR2X1 U478 ( .A(n858), .B(B[14]), .Y(n535) );
  XNOR2XL U479 ( .A(n1102), .B(B[10]), .Y(n538) );
  XNOR2XL U480 ( .A(n1062), .B(B[11]), .Y(n578) );
  XNOR2X1 U481 ( .A(n866), .B(B[15]), .Y(n579) );
  XNOR2XL U482 ( .A(n1102), .B(B[9]), .Y(n573) );
  XNOR2XL U483 ( .A(n858), .B(B[12]), .Y(n607) );
  XNOR2XL U484 ( .A(n1102), .B(B[8]), .Y(n609) );
  XNOR2XL U485 ( .A(n895), .B(B[6]), .Y(n959) );
  XOR2XL U486 ( .A(B[4]), .B(n14), .Y(n91) );
  XNOR2XL U487 ( .A(n908), .B(B[8]), .Y(n963) );
  XNOR2XL U488 ( .A(n866), .B(B[5]), .Y(n835) );
  XNOR2XL U489 ( .A(B[11]), .B(n905), .Y(n107) );
  XNOR2XL U490 ( .A(n895), .B(B[8]), .Y(n162) );
  XNOR2XL U491 ( .A(n858), .B(B[4]), .Y(n175) );
  XNOR2XL U492 ( .A(n858), .B(B[3]), .Y(n840) );
  XNOR2XL U493 ( .A(n895), .B(B[24]), .Y(n328) );
  NAND2BXL U494 ( .AN(B[0]), .B(n1148), .Y(n150) );
  XNOR2XL U495 ( .A(n908), .B(n856), .Y(n965) );
  XNOR2XL U496 ( .A(n895), .B(B[3]), .Y(n865) );
  XNOR2XL U497 ( .A(n908), .B(B[5]), .Y(n869) );
  AOI21XL U498 ( .A0(n235), .A1(n227), .B0(n216), .Y(n217) );
  INVXL U499 ( .A(n1210), .Y(n216) );
  AOI21XL U500 ( .A0(n1195), .A1(n1188), .B0(n1191), .Y(n1130) );
  XNOR2X1 U501 ( .A(A[15]), .B(B[22]), .Y(n1107) );
  XNOR2XL U502 ( .A(A[15]), .B(B[19]), .Y(n264) );
  XNOR2XL U503 ( .A(n1102), .B(B[21]), .Y(n263) );
  OAI22X1 U504 ( .A0(n713), .A1(n461), .B0(n429), .B1(n1042), .Y(n460) );
  OAI22XL U505 ( .A0(n1114), .A1(n432), .B0(n1141), .B1(n398), .Y(n439) );
  OAI22X1 U506 ( .A0(n397), .A1(n964), .B0(n966), .B1(n94), .Y(n440) );
  OAI22X1 U507 ( .A0(n1060), .A1(n431), .B0(n1061), .B1(n396), .Y(n441) );
  OAI22XL U508 ( .A0(n962), .A1(n436), .B0(n960), .B1(n402), .Y(n444) );
  CMPR32X1 U509 ( .A(n552), .B(n551), .C(n550), .CO(n566), .S(n600) );
  OAI22XL U510 ( .A0(n1083), .A1(n545), .B0(n1081), .B1(n501), .Y(n551) );
  ADDFX2 U511 ( .A(n612), .B(n611), .CI(n610), .CO(n624), .S(n657) );
  OAI22XL U512 ( .A0(n1114), .A1(n644), .B0(n1141), .B1(n609), .Y(n651) );
  OAI22XL U513 ( .A0(n1060), .A1(n642), .B0(n1061), .B1(n607), .Y(n652) );
  OAI22XL U514 ( .A0(n958), .A1(n650), .B0(n956), .B1(n615), .Y(n653) );
  OAI22XL U515 ( .A0(n958), .A1(n685), .B0(n956), .B1(n650), .Y(n689) );
  OAI22XL U516 ( .A0(n1114), .A1(n679), .B0(n1141), .B1(n644), .Y(n686) );
  OAI22XL U517 ( .A0(n958), .A1(n729), .B0(n956), .B1(n685), .Y(n734) );
  XNOR2XL U518 ( .A(n908), .B(B[11]), .Y(n159) );
  XNOR2XL U519 ( .A(n858), .B(B[6]), .Y(n123) );
  XNOR2XL U520 ( .A(n866), .B(B[6]), .Y(n145) );
  XNOR2XL U521 ( .A(n1062), .B(B[3]), .Y(n137) );
  NOR2BXL U522 ( .AN(B[0]), .B(n1150), .Y(n157) );
  OAI22XL U523 ( .A0(n1114), .A1(n154), .B0(n1141), .B1(n153), .Y(n155) );
  XNOR2XL U524 ( .A(n895), .B(B[9]), .Y(n161) );
  XNOR2XL U525 ( .A(n895), .B(B[10]), .Y(n149) );
  OAI2BB1XL U526 ( .A0N(n964), .A1N(n537), .B0(n316), .Y(n332) );
  CMPR32X1 U527 ( .A(n373), .B(n372), .C(n371), .CO(n391), .S(n424) );
  OAI22XL U528 ( .A0(n1060), .A1(n359), .B0(n1061), .B1(n331), .Y(n371) );
  OAI22XL U529 ( .A0(n1152), .A1(n360), .B0(n1150), .B1(n330), .Y(n372) );
  OAI22XL U530 ( .A0(n958), .A1(n357), .B0(n956), .B1(n329), .Y(n373) );
  OAI22XL U531 ( .A0(n1110), .A1(n403), .B0(n1081), .B1(n366), .Y(n409) );
  OAI22XL U532 ( .A0(n1140), .A1(n358), .B0(n1141), .B1(n356), .Y(n401) );
  OAI22XL U533 ( .A0(n958), .A1(n730), .B0(n956), .B1(n729), .Y(n766) );
  OAI22XL U534 ( .A0(n1114), .A1(n721), .B0(n1141), .B1(n720), .Y(n763) );
  OAI22XL U535 ( .A0(n958), .A1(n148), .B0(n956), .B1(n190), .Y(n183) );
  OAI22XL U536 ( .A0(n958), .A1(n190), .B0(n956), .B1(n730), .Y(n760) );
  OAI22XL U537 ( .A0(n1114), .A1(n187), .B0(n1141), .B1(n721), .Y(n754) );
  OAI22XL U538 ( .A0(n1060), .A1(n113), .B0(n717), .B1(n1061), .Y(n756) );
  OAI22XL U539 ( .A0(n1060), .A1(n325), .B0(n1061), .B1(n290), .Y(n317) );
  OAI22XL U540 ( .A0(n1140), .A1(n289), .B0(n1141), .B1(n255), .Y(n292) );
  OAI22XL U541 ( .A0(n958), .A1(n287), .B0(n956), .B1(n254), .Y(n293) );
  OAI22XL U542 ( .A0(n1140), .A1(n255), .B0(n1141), .B1(n251), .Y(n259) );
  XNOR2XL U543 ( .A(n905), .B(B[3]), .Y(n915) );
  XNOR2XL U544 ( .A(n908), .B(B[4]), .Y(n886) );
  OAI22XL U545 ( .A0(n962), .A1(n9), .B0(n960), .B1(n887), .Y(n899) );
  XNOR2XL U546 ( .A(n908), .B(B[3]), .Y(n894) );
  NOR2BXL U547 ( .AN(B[0]), .B(n956), .Y(n890) );
  OAI22XL U548 ( .A0(n962), .A1(n896), .B0(n960), .B1(n882), .Y(n888) );
  OAI22XL U549 ( .A0(n958), .A1(n14), .B0(n956), .B1(n855), .Y(n876) );
  NAND2BXL U550 ( .AN(B[0]), .B(n866), .Y(n855) );
  CMPR32X1 U551 ( .A(n952), .B(n951), .C(n950), .CO(n976), .S(n984) );
  OAI22XL U552 ( .A0(n1060), .A1(n853), .B0(n1061), .B1(n949), .Y(n951) );
  OAI22XL U553 ( .A0(n962), .A1(n854), .B0(n960), .B1(n961), .Y(n950) );
  NOR2BXL U554 ( .AN(B[0]), .B(n1061), .Y(n864) );
  OAI22XL U555 ( .A0(n958), .A1(n867), .B0(n956), .B1(n861), .Y(n862) );
  INVX1 U556 ( .A(A[0]), .Y(n133) );
  OAI22XL U557 ( .A0(n1083), .A1(n266), .B0(n1111), .B1(n1063), .Y(n1070) );
  OAI22XL U558 ( .A0(n1114), .A1(n1064), .B0(n1141), .B1(n1079), .Y(n1085) );
  OAI22XL U559 ( .A0(n1083), .A1(n1063), .B0(n1111), .B1(n1082), .Y(n1086) );
  OAI2BB1XL U560 ( .A0N(n1061), .A1N(n1060), .B0(n1059), .Y(n1076) );
  OAI22XL U561 ( .A0(n1152), .A1(n1057), .B0(n1150), .B1(n1080), .Y(n1078) );
  INVXL U562 ( .A(n1058), .Y(n1059) );
  NAND2X1 U563 ( .A(n541), .B(n540), .Y(n589) );
  NAND2XL U564 ( .A(n575), .B(n576), .Y(n540) );
  NAND2XL U565 ( .A(n539), .B(n574), .Y(n541) );
  ADDFX2 U566 ( .A(n749), .B(n748), .CI(n747), .CO(n737), .S(n777) );
  ADDFX2 U567 ( .A(n792), .B(n791), .CI(n790), .CO(n776), .S(n808) );
  NAND2X1 U568 ( .A(n89), .B(n88), .Y(n1006) );
  NAND2X1 U569 ( .A(n1001), .B(n1000), .Y(n88) );
  OAI21XL U570 ( .A0(n1001), .A1(n1000), .B0(n999), .Y(n89) );
  ADDFX2 U571 ( .A(n413), .B(n412), .CI(n411), .CO(n387), .S(n421) );
  CMPR32X1 U572 ( .A(n193), .B(n192), .C(n191), .CO(n806), .S(n207) );
  ADDFX2 U573 ( .A(n801), .B(n800), .CI(n799), .CO(n812), .S(n805) );
  OAI21XL U574 ( .A0(n205), .A1(n206), .B0(n204), .Y(n112) );
  OAI22XL U575 ( .A0(n1083), .A1(n256), .B0(n1081), .B1(n252), .Y(n262) );
  OAI22XL U576 ( .A0(n1152), .A1(n245), .B0(n1150), .B1(n248), .Y(n261) );
  ADDFX2 U577 ( .A(n299), .B(n298), .CI(n297), .CO(n343), .S(n338) );
  OAI22XL U578 ( .A0(n1060), .A1(n290), .B0(n1061), .B1(n285), .Y(n299) );
  ADDFX2 U579 ( .A(n340), .B(n339), .CI(n338), .CO(n342), .S(n350) );
  ADDFX2 U580 ( .A(n302), .B(n301), .CI(n300), .CO(n303), .S(n341) );
  OAI22XL U581 ( .A0(n947), .A1(n901), .B0(n906), .B1(n1042), .Y(n904) );
  NOR2BXL U582 ( .AN(B[0]), .B(n964), .Y(n903) );
  OAI22XL U583 ( .A0(n966), .A1(n114), .B0(n964), .B1(n909), .Y(n911) );
  NAND2BXL U584 ( .AN(B[0]), .B(n908), .Y(n909) );
  NAND2XL U585 ( .A(n213), .B(n1194), .Y(n1197) );
  AOI21XL U586 ( .A0(n1195), .A1(n1194), .B0(n1193), .Y(n1196) );
  NOR2XL U587 ( .A(n1013), .B(n1012), .Y(n1011) );
  ADDFX2 U588 ( .A(n487), .B(n486), .CI(n485), .CO(n481), .S(n513) );
  NAND2X1 U589 ( .A(n511), .B(n510), .Y(n92) );
  INVXL U590 ( .A(n1011), .Y(n1018) );
  NAND2X1 U591 ( .A(n1013), .B(n1012), .Y(n1016) );
  OAI22XL U592 ( .A0(n1152), .A1(n1112), .B0(n1150), .B1(n1137), .Y(n1136) );
  INVXL U593 ( .A(n1146), .Y(n1135) );
  OAI22XL U594 ( .A0(n1114), .A1(n1103), .B0(n1141), .B1(n1113), .Y(n1125) );
  ADDFX2 U595 ( .A(n1056), .B(n1055), .CI(n1054), .CO(n1072), .S(n276) );
  ADDFX2 U596 ( .A(n1075), .B(n1074), .CI(n1073), .CO(n1088), .S(n1071) );
  XOR3X2 U597 ( .A(n388), .B(n387), .C(n386), .Y(n415) );
  XOR2X1 U598 ( .A(n509), .B(n93), .Y(n525) );
  XOR2X1 U599 ( .A(n510), .B(n511), .Y(n93) );
  NAND2X1 U600 ( .A(n102), .B(n101), .Y(n659) );
  OAI21XL U601 ( .A0(n668), .A1(n669), .B0(n667), .Y(n102) );
  XOR2X1 U602 ( .A(n668), .B(n669), .Y(n103) );
  XOR3X2 U603 ( .A(n206), .B(n204), .C(n205), .Y(n209) );
  OAI2BB1X2 U604 ( .A0N(n109), .A1N(n180), .B0(n108), .Y(n208) );
  NAND2X1 U605 ( .A(n181), .B(n182), .Y(n108) );
  OAI21XL U606 ( .A0(n117), .A1(n116), .B0(n115), .Y(n377) );
  OAI21XL U607 ( .A0(n387), .A1(n388), .B0(n386), .Y(n115) );
  NOR2XL U608 ( .A(n904), .B(n903), .Y(n1176) );
  NAND2XL U609 ( .A(n904), .B(n903), .Y(n1177) );
  NAND2XL U610 ( .A(n912), .B(n911), .Y(n1173) );
  OAI21XL U611 ( .A0(n823), .A1(mult_x_1_n313), .B0(n824), .Y(mult_x_1_n306)
         );
  NAND2XL U612 ( .A(n1157), .B(n1156), .Y(mult_x_1_n54) );
  NAND2XL U613 ( .A(n1155), .B(n1154), .Y(n1156) );
  INVXL U614 ( .A(n1153), .Y(n1154) );
  NOR2BXL U615 ( .AN(B[0]), .B(n1042), .Y(n1284) );
  NOR2XL U616 ( .A(n414), .B(n415), .Y(mult_x_1_n202) );
  NOR2XL U617 ( .A(n1143), .B(n1142), .Y(mult_x_1_n105) );
  NAND2XL U618 ( .A(n1143), .B(n1142), .Y(mult_x_1_n106) );
  NOR2XL U619 ( .A(n1119), .B(n1118), .Y(mult_x_1_n114) );
  NAND2XL U620 ( .A(n1119), .B(n1118), .Y(mult_x_1_n115) );
  NOR2XL U621 ( .A(n1127), .B(n1126), .Y(mult_x_1_n125) );
  NAND2XL U622 ( .A(n1127), .B(n1126), .Y(mult_x_1_n126) );
  NOR2XL U623 ( .A(n1088), .B(n1087), .Y(mult_x_1_n134) );
  NAND2XL U624 ( .A(n1088), .B(n1087), .Y(mult_x_1_n135) );
  NOR2XL U625 ( .A(n1072), .B(n1071), .Y(mult_x_1_n149) );
  NAND2XL U626 ( .A(n1072), .B(n1071), .Y(mult_x_1_n150) );
  NAND2XL U627 ( .A(n415), .B(n414), .Y(mult_x_1_n203) );
  XOR2XL U628 ( .A(n1179), .B(n1182), .Y(n1282) );
  NAND2XL U629 ( .A(n1178), .B(n1177), .Y(n1179) );
  INVXL U630 ( .A(n1176), .Y(n1178) );
  XNOR2XL U631 ( .A(n1175), .B(n1174), .Y(n1281) );
  NAND2XL U632 ( .A(n910), .B(n1173), .Y(n1175) );
  XOR2XL U633 ( .A(n1172), .B(n1171), .Y(n1280) );
  NAND2XL U634 ( .A(n1170), .B(n1169), .Y(n1172) );
  INVXL U635 ( .A(n1168), .Y(n1170) );
  NAND2XL U636 ( .A(n1185), .B(n1184), .Y(n1187) );
  NAND2XL U637 ( .A(n1165), .B(n1164), .Y(n1167) );
  AOI21XL U638 ( .A0(n1166), .A1(n1165), .B0(n1159), .Y(n1163) );
  NAND2XL U639 ( .A(n1161), .B(n1160), .Y(n1162) );
  NAND2XL U640 ( .A(n1039), .B(n1038), .Y(n1040) );
  NAND2XL U641 ( .A(n1034), .B(n1033), .Y(n1035) );
  INVX1 U642 ( .A(n225), .Y(n346) );
  NOR2X1 U643 ( .A(n219), .B(n347), .Y(n213) );
  XNOR2X1 U644 ( .A(n905), .B(B[25]), .Y(n429) );
  XNOR2X1 U645 ( .A(n905), .B(B[24]), .Y(n461) );
  OAI22X1 U646 ( .A0(n713), .A1(n197), .B0(n712), .B1(n1042), .Y(n753) );
  OAI22X1 U647 ( .A0(n1152), .A1(n532), .B0(n1150), .B1(n493), .Y(n533) );
  OAI22X1 U648 ( .A0(n641), .A1(n570), .B0(n1150), .B1(n532), .Y(n567) );
  OAI22X1 U649 ( .A0(n1060), .A1(n677), .B0(n1061), .B1(n642), .Y(n688) );
  OAI22X1 U650 ( .A0(n966), .A1(n857), .B0(n964), .B1(n965), .Y(n975) );
  OAI22X1 U651 ( .A0(n962), .A1(n323), .B0(n960), .B1(n246), .Y(n295) );
  OAI22X1 U652 ( .A0(n580), .A1(n254), .B0(n956), .B1(n249), .Y(n268) );
  XOR2X1 U653 ( .A(B[25]), .B(n14), .Y(n254) );
  BUFX1 U654 ( .A(n892), .Y(n84) );
  OAI22X1 U655 ( .A0(n1114), .A1(n398), .B0(n1141), .B1(n358), .Y(n394) );
  OAI22X1 U656 ( .A0(n1152), .A1(n430), .B0(n1150), .B1(n393), .Y(n427) );
  OAI22X1 U657 ( .A0(n1152), .A1(n606), .B0(n1150), .B1(n570), .Y(n603) );
  OAI22X1 U658 ( .A0(n641), .A1(n493), .B0(n1150), .B1(n462), .Y(n491) );
  CMPR22X1 U659 ( .A(n751), .B(n750), .CO(n758), .S(n786) );
  NAND2X1 U660 ( .A(n662), .B(n1238), .Y(n701) );
  NAND2X1 U661 ( .A(n742), .B(n1240), .Y(n743) );
  OAI22X2 U662 ( .A0(n1083), .A1(n578), .B0(n1081), .B1(n545), .Y(n585) );
  OAI22X1 U663 ( .A0(n123), .A1(n841), .B0(n1061), .B1(n113), .Y(n203) );
  OAI22XL U664 ( .A0(n841), .A1(n158), .B0(n1061), .B1(n123), .Y(n165) );
  XNOR2X1 U665 ( .A(n866), .B(B[24]), .Y(n287) );
  XNOR2X1 U666 ( .A(A[9]), .B(B[17]), .Y(n431) );
  XNOR2X1 U667 ( .A(n905), .B(B[17]), .Y(n711) );
  XNOR2X1 U668 ( .A(n895), .B(B[17]), .Y(n577) );
  NAND2X1 U669 ( .A(n1254), .B(n1243), .Y(n85) );
  NAND2BX2 U670 ( .AN(n1244), .B(n53), .Y(n86) );
  NAND3BX2 U671 ( .AN(n1255), .B(n1243), .C(n1248), .Y(n87) );
  XNOR2X1 U672 ( .A(B[20]), .B(n908), .Y(n536) );
  XOR2X1 U673 ( .A(n90), .B(n999), .Y(n1008) );
  XOR2X1 U674 ( .A(n1001), .B(n1000), .Y(n90) );
  OAI22X1 U675 ( .A0(n464), .A1(n966), .B0(n964), .B1(n94), .Y(n473) );
  XOR2X1 U676 ( .A(B[18]), .B(n114), .Y(n608) );
  XOR2X1 U677 ( .A(B[18]), .B(n13), .Y(n327) );
  XOR2X1 U678 ( .A(B[18]), .B(n14), .Y(n471) );
  XOR2X1 U679 ( .A(B[18]), .B(n98), .Y(n248) );
  OAI22X1 U680 ( .A0(n461), .A1(n1042), .B0(n947), .B1(n99), .Y(n492) );
  OAI22X1 U681 ( .A0(n531), .A1(n947), .B0(n1042), .B1(n99), .Y(n534) );
  XNOR2X1 U682 ( .A(B[23]), .B(n905), .Y(n99) );
  AOI21X1 U683 ( .A0(n1024), .A1(n1022), .B0(n990), .Y(n991) );
  XNOR2X1 U684 ( .A(B[20]), .B(n905), .Y(n605) );
  OAI22X1 U685 ( .A0(n947), .A1(n151), .B0(n197), .B1(n1042), .Y(n200) );
  OAI22X1 U686 ( .A0(n947), .A1(n946), .B0(n945), .B1(n1042), .Y(n954) );
  OAI21XL U687 ( .A0(n1227), .A1(n1230), .B0(n1228), .Y(n104) );
  OAI21XL U688 ( .A0(n1235), .A1(n1238), .B0(n1236), .Y(n105) );
  OAI22X1 U689 ( .A0(n945), .A1(n947), .B0(n1042), .B1(n107), .Y(n843) );
  XOR2X1 U690 ( .A(n180), .B(n111), .Y(n829) );
  XOR2X1 U691 ( .A(n181), .B(n182), .Y(n111) );
  OAI22X1 U692 ( .A0(n947), .A1(n711), .B0(n675), .B1(n1042), .Y(n710) );
  AOI21XL U693 ( .A0(n628), .A1(n519), .B0(n518), .Y(n520) );
  ADDFHX1 U694 ( .A(n544), .B(n543), .CI(n542), .CO(n555), .S(n588) );
  INVX1 U695 ( .A(n698), .Y(n699) );
  OAI22X1 U696 ( .A0(n947), .A1(n605), .B0(n569), .B1(n1042), .Y(n604) );
  OAI22X1 U697 ( .A0(n966), .A1(n718), .B0(n964), .B1(n678), .Y(n732) );
  AOI21X1 U698 ( .A0(n346), .A1(n348), .B0(n309), .Y(n310) );
  CMPR22X1 U699 ( .A(n428), .B(n427), .CO(n435), .S(n468) );
  OAI22X1 U700 ( .A0(n713), .A1(n429), .B0(n392), .B1(n1042), .Y(n428) );
  CMPR22X1 U701 ( .A(n142), .B(n141), .CO(n138), .S(n834) );
  OAI22X1 U702 ( .A0(n947), .A1(n143), .B0(n152), .B1(n1042), .Y(n142) );
  XNOR2X4 U703 ( .A(n420), .B(n419), .Y(PRODUCT[29]) );
  OAI22X1 U704 ( .A0(n537), .A1(n536), .B0(n964), .B1(n495), .Y(n548) );
  OAI22X1 U705 ( .A0(n966), .A1(n160), .B0(n964), .B1(n159), .Y(n173) );
  XNOR2X1 U706 ( .A(n905), .B(B[14]), .Y(n151) );
  NAND2X1 U707 ( .A(n308), .B(n348), .Y(n311) );
  INVX1 U708 ( .A(n1048), .Y(n1020) );
  XOR2XL U709 ( .A(A[8]), .B(A[9]), .Y(n118) );
  XNOR2XL U710 ( .A(A[8]), .B(A[7]), .Y(n119) );
  NAND2X1 U711 ( .A(n118), .B(n119), .Y(n841) );
  XNOR2X1 U712 ( .A(n858), .B(B[5]), .Y(n158) );
  BUFX3 U713 ( .A(n119), .Y(n1061) );
  XOR2XL U714 ( .A(A[10]), .B(A[11]), .Y(n120) );
  BUFX3 U715 ( .A(n1110), .Y(n1083) );
  BUFX3 U716 ( .A(n1111), .Y(n1081) );
  OAI22XL U717 ( .A0(n1083), .A1(n137), .B0(n1081), .B1(n147), .Y(n164) );
  XOR2XL U718 ( .A(A[2]), .B(A[3]), .Y(n121) );
  XNOR2XL U719 ( .A(A[2]), .B(A[1]), .Y(n122) );
  NAND2X1 U720 ( .A(n121), .B(n122), .Y(n537) );
  BUFX3 U721 ( .A(n537), .Y(n966) );
  BUFX3 U722 ( .A(n122), .Y(n964) );
  OAI22XL U723 ( .A0(n966), .A1(n159), .B0(n964), .B1(n146), .Y(n163) );
  BUFX3 U724 ( .A(B[7]), .Y(n856) );
  XOR2XL U725 ( .A(A[14]), .B(A[15]), .Y(n124) );
  NAND2X1 U726 ( .A(n124), .B(n125), .Y(n641) );
  BUFX3 U727 ( .A(n641), .Y(n1152) );
  CLKINVX3 U728 ( .A(n98), .Y(n1148) );
  XNOR2XL U729 ( .A(n1148), .B(B[0]), .Y(n126) );
  BUFX3 U730 ( .A(n125), .Y(n1150) );
  XNOR2XL U731 ( .A(n1148), .B(B[1]), .Y(n198) );
  XOR2XL U732 ( .A(A[12]), .B(A[13]), .Y(n127) );
  BUFX3 U733 ( .A(n1140), .Y(n1114) );
  XNOR2XL U734 ( .A(n1102), .B(B[2]), .Y(n153) );
  BUFX3 U735 ( .A(n128), .Y(n1141) );
  XOR2XL U736 ( .A(A[4]), .B(A[5]), .Y(n129) );
  XNOR2XL U737 ( .A(A[4]), .B(A[3]), .Y(n130) );
  BUFX3 U738 ( .A(n898), .Y(n962) );
  BUFX3 U739 ( .A(n130), .Y(n960) );
  OAI22XL U740 ( .A0(n962), .A1(n161), .B0(n960), .B1(n149), .Y(n140) );
  XOR2XL U741 ( .A(A[6]), .B(A[7]), .Y(n131) );
  XNOR2XL U742 ( .A(A[6]), .B(A[5]), .Y(n132) );
  NAND2X1 U743 ( .A(n131), .B(n132), .Y(n580) );
  BUFX3 U744 ( .A(n580), .Y(n958) );
  BUFX3 U745 ( .A(n132), .Y(n956) );
  OAI22XL U746 ( .A0(n958), .A1(n135), .B0(n956), .B1(n148), .Y(n139) );
  NAND2X1 U747 ( .A(A[1]), .B(n133), .Y(n713) );
  BUFX3 U748 ( .A(n713), .Y(n947) );
  XNOR2X1 U749 ( .A(n905), .B(B[13]), .Y(n152) );
  BUFX3 U750 ( .A(n133), .Y(n1042) );
  OAI22X1 U751 ( .A0(n1114), .A1(n12), .B0(n1141), .B1(n134), .Y(n141) );
  OAI22X1 U752 ( .A0(n958), .A1(n145), .B0(n956), .B1(n135), .Y(n171) );
  XNOR2XL U753 ( .A(n1102), .B(B[0]), .Y(n136) );
  XNOR2XL U754 ( .A(n1102), .B(B[1]), .Y(n154) );
  XNOR2XL U755 ( .A(n1062), .B(B[2]), .Y(n144) );
  XNOR2XL U756 ( .A(n1062), .B(B[1]), .Y(n836) );
  OAI22X1 U757 ( .A0(n958), .A1(n835), .B0(n956), .B1(n145), .Y(n846) );
  XNOR2X1 U758 ( .A(n908), .B(B[9]), .Y(n838) );
  XNOR2X1 U759 ( .A(n908), .B(B[10]), .Y(n160) );
  OAI22XL U760 ( .A0(n966), .A1(n838), .B0(n964), .B1(n160), .Y(n845) );
  XNOR2X1 U761 ( .A(n895), .B(n856), .Y(n839) );
  OAI22XL U762 ( .A0(n962), .A1(n839), .B0(n960), .B1(n162), .Y(n844) );
  XNOR2X1 U763 ( .A(n908), .B(B[13]), .Y(n186) );
  OAI22XL U764 ( .A0(n966), .A1(n146), .B0(n964), .B1(n186), .Y(n185) );
  OAI22XL U765 ( .A0(n1083), .A1(n147), .B0(n1081), .B1(n189), .Y(n184) );
  OAI22XL U766 ( .A0(n962), .A1(n149), .B0(n960), .B1(n188), .Y(n196) );
  OAI22X1 U767 ( .A0(n1152), .A1(n98), .B0(n1150), .B1(n150), .Y(n199) );
  OAI22X1 U768 ( .A0(n947), .A1(n152), .B0(n151), .B1(n1042), .Y(n156) );
  ADDFHX1 U769 ( .A(n157), .B(n156), .CI(n155), .CO(n194), .S(n168) );
  BUFX3 U770 ( .A(n841), .Y(n1060) );
  OAI22XL U771 ( .A0(n1060), .A1(n175), .B0(n1061), .B1(n158), .Y(n174) );
  OAI22XL U772 ( .A0(n898), .A1(n162), .B0(n960), .B1(n161), .Y(n172) );
  CMPR32X1 U773 ( .A(n168), .B(n167), .C(n166), .CO(n191), .S(n831) );
  CMPR32X1 U774 ( .A(n171), .B(n170), .C(n169), .CO(n182), .S(n849) );
  ADDFHX1 U775 ( .A(n174), .B(n173), .CI(n172), .CO(n167), .S(n848) );
  XNOR2X1 U776 ( .A(n905), .B(B[10]), .Y(n945) );
  OAI22X1 U777 ( .A0(n1083), .A1(n13), .B0(n1081), .B1(n176), .Y(n842) );
  NAND2XL U778 ( .A(n822), .B(n821), .Y(mult_x_1_n313) );
  CMPR32X1 U779 ( .A(n185), .B(n184), .C(n183), .CO(n789), .S(n193) );
  XNOR2X1 U780 ( .A(n908), .B(B[14]), .Y(n719) );
  OAI22XL U781 ( .A0(n966), .A1(n186), .B0(n964), .B1(n719), .Y(n755) );
  OAI22XL U782 ( .A0(n962), .A1(n188), .B0(n960), .B1(n726), .Y(n762) );
  XNOR2X1 U783 ( .A(n1062), .B(B[6]), .Y(n728) );
  OAI22XL U784 ( .A0(n1083), .A1(n189), .B0(n1081), .B1(n728), .Y(n761) );
  CMPR32X1 U785 ( .A(n196), .B(n195), .C(n194), .CO(n801), .S(n192) );
  XNOR2XL U786 ( .A(n1148), .B(B[2]), .Y(n715) );
  OAI22X1 U787 ( .A0(n1152), .A1(n198), .B0(n1150), .B1(n715), .Y(n752) );
  CMPR22X1 U788 ( .A(n200), .B(n199), .CO(n782), .S(n195) );
  CMPR32X1 U789 ( .A(n203), .B(n202), .C(n201), .CO(n781), .S(n205) );
  CMPR32X1 U790 ( .A(n209), .B(n208), .C(n207), .CO(n210), .S(n822) );
  NAND2XL U791 ( .A(n242), .B(n235), .Y(n218) );
  NAND2XL U792 ( .A(n213), .B(n1091), .Y(n221) );
  OAI21XL U793 ( .A0(n1219), .A1(n1222), .B0(n1220), .Y(n214) );
  OAI21XL U794 ( .A0(n1215), .A1(n1218), .B0(n1216), .Y(n226) );
  AOI21XL U795 ( .A0(n1195), .A1(n1091), .B0(n1094), .Y(n220) );
  OAI21XL U796 ( .A0(n1198), .A1(n221), .B0(n220), .Y(n223) );
  INVX1 U797 ( .A(n347), .Y(n308) );
  INVXL U798 ( .A(n224), .Y(n278) );
  INVXL U799 ( .A(n1213), .Y(n282) );
  NAND2XL U800 ( .A(n282), .B(n242), .Y(n230) );
  NOR2XL U801 ( .A(n278), .B(n230), .Y(n232) );
  NAND2XL U802 ( .A(n308), .B(n232), .Y(n234) );
  AOI21XL U803 ( .A0(n228), .A1(n242), .B0(n227), .Y(n229) );
  OAI21XL U804 ( .A0(n279), .A1(n230), .B0(n229), .Y(n231) );
  AOI21XL U805 ( .A0(n346), .A1(n232), .B0(n231), .Y(n233) );
  OAI21XL U806 ( .A0(n1198), .A1(n234), .B0(n233), .Y(n237) );
  XNOR2X1 U807 ( .A(n237), .B(n236), .Y(PRODUCT[35]) );
  NOR2XL U808 ( .A(n278), .B(n1213), .Y(n239) );
  NAND2XL U809 ( .A(n308), .B(n239), .Y(n241) );
  OAI21XL U810 ( .A0(n279), .A1(n1213), .B0(n1214), .Y(n238) );
  AOI21XL U811 ( .A0(n346), .A1(n239), .B0(n238), .Y(n240) );
  XNOR2X2 U812 ( .A(n244), .B(n243), .Y(PRODUCT[34]) );
  XNOR2X1 U813 ( .A(A[15]), .B(B[17]), .Y(n245) );
  XNOR2X1 U814 ( .A(A[15]), .B(B[16]), .Y(n288) );
  XNOR2X1 U815 ( .A(n895), .B(n1147), .Y(n246) );
  XNOR2X1 U816 ( .A(A[9]), .B(B[23]), .Y(n285) );
  XNOR2X1 U817 ( .A(A[9]), .B(B[24]), .Y(n253) );
  OAI22XL U818 ( .A0(n1060), .A1(n285), .B0(n1061), .B1(n253), .Y(n258) );
  INVXL U819 ( .A(n268), .Y(n257) );
  OAI22X1 U820 ( .A0(n1152), .A1(n248), .B0(n1150), .B1(n264), .Y(n269) );
  OAI22XL U821 ( .A0(n1110), .A1(n252), .B0(n1081), .B1(n266), .Y(n271) );
  OAI22XL U822 ( .A0(n1083), .A1(n286), .B0(n1081), .B1(n256), .Y(n291) );
  CMPR32X1 U823 ( .A(n259), .B(n258), .C(n257), .CO(n275), .S(n301) );
  CMPR32X1 U824 ( .A(n262), .B(n261), .C(n260), .CO(n305), .S(n300) );
  OAI22X1 U825 ( .A0(n1060), .A1(n265), .B0(n1061), .B1(n1058), .Y(n1077) );
  CMPR32X1 U826 ( .A(n269), .B(n268), .C(n267), .CO(n1069), .S(n274) );
  CMPR32X1 U827 ( .A(n272), .B(n271), .C(n270), .CO(n1068), .S(n273) );
  CMPR32X1 U828 ( .A(n275), .B(n274), .C(n273), .CO(n1054), .S(n304) );
  NOR2XL U829 ( .A(n277), .B(n276), .Y(mult_x_1_n162) );
  NAND2XL U830 ( .A(n277), .B(n276), .Y(mult_x_1_n163) );
  NAND2XL U831 ( .A(n308), .B(n224), .Y(n281) );
  AOI21XL U832 ( .A0(n346), .A1(n224), .B0(n226), .Y(n280) );
  NAND2X1 U833 ( .A(n282), .B(n1214), .Y(n283) );
  XNOR2X4 U834 ( .A(n284), .B(n283), .Y(PRODUCT[33]) );
  XNOR2X1 U835 ( .A(A[9]), .B(B[22]), .Y(n290) );
  XNOR2X1 U836 ( .A(n1062), .B(B[19]), .Y(n326) );
  OAI22XL U837 ( .A0(n1110), .A1(n326), .B0(n1081), .B1(n286), .Y(n322) );
  INVXL U838 ( .A(n295), .Y(n320) );
  OAI22XL U839 ( .A0(n1152), .A1(n314), .B0(n1150), .B1(n288), .Y(n319) );
  OAI22XL U840 ( .A0(n1140), .A1(n324), .B0(n1141), .B1(n289), .Y(n318) );
  CMPR32X1 U841 ( .A(n293), .B(n292), .C(n291), .CO(n302), .S(n340) );
  CMPR32X1 U842 ( .A(n296), .B(n295), .C(n294), .CO(n260), .S(n339) );
  CMPR32X1 U843 ( .A(n305), .B(n304), .C(n303), .CO(n277), .S(n306) );
  NOR2XL U844 ( .A(n307), .B(n306), .Y(mult_x_1_n173) );
  NAND2XL U845 ( .A(n307), .B(n306), .Y(mult_x_1_n174) );
  OAI22XL U846 ( .A0(n1152), .A1(n330), .B0(n1150), .B1(n314), .Y(n334) );
  XNOR2X1 U847 ( .A(n908), .B(n1147), .Y(n315) );
  INVXL U848 ( .A(n315), .Y(n316) );
  CMPR32X1 U849 ( .A(n319), .B(n318), .C(n317), .CO(n297), .S(n354) );
  CMPR32X1 U850 ( .A(n322), .B(n321), .C(n320), .CO(n298), .S(n353) );
  OAI22XL U851 ( .A0(n962), .A1(n328), .B0(n960), .B1(n323), .Y(n337) );
  OAI22XL U852 ( .A0(n1114), .A1(n356), .B0(n1141), .B1(n324), .Y(n336) );
  XNOR2X1 U853 ( .A(A[9]), .B(B[20]), .Y(n331) );
  OAI22XL U854 ( .A0(n1060), .A1(n331), .B0(n1061), .B1(n325), .Y(n364) );
  OAI22XL U855 ( .A0(n1110), .A1(n327), .B0(n1081), .B1(n326), .Y(n363) );
  XNOR2X1 U856 ( .A(n1062), .B(B[17]), .Y(n366) );
  OAI22X1 U857 ( .A0(n1083), .A1(n366), .B0(n1081), .B1(n327), .Y(n370) );
  XNOR2X1 U858 ( .A(n895), .B(B[23]), .Y(n367) );
  OAI22X1 U859 ( .A0(n962), .A1(n367), .B0(n960), .B1(n328), .Y(n369) );
  INVXL U860 ( .A(n333), .Y(n368) );
  XNOR2X1 U861 ( .A(n1148), .B(B[13]), .Y(n360) );
  XNOR2X1 U862 ( .A(A[9]), .B(B[19]), .Y(n359) );
  CMPR32X1 U863 ( .A(n337), .B(n336), .C(n335), .CO(n376), .S(n389) );
  CMPR32X1 U864 ( .A(n343), .B(n342), .C(n341), .CO(n307), .S(n344) );
  NOR2XL U865 ( .A(n345), .B(n344), .Y(mult_x_1_n184) );
  NAND2XL U866 ( .A(n345), .B(n344), .Y(mult_x_1_n185) );
  CMPR32X1 U867 ( .A(n352), .B(n351), .C(n350), .CO(n345), .S(n378) );
  CMPR32X1 U868 ( .A(n355), .B(n354), .C(n353), .CO(n352), .S(n388) );
  XNOR2X1 U869 ( .A(B[15]), .B(n1102), .Y(n358) );
  OAI22X1 U870 ( .A0(n958), .A1(n404), .B0(n956), .B1(n357), .Y(n395) );
  OR2X2 U871 ( .A(n395), .B(n394), .Y(n400) );
  CMPR32X1 U872 ( .A(n364), .B(n363), .C(n362), .CO(n375), .S(n412) );
  OAI22X1 U873 ( .A0(n966), .A1(n397), .B0(n964), .B1(n365), .Y(n410) );
  XNOR2X1 U874 ( .A(n1062), .B(B[16]), .Y(n403) );
  OAI22XL U875 ( .A0(n962), .A1(n402), .B0(n960), .B1(n367), .Y(n408) );
  NOR2XL U876 ( .A(n378), .B(n377), .Y(mult_x_1_n191) );
  NAND2XL U877 ( .A(n378), .B(n377), .Y(mult_x_1_n192) );
  INVXL U878 ( .A(n379), .Y(n417) );
  CMPR32X1 U879 ( .A(n391), .B(n390), .C(n389), .CO(n374), .S(n423) );
  XNOR2X1 U880 ( .A(n395), .B(n394), .Y(n434) );
  CMPR32X1 U881 ( .A(n401), .B(n400), .C(n399), .CO(n413), .S(n446) );
  OAI22XL U882 ( .A0(n1083), .A1(n437), .B0(n1081), .B1(n403), .Y(n443) );
  OAI22XL U883 ( .A0(n958), .A1(n438), .B0(n956), .B1(n404), .Y(n442) );
  CMPR32X1 U884 ( .A(n410), .B(n409), .C(n408), .CO(n426), .S(n456) );
  OAI21X2 U885 ( .A0(n1198), .A1(n417), .B0(n416), .Y(n420) );
  NAND2X1 U886 ( .A(n418), .B(n1222), .Y(n419) );
  CMPR32X1 U887 ( .A(n423), .B(n422), .C(n421), .CO(n414), .S(n449) );
  CMPR32X1 U888 ( .A(n426), .B(n425), .C(n424), .CO(n411), .S(n455) );
  XNOR2X1 U889 ( .A(n1148), .B(B[10]), .Y(n462) );
  OAI22XL U890 ( .A0(n641), .A1(n462), .B0(n1150), .B1(n430), .Y(n459) );
  XNOR2X1 U891 ( .A(A[9]), .B(B[16]), .Y(n463) );
  CMPR32X1 U892 ( .A(n435), .B(n434), .C(n433), .CO(n447), .S(n479) );
  XNOR2X1 U893 ( .A(n895), .B(B[20]), .Y(n469) );
  OAI22XL U894 ( .A0(n1083), .A1(n470), .B0(n1081), .B1(n437), .Y(n476) );
  ADDFHX1 U895 ( .A(n441), .B(n440), .CI(n439), .CO(n433), .S(n489) );
  CMPR32X1 U896 ( .A(n444), .B(n443), .C(n442), .CO(n458), .S(n488) );
  NOR2XL U897 ( .A(n449), .B(n448), .Y(mult_x_1_n209) );
  NAND2XL U898 ( .A(n449), .B(n448), .Y(mult_x_1_n210) );
  INVXL U899 ( .A(n1223), .Y(n450) );
  NAND2X1 U900 ( .A(n450), .B(n1224), .Y(n451) );
  XNOR2X4 U901 ( .A(n452), .B(n451), .Y(PRODUCT[28]) );
  CMPR32X1 U902 ( .A(n455), .B(n454), .C(n453), .CO(n448), .S(n482) );
  CMPR32X1 U903 ( .A(n458), .B(n457), .C(n456), .CO(n445), .S(n487) );
  ADDHXL U904 ( .A(n460), .B(n459), .CO(n467), .S(n499) );
  XNOR2X1 U905 ( .A(A[9]), .B(B[15]), .Y(n494) );
  OAI22XL U906 ( .A0(n1060), .A1(n494), .B0(n1061), .B1(n463), .Y(n505) );
  XNOR2X1 U907 ( .A(n908), .B(B[21]), .Y(n495) );
  XNOR2X1 U908 ( .A(n895), .B(B[19]), .Y(n500) );
  OAI22X1 U909 ( .A0(n962), .A1(n500), .B0(n960), .B1(n469), .Y(n508) );
  XNOR2X1 U910 ( .A(n1062), .B(B[13]), .Y(n501) );
  OAI22XL U911 ( .A0(n580), .A1(n502), .B0(n956), .B1(n471), .Y(n506) );
  CMPR32X1 U912 ( .A(n477), .B(n476), .C(n475), .CO(n490), .S(n528) );
  NOR2XL U913 ( .A(n482), .B(n481), .Y(mult_x_1_n220) );
  NAND2XL U914 ( .A(n482), .B(n481), .Y(mult_x_1_n221) );
  INVXL U915 ( .A(n1225), .Y(n483) );
  XOR2X2 U916 ( .A(n1198), .B(n484), .Y(PRODUCT[27]) );
  CMPR32X1 U917 ( .A(n490), .B(n489), .C(n488), .CO(n478), .S(n527) );
  CMPR22X1 U918 ( .A(n492), .B(n491), .CO(n498), .S(n544) );
  XNOR2X1 U919 ( .A(n905), .B(B[22]), .Y(n531) );
  OAI22XL U920 ( .A0(n1060), .A1(n535), .B0(n1061), .B1(n494), .Y(n549) );
  OAI22XL U921 ( .A0(n580), .A1(n546), .B0(n956), .B1(n502), .Y(n550) );
  NOR2XL U922 ( .A(n513), .B(n512), .Y(mult_x_1_n223) );
  NAND2XL U923 ( .A(n519), .B(n627), .Y(n521) );
  OAI21XL U924 ( .A0(n11), .A1(n1229), .B0(n1230), .Y(n518) );
  CMPR32X1 U925 ( .A(n530), .B(n529), .C(n528), .CO(n509), .S(n563) );
  OAI22X1 U926 ( .A0(n947), .A1(n569), .B0(n531), .B1(n1042), .Y(n568) );
  CMPR22X1 U927 ( .A(n534), .B(n533), .CO(n543), .S(n576) );
  OR2X2 U928 ( .A(n575), .B(n576), .Y(n539) );
  XNOR2X1 U929 ( .A(n858), .B(B[13]), .Y(n571) );
  OAI22XL U930 ( .A0(n1060), .A1(n571), .B0(n1061), .B1(n535), .Y(n583) );
  XNOR2X1 U931 ( .A(n908), .B(B[19]), .Y(n572) );
  OAI22X1 U932 ( .A0(n537), .A1(n572), .B0(n964), .B1(n536), .Y(n582) );
  OAI22X1 U933 ( .A0(n958), .A1(n579), .B0(n956), .B1(n546), .Y(n584) );
  ADDFHX1 U934 ( .A(n549), .B(n548), .CI(n547), .CO(n542), .S(n601) );
  NOR2XL U935 ( .A(n557), .B(n556), .Y(mult_x_1_n232) );
  NAND2XL U936 ( .A(n627), .B(n514), .Y(n559) );
  CMPR32X1 U937 ( .A(n563), .B(n562), .C(n561), .CO(n556), .S(n591) );
  CMPR32X1 U938 ( .A(n566), .B(n565), .C(n564), .CO(n553), .S(n599) );
  CMPR22X1 U939 ( .A(n568), .B(n567), .CO(n575), .S(n612) );
  OAI22XL U940 ( .A0(n1060), .A1(n607), .B0(n1061), .B1(n571), .Y(n618) );
  OAI22X1 U941 ( .A0(n966), .A1(n608), .B0(n964), .B1(n572), .Y(n617) );
  OAI22X1 U942 ( .A0(n1114), .A1(n609), .B0(n1141), .B1(n573), .Y(n616) );
  XOR3X2 U943 ( .A(n576), .B(n575), .C(n574), .Y(n623) );
  OAI22X1 U944 ( .A0(n962), .A1(n613), .B0(n960), .B1(n577), .Y(n621) );
  XNOR2X1 U945 ( .A(n1062), .B(B[10]), .Y(n614) );
  CMPR32X1 U946 ( .A(n589), .B(n588), .C(n587), .CO(n562), .S(n597) );
  NOR2XL U947 ( .A(n591), .B(n590), .Y(mult_x_1_n241) );
  NAND2XL U948 ( .A(n591), .B(n590), .Y(mult_x_1_n242) );
  CMPR32X1 U949 ( .A(n602), .B(n601), .C(n600), .CO(n587), .S(n633) );
  CMPR22X1 U950 ( .A(n604), .B(n603), .CO(n611), .S(n647) );
  XNOR2X1 U951 ( .A(n905), .B(B[19]), .Y(n639) );
  OAI22X1 U952 ( .A0(n947), .A1(n639), .B0(n605), .B1(n1042), .Y(n638) );
  OAI22X1 U953 ( .A0(n1152), .A1(n640), .B0(n1150), .B1(n606), .Y(n637) );
  OAI22XL U954 ( .A0(n962), .A1(n648), .B0(n960), .B1(n613), .Y(n655) );
  OAI22XL U955 ( .A0(n1083), .A1(n649), .B0(n1081), .B1(n614), .Y(n654) );
  CMPR32X1 U956 ( .A(n618), .B(n617), .C(n616), .CO(n610), .S(n671) );
  CMPR32X1 U957 ( .A(n624), .B(n623), .C(n622), .CO(n598), .S(n631) );
  NOR2XL U958 ( .A(n626), .B(n625), .Y(mult_x_1_n252) );
  NAND2XL U959 ( .A(n626), .B(n625), .Y(mult_x_1_n253) );
  CMPR32X1 U960 ( .A(n633), .B(n632), .C(n631), .CO(n625), .S(n660) );
  CMPR32X1 U961 ( .A(n636), .B(n635), .C(n634), .CO(n622), .S(n669) );
  CMPR22X1 U962 ( .A(n638), .B(n637), .CO(n646), .S(n682) );
  OAI22X1 U963 ( .A0(n947), .A1(n675), .B0(n639), .B1(n1042), .Y(n674) );
  OAI22X1 U964 ( .A0(n641), .A1(n676), .B0(n1150), .B1(n640), .Y(n673) );
  XNOR2X1 U965 ( .A(n858), .B(B[10]), .Y(n677) );
  XNOR2X1 U966 ( .A(n908), .B(B[16]), .Y(n678) );
  XNOR2X1 U967 ( .A(n895), .B(B[14]), .Y(n683) );
  OAI22XL U968 ( .A0(n962), .A1(n683), .B0(n960), .B1(n648), .Y(n691) );
  OAI22XL U969 ( .A0(n1083), .A1(n684), .B0(n1081), .B1(n649), .Y(n690) );
  CMPR32X1 U970 ( .A(n655), .B(n654), .C(n653), .CO(n672), .S(n706) );
  NAND2XL U971 ( .A(n660), .B(n659), .Y(mult_x_1_n260) );
  NAND2XL U972 ( .A(n697), .B(n662), .Y(n664) );
  CMPR32X1 U973 ( .A(n672), .B(n671), .C(n670), .CO(n656), .S(n705) );
  CMPR22X1 U974 ( .A(n674), .B(n673), .CO(n681), .S(n724) );
  OAI22X1 U975 ( .A0(n1152), .A1(n714), .B0(n1150), .B1(n676), .Y(n709) );
  XNOR2X1 U976 ( .A(n858), .B(B[9]), .Y(n716) );
  OAI22XL U977 ( .A0(n1060), .A1(n716), .B0(n1061), .B1(n677), .Y(n733) );
  XNOR2X1 U978 ( .A(n908), .B(B[15]), .Y(n718) );
  XNOR2X1 U979 ( .A(n895), .B(B[13]), .Y(n725) );
  OAI22XL U980 ( .A0(n962), .A1(n725), .B0(n960), .B1(n683), .Y(n736) );
  XNOR2X1 U981 ( .A(n1062), .B(n856), .Y(n727) );
  OAI22XL U982 ( .A0(n1083), .A1(n727), .B0(n1081), .B1(n684), .Y(n735) );
  CMPR32X1 U983 ( .A(n691), .B(n690), .C(n689), .CO(n708), .S(n747) );
  NOR2XL U984 ( .A(n696), .B(n695), .Y(mult_x_1_n270) );
  NAND2XL U985 ( .A(n696), .B(n695), .Y(mult_x_1_n271) );
  CMPR32X1 U986 ( .A(n705), .B(n704), .C(n703), .CO(n695), .S(n741) );
  CMPR22X1 U987 ( .A(n710), .B(n709), .CO(n723), .S(n759) );
  OAI22X1 U988 ( .A0(n713), .A1(n712), .B0(n711), .B1(n1042), .Y(n751) );
  OAI22X1 U989 ( .A0(n1152), .A1(n715), .B0(n1150), .B1(n714), .Y(n750) );
  OAI22XL U990 ( .A0(n841), .A1(n717), .B0(n1061), .B1(n716), .Y(n765) );
  OAI22XL U991 ( .A0(n966), .A1(n719), .B0(n964), .B1(n718), .Y(n764) );
  CMPR32X1 U992 ( .A(n724), .B(n723), .C(n722), .CO(n739), .S(n770) );
  OAI22XL U993 ( .A0(n962), .A1(n726), .B0(n960), .B1(n725), .Y(n768) );
  OAI22XL U994 ( .A0(n1083), .A1(n728), .B0(n1081), .B1(n727), .Y(n767) );
  CMPR32X1 U995 ( .A(n733), .B(n732), .C(n731), .CO(n722), .S(n779) );
  CMPR32X1 U996 ( .A(n736), .B(n735), .C(n734), .CO(n749), .S(n778) );
  CMPR32X1 U997 ( .A(n739), .B(n738), .C(n737), .CO(n704), .S(n744) );
  NOR2XL U998 ( .A(n741), .B(n740), .Y(mult_x_1_n277) );
  NAND2XL U999 ( .A(n741), .B(n740), .Y(mult_x_1_n278) );
  CMPR32X1 U1000 ( .A(n746), .B(n745), .C(n744), .CO(n740), .S(n773) );
  CMPR22X1 U1001 ( .A(n753), .B(n752), .CO(n785), .S(n783) );
  CMPR32X1 U1002 ( .A(n756), .B(n755), .C(n754), .CO(n784), .S(n788) );
  CMPR32X1 U1003 ( .A(n762), .B(n761), .C(n760), .CO(n798), .S(n787) );
  CMPR32X1 U1004 ( .A(n765), .B(n764), .C(n763), .CO(n757), .S(n797) );
  CMPR32X1 U1005 ( .A(n768), .B(n767), .C(n766), .CO(n780), .S(n796) );
  NOR2XL U1006 ( .A(n773), .B(n772), .Y(mult_x_1_n288) );
  NAND2XL U1007 ( .A(n773), .B(n772), .Y(mult_x_1_n289) );
  CMPR32X1 U1008 ( .A(n780), .B(n779), .C(n778), .CO(n769), .S(n810) );
  CMPR32X1 U1009 ( .A(n783), .B(n782), .C(n781), .CO(n804), .S(n800) );
  CMPR32X1 U1010 ( .A(n789), .B(n788), .C(n787), .CO(n802), .S(n807) );
  NOR2XL U1011 ( .A(n794), .B(n793), .Y(mult_x_1_n291) );
  NAND2XL U1012 ( .A(n794), .B(n793), .Y(mult_x_1_n292) );
  INVXL U1013 ( .A(n1244), .Y(n795) );
  CMPR32X1 U1014 ( .A(n798), .B(n797), .C(n796), .CO(n790), .S(n813) );
  NOR2XL U1015 ( .A(mult_x_1_n302), .B(mult_x_1_n299), .Y(mult_x_1_n297) );
  NAND2XL U1016 ( .A(n815), .B(n814), .Y(mult_x_1_n300) );
  NAND2XL U1017 ( .A(n818), .B(n817), .Y(mult_x_1_n303) );
  INVXL U1018 ( .A(n1251), .Y(n819) );
  XOR2X1 U1019 ( .A(n820), .B(n1249), .Y(PRODUCT[16]) );
  NOR2XL U1020 ( .A(n823), .B(mult_x_1_n312), .Y(mult_x_1_n305) );
  NAND2XL U1021 ( .A(n825), .B(n824), .Y(mult_x_1_n78) );
  NAND2XL U1022 ( .A(n826), .B(n1251), .Y(n827) );
  XNOR2X1 U1023 ( .A(n828), .B(n827), .Y(PRODUCT[15]) );
  XNOR2X1 U1024 ( .A(n1256), .B(n1252), .Y(PRODUCT[14]) );
  CMPR32X1 U1025 ( .A(n834), .B(n833), .C(n832), .CO(n180), .S(n995) );
  XNOR2XL U1026 ( .A(n1062), .B(B[0]), .Y(n837) );
  OAI22XL U1027 ( .A0(n898), .A1(n959), .B0(n960), .B1(n839), .Y(n942) );
  XNOR2XL U1028 ( .A(n858), .B(B[2]), .Y(n948) );
  OAI22X1 U1029 ( .A0(n841), .A1(n948), .B0(n1061), .B1(n840), .Y(n941) );
  CMPR22X1 U1030 ( .A(n843), .B(n842), .CO(n997), .S(n940) );
  CMPR32X1 U1031 ( .A(n846), .B(n845), .C(n844), .CO(n832), .S(n1002) );
  CMPR32X1 U1032 ( .A(n849), .B(n848), .C(n847), .CO(n830), .S(n993) );
  INVXL U1033 ( .A(n1045), .Y(n852) );
  NAND2XL U1034 ( .A(n852), .B(n1044), .Y(mult_x_1_n80) );
  XNOR2X1 U1035 ( .A(n1257), .B(n1253), .Y(PRODUCT[13]) );
  XNOR2XL U1036 ( .A(n866), .B(B[2]), .Y(n861) );
  OAI22XL U1037 ( .A0(n958), .A1(n861), .B0(n956), .B1(n957), .Y(n952) );
  XNOR2XL U1038 ( .A(n858), .B(B[0]), .Y(n853) );
  XNOR2XL U1039 ( .A(n858), .B(B[1]), .Y(n949) );
  XNOR2X1 U1040 ( .A(n908), .B(B[6]), .Y(n857) );
  OAI22XL U1041 ( .A0(n966), .A1(n869), .B0(n964), .B1(n857), .Y(n872) );
  OAI22XL U1042 ( .A0(n898), .A1(n865), .B0(n960), .B1(n854), .Y(n871) );
  XNOR2X1 U1043 ( .A(n905), .B(B[6]), .Y(n881) );
  XNOR2X1 U1044 ( .A(n905), .B(B[8]), .Y(n860) );
  XNOR2X1 U1045 ( .A(n905), .B(B[9]), .Y(n946) );
  OAI22X1 U1046 ( .A0(n947), .A1(n860), .B0(n946), .B1(n1042), .Y(n944) );
  OAI22X1 U1047 ( .A0(n1060), .A1(n97), .B0(n1061), .B1(n859), .Y(n943) );
  XNOR2XL U1048 ( .A(n866), .B(B[1]), .Y(n867) );
  CMPR32X1 U1049 ( .A(n864), .B(n863), .C(n862), .CO(n973), .S(n875) );
  XNOR2XL U1050 ( .A(n895), .B(B[2]), .Y(n882) );
  OAI22X1 U1051 ( .A0(n962), .A1(n882), .B0(n960), .B1(n865), .Y(n880) );
  XNOR2XL U1052 ( .A(n866), .B(B[0]), .Y(n868) );
  OAI22X1 U1053 ( .A0(n958), .A1(n868), .B0(n956), .B1(n867), .Y(n879) );
  OAI22XL U1054 ( .A0(n966), .A1(n886), .B0(n964), .B1(n869), .Y(n878) );
  CMPR32X1 U1055 ( .A(n872), .B(n871), .C(n870), .CO(n983), .S(n873) );
  ADDHXL U1056 ( .A(n877), .B(n876), .CO(n870), .S(n885) );
  CMPR32X1 U1057 ( .A(n880), .B(n879), .C(n878), .CO(n874), .S(n884) );
  XNOR2XL U1058 ( .A(n895), .B(B[1]), .Y(n896) );
  CMPR32X1 U1059 ( .A(n883), .B(n884), .C(n885), .CO(n936), .S(n934) );
  CMPR32X1 U1060 ( .A(n890), .B(n889), .C(n888), .CO(n883), .S(n891) );
  NOR2X1 U1061 ( .A(n934), .B(n933), .Y(n935) );
  XNOR2XL U1062 ( .A(n908), .B(B[2]), .Y(n916) );
  XNOR2XL U1063 ( .A(n895), .B(B[0]), .Y(n897) );
  ADDHXL U1064 ( .A(n900), .B(n899), .CO(n892), .S(n922) );
  OR2X2 U1065 ( .A(n932), .B(n931), .Y(n1165) );
  XNOR2XL U1066 ( .A(n905), .B(B[1]), .Y(n901) );
  XNOR2XL U1067 ( .A(n905), .B(B[2]), .Y(n906) );
  OAI21XL U1068 ( .A0(n1176), .A1(n1182), .B0(n1177), .Y(n1174) );
  OAI22X1 U1069 ( .A0(n947), .A1(n906), .B0(n915), .B1(n1042), .Y(n919) );
  XNOR2XL U1070 ( .A(n908), .B(B[0]), .Y(n907) );
  XNOR2XL U1071 ( .A(n908), .B(B[1]), .Y(n917) );
  OAI22X1 U1072 ( .A0(n966), .A1(n907), .B0(n964), .B1(n917), .Y(n918) );
  CMPR22X1 U1073 ( .A(n919), .B(n918), .CO(n920), .S(n912) );
  OAI21XL U1074 ( .A0(n1171), .A1(n1168), .B0(n1169), .Y(n1186) );
  CMPR32X1 U1075 ( .A(n924), .B(n923), .C(n922), .CO(n931), .S(n929) );
  CMPR32X1 U1076 ( .A(n927), .B(n926), .C(n925), .CO(n928), .S(n921) );
  OR2X2 U1077 ( .A(n929), .B(n928), .Y(n1185) );
  ADDFHX1 U1078 ( .A(n942), .B(n941), .CI(n940), .CO(n1003), .S(n1010) );
  CMPR22X1 U1079 ( .A(n944), .B(n943), .CO(n978), .S(n974) );
  ADDFHX1 U1080 ( .A(n955), .B(n954), .CI(n953), .CO(n1001), .S(n977) );
  OAI22X1 U1081 ( .A0(n962), .A1(n961), .B0(n960), .B1(n959), .Y(n971) );
  OAI22XL U1082 ( .A0(n966), .A1(n965), .B0(n964), .B1(n963), .Y(n970) );
  CMPR32X1 U1083 ( .A(n969), .B(n968), .C(n967), .CO(n1004), .S(n999) );
  ADDFHX1 U1084 ( .A(n978), .B(n977), .CI(n976), .CO(n1009), .S(n979) );
  CMPR32X1 U1085 ( .A(n981), .B(n980), .C(n979), .CO(n988), .S(n987) );
  CMPR32X1 U1086 ( .A(n984), .B(n983), .C(n982), .CO(n986), .S(n939) );
  NOR2XL U1087 ( .A(n987), .B(n986), .Y(n985) );
  NAND2XL U1088 ( .A(n1024), .B(n1028), .Y(n992) );
  NAND2XL U1089 ( .A(n989), .B(n988), .Y(n1023) );
  INVXL U1090 ( .A(n1023), .Y(n990) );
  OAI21X1 U1091 ( .A0(n1021), .A1(n992), .B0(n991), .Y(n1048) );
  CMPR32X1 U1092 ( .A(n998), .B(n997), .C(n996), .CO(n847), .S(n1007) );
  CMPR32X1 U1093 ( .A(n1004), .B(n1003), .C(n1002), .CO(n994), .S(n1005) );
  CMPR32X1 U1094 ( .A(n1007), .B(n1006), .C(n1005), .CO(n1014), .S(n1013) );
  NAND2XL U1095 ( .A(n1090), .B(n1018), .Y(n1043) );
  INVXL U1096 ( .A(n1016), .Y(n1019) );
  OAI21XL U1097 ( .A0(n1020), .A1(n1043), .B0(n1046), .Y(mult_x_1_n320) );
  NAND2XL U1098 ( .A(n1018), .B(n1016), .Y(n1017) );
  OAI21XL U1099 ( .A0(n1020), .A1(n1011), .B0(n1016), .Y(mult_x_1_n327) );
  AOI21X1 U1100 ( .A0(n1030), .A1(n1028), .B0(n1022), .Y(n1026) );
  NAND2XL U1101 ( .A(n1024), .B(n1023), .Y(n1025) );
  XOR2X1 U1102 ( .A(n1026), .B(n1025), .Y(n1273) );
  NAND2XL U1103 ( .A(n1028), .B(n1027), .Y(n1029) );
  OAI21XL U1104 ( .A0(n1041), .A1(n1037), .B0(n1038), .Y(n1036) );
  INVXL U1105 ( .A(n1032), .Y(n1034) );
  INVXL U1106 ( .A(n1037), .Y(n1039) );
  NOR2XL U1107 ( .A(n1043), .B(n1045), .Y(n1049) );
  OAI21XL U1108 ( .A0(n1046), .A1(n1045), .B0(n1044), .Y(n1047) );
  AOI21XL U1109 ( .A0(n1049), .A1(n1048), .B0(n1047), .Y(mult_x_1_n315) );
  OAI21XL U1110 ( .A0(n1198), .A1(n1051), .B0(n1050), .Y(n1053) );
  CMPR32X1 U1111 ( .A(n1067), .B(n1066), .C(n1065), .CO(n1084), .S(n1056) );
  CMPR32X1 U1112 ( .A(n1070), .B(n1069), .C(n1068), .CO(n1073), .S(n1055) );
  CMPR32X1 U1113 ( .A(n1078), .B(n1077), .C(n1076), .CO(n1122), .S(n1075) );
  OAI22X1 U1114 ( .A0(n1083), .A1(n1082), .B0(n1081), .B1(n1108), .Y(n1117) );
  CMPR32X1 U1115 ( .A(n1086), .B(n1085), .C(n1084), .CO(n1120), .S(n1074) );
  NAND2XL U1116 ( .A(n1090), .B(n1089), .Y(mult_x_1_n81) );
  OAI21XL U1117 ( .A0(n1198), .A1(n1098), .B0(n1097), .Y(n1101) );
  CMPR32X1 U1118 ( .A(n1106), .B(n1105), .C(n1104), .CO(n1124), .S(n1121) );
  OAI22X1 U1119 ( .A0(n1114), .A1(n1113), .B0(n1141), .B1(n1138), .Y(n1146) );
  CMPR32X1 U1120 ( .A(n1117), .B(n1116), .C(n1115), .CO(n1134), .S(n1123) );
  CMPR32X1 U1121 ( .A(n1122), .B(n1121), .C(n1120), .CO(n1127), .S(n1087) );
  CMPR32X1 U1122 ( .A(n1125), .B(n1124), .C(n1123), .CO(n1119), .S(n1126) );
  OAI21XL U1123 ( .A0(n1129), .A1(n1203), .B0(n1204), .Y(n1191) );
  OAI21XL U1124 ( .A0(n1198), .A1(n1131), .B0(n1130), .Y(n1133) );
  CMPR32X1 U1125 ( .A(n1136), .B(n1135), .C(n1134), .CO(n1143), .S(n1118) );
  CMPR32X1 U1126 ( .A(n1146), .B(n1145), .C(n1144), .CO(n1155), .S(n1142) );
  XNOR2XL U1127 ( .A(n1148), .B(n1147), .Y(n1149) );
  INVXL U1128 ( .A(n1164), .Y(n1159) );
  XNOR2XL U1129 ( .A(n1187), .B(n1186), .Y(n1279) );
  OAI21XL U1130 ( .A0(n1198), .A1(n1197), .B0(n1196), .Y(n1199) );
endmodule


module FFT2048_DW02_mult_2_stage_J1_14 ( A, B, TC, CLK, PRODUCT );
  input [15:0] A;
  input [26:0] B;
  output [42:0] PRODUCT;
  input TC, CLK;
  wire   n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, mult_x_1_n335, mult_x_1_n327, mult_x_1_n320,
         mult_x_1_n317, mult_x_1_n316, mult_x_1_n313, mult_x_1_n312,
         mult_x_1_n306, mult_x_1_n305, mult_x_1_n303, mult_x_1_n302,
         mult_x_1_n300, mult_x_1_n299, mult_x_1_n297, mult_x_1_n292,
         mult_x_1_n291, mult_x_1_n289, mult_x_1_n288, mult_x_1_n278,
         mult_x_1_n277, mult_x_1_n271, mult_x_1_n270, mult_x_1_n260,
         mult_x_1_n259, mult_x_1_n253, mult_x_1_n252, mult_x_1_n242,
         mult_x_1_n241, mult_x_1_n233, mult_x_1_n232, mult_x_1_n224,
         mult_x_1_n223, mult_x_1_n221, mult_x_1_n220, mult_x_1_n210,
         mult_x_1_n209, mult_x_1_n203, mult_x_1_n202, mult_x_1_n192,
         mult_x_1_n191, mult_x_1_n185, mult_x_1_n184, mult_x_1_n174,
         mult_x_1_n173, mult_x_1_n163, mult_x_1_n162, mult_x_1_n150,
         mult_x_1_n149, mult_x_1_n135, mult_x_1_n134, mult_x_1_n126,
         mult_x_1_n125, mult_x_1_n115, mult_x_1_n114, mult_x_1_n106,
         mult_x_1_n105, mult_x_1_n81, mult_x_1_n80, mult_x_1_n78, mult_x_1_n54,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290;

  DFFHQXL mult_x_1_clk_r_REG20_S1 ( .D(mult_x_1_n223), .CK(CLK), .Q(n1256) );
  DFFHQXL mult_x_1_clk_r_REG22_S1 ( .D(mult_x_1_n220), .CK(CLK), .Q(n1254) );
  DFFHQXL mult_x_1_clk_r_REG19_S1 ( .D(mult_x_1_n224), .CK(CLK), .Q(n1257) );
  DFFHQXL mult_x_1_clk_r_REG40_S1 ( .D(mult_x_1_n173), .CK(CLK), .Q(n1244) );
  DFFHQXL mult_x_1_clk_r_REG36_S1 ( .D(mult_x_1_n191), .CK(CLK), .Q(n1248) );
  DFFHQX1 mult_x_1_clk_r_REG57_S1 ( .D(mult_x_1_n320), .CK(CLK), .Q(n1288) );
  DFFHQX4 mult_x_1_clk_r_REG54_S1 ( .D(mult_x_1_n317), .CK(CLK), .Q(n1287) );
  DFFHQX4 mult_x_1_clk_r_REG55_S1 ( .D(mult_x_1_n316), .CK(CLK), .Q(n1283) );
  DFFHQX4 mult_x_1_clk_r_REG7_S1 ( .D(mult_x_1_n297), .CK(CLK), .Q(n1274) );
  DFFHQX4 mult_x_1_clk_r_REG32_S1 ( .D(mult_x_1_n288), .CK(CLK), .Q(n1270) );
  DFFHQX1 mult_x_1_clk_r_REG27_S1 ( .D(mult_x_1_n271), .CK(CLK), .Q(n1267) );
  DFFHQX4 mult_x_1_clk_r_REG16_S1 ( .D(mult_x_1_n241), .CK(CLK), .Q(n1260) );
  DFFHQX4 mult_x_1_clk_r_REG1_S1 ( .D(mult_x_1_n306), .CK(CLK), .Q(n1286) );
  DFFHQXL mult_x_1_clk_r_REG37_S1 ( .D(mult_x_1_n185), .CK(CLK), .Q(n1247) );
  DFFHQXL clk_r_REG58_S1 ( .D(n1304), .CK(CLK), .Q(PRODUCT[12]) );
  DFFHQXL clk_r_REG60_S1 ( .D(n1305), .CK(CLK), .Q(PRODUCT[11]) );
  DFFHQX4 mult_x_1_clk_r_REG31_S1 ( .D(mult_x_1_n289), .CK(CLK), .Q(n1271) );
  DFFHQXL clk_r_REG62_S1 ( .D(n1306), .CK(CLK), .Q(PRODUCT[10]) );
  DFFHQXL mult_x_1_clk_r_REG59_S1 ( .D(mult_x_1_n327), .CK(CLK), .Q(n1289) );
  DFFHQXL mult_x_1_clk_r_REG42_S1 ( .D(mult_x_1_n162), .CK(CLK), .Q(n1242) );
  DFFHQXL mult_x_1_clk_r_REG33_S1 ( .D(mult_x_1_n203), .CK(CLK), .Q(n1251) );
  DFFHQXL clk_r_REG63_S1 ( .D(n1307), .CK(CLK), .Q(PRODUCT[9]) );
  DFFHQXL mult_x_1_clk_r_REG34_S1 ( .D(mult_x_1_n202), .CK(CLK), .Q(n1250) );
  DFFHQXL mult_x_1_clk_r_REG47_S1 ( .D(mult_x_1_n126), .CK(CLK), .Q(n1237) );
  DFFHQXL mult_x_1_clk_r_REG24_S1 ( .D(mult_x_1_n209), .CK(CLK), .Q(n1252) );
  DFFHQXL mult_x_1_clk_r_REG39_S1 ( .D(mult_x_1_n174), .CK(CLK), .Q(n1245) );
  DFFHQXL mult_x_1_clk_r_REG17_S1 ( .D(mult_x_1_n233), .CK(CLK), .Q(n1259) );
  DFFHQXL clk_r_REG64_S1 ( .D(n1308), .CK(CLK), .Q(PRODUCT[8]) );
  DFFHQXL clk_r_REG65_S1 ( .D(n1309), .CK(CLK), .Q(PRODUCT[7]) );
  DFFHQXL clk_r_REG66_S1 ( .D(n1310), .CK(CLK), .Q(PRODUCT[6]) );
  DFFHQXL clk_r_REG67_S1 ( .D(n1311), .CK(CLK), .Q(PRODUCT[5]) );
  DFFHQXL clk_r_REG68_S1 ( .D(n1312), .CK(CLK), .Q(PRODUCT[4]) );
  DFFHQXL clk_r_REG69_S1 ( .D(n1313), .CK(CLK), .Q(PRODUCT[3]) );
  DFFHQXL clk_r_REG70_S1 ( .D(n1314), .CK(CLK), .Q(PRODUCT[2]) );
  DFFHQXL clk_r_REG71_S1 ( .D(n1315), .CK(CLK), .Q(PRODUCT[1]) );
  DFFHQXL clk_r_REG72_S1 ( .D(n1316), .CK(CLK), .Q(PRODUCT[0]) );
  DFFHQXL mult_x_1_clk_r_REG44_S1 ( .D(mult_x_1_n149), .CK(CLK), .Q(n1240) );
  DFFHQXL mult_x_1_clk_r_REG56_S1 ( .D(mult_x_1_n81), .CK(CLK), .Q(n1285) );
  DFFHQX1 mult_x_1_clk_r_REG53_S1 ( .D(mult_x_1_n80), .CK(CLK), .Q(n1284) );
  DFFHQXL mult_x_1_clk_r_REG0_S1 ( .D(mult_x_1_n313), .CK(CLK), .Q(n1282) );
  DFFHQX1 mult_x_1_clk_r_REG2_S1 ( .D(mult_x_1_n312), .CK(CLK), .Q(n1281) );
  DFFHQXL mult_x_1_clk_r_REG4_S1 ( .D(mult_x_1_n78), .CK(CLK), .Q(n1280) );
  DFFHQXL mult_x_1_clk_r_REG6_S1 ( .D(mult_x_1_n302), .CK(CLK), .Q(n1277) );
  DFFHQX2 mult_x_1_clk_r_REG9_S1 ( .D(mult_x_1_n299), .CK(CLK), .Q(n1275) );
  DFFHQX1 mult_x_1_clk_r_REG25_S1 ( .D(mult_x_1_n260), .CK(CLK), .Q(n1265) );
  DFFHQXL mult_x_1_clk_r_REG15_S1 ( .D(mult_x_1_n242), .CK(CLK), .Q(n1261) );
  DFFHQXL mult_x_1_clk_r_REG21_S1 ( .D(mult_x_1_n221), .CK(CLK), .Q(n1255) );
  DFFHQXL mult_x_1_clk_r_REG23_S1 ( .D(mult_x_1_n210), .CK(CLK), .Q(n1253) );
  DFFHQXL mult_x_1_clk_r_REG35_S1 ( .D(mult_x_1_n192), .CK(CLK), .Q(n1249) );
  DFFHQXL mult_x_1_clk_r_REG38_S1 ( .D(mult_x_1_n184), .CK(CLK), .Q(n1246) );
  DFFHQXL mult_x_1_clk_r_REG41_S1 ( .D(mult_x_1_n163), .CK(CLK), .Q(n1243) );
  DFFHQXL mult_x_1_clk_r_REG43_S1 ( .D(mult_x_1_n150), .CK(CLK), .Q(n1241) );
  DFFHQXL mult_x_1_clk_r_REG45_S1 ( .D(mult_x_1_n135), .CK(CLK), .Q(n1239) );
  DFFHQXL mult_x_1_clk_r_REG46_S1 ( .D(mult_x_1_n134), .CK(CLK), .Q(n1238) );
  DFFHQXL mult_x_1_clk_r_REG48_S1 ( .D(mult_x_1_n125), .CK(CLK), .Q(n1236) );
  DFFHQXL mult_x_1_clk_r_REG49_S1 ( .D(mult_x_1_n115), .CK(CLK), .Q(n1235) );
  DFFHQXL mult_x_1_clk_r_REG50_S1 ( .D(mult_x_1_n114), .CK(CLK), .Q(n1234) );
  DFFHQXL mult_x_1_clk_r_REG51_S1 ( .D(mult_x_1_n106), .CK(CLK), .Q(n1233) );
  DFFHQXL mult_x_1_clk_r_REG52_S1 ( .D(mult_x_1_n105), .CK(CLK), .Q(n1232) );
  DFFHQXL mult_x_1_clk_r_REG12_S1 ( .D(mult_x_1_n54), .CK(CLK), .Q(n1231) );
  DFFHQX2 mult_x_1_clk_r_REG8_S1 ( .D(mult_x_1_n300), .CK(CLK), .Q(n1276) );
  DFFHQX1 mult_x_1_clk_r_REG13_S1 ( .D(mult_x_1_n253), .CK(CLK), .Q(n1263) );
  DFFHQX4 mult_x_1_clk_r_REG61_S1 ( .D(mult_x_1_n335), .CK(CLK), .Q(n1290) );
  DFFHQX1 mult_x_1_clk_r_REG11_S1 ( .D(mult_x_1_n291), .CK(CLK), .Q(n1272) );
  DFFHQX2 mult_x_1_clk_r_REG3_S1 ( .D(mult_x_1_n305), .CK(CLK), .Q(n1279) );
  DFFHQX2 mult_x_1_clk_r_REG5_S1 ( .D(mult_x_1_n303), .CK(CLK), .Q(n1278) );
  DFFHQX1 mult_x_1_clk_r_REG30_S1 ( .D(mult_x_1_n277), .CK(CLK), .Q(n1268) );
  DFFHQX2 mult_x_1_clk_r_REG29_S1 ( .D(mult_x_1_n278), .CK(CLK), .Q(n1269) );
  DFFHQX2 mult_x_1_clk_r_REG28_S1 ( .D(mult_x_1_n270), .CK(CLK), .Q(n1266) );
  DFFHQX2 mult_x_1_clk_r_REG10_S1 ( .D(mult_x_1_n292), .CK(CLK), .Q(n1273) );
  DFFHQX1 mult_x_1_clk_r_REG18_S1 ( .D(mult_x_1_n232), .CK(CLK), .Q(n1258) );
  DFFHQX1 mult_x_1_clk_r_REG26_S1 ( .D(mult_x_1_n259), .CK(CLK), .Q(n1264) );
  DFFHQX2 mult_x_1_clk_r_REG14_S1 ( .D(mult_x_1_n252), .CK(CLK), .Q(n1262) );
  XOR2X1 U1 ( .A(n56), .B(n880), .Y(n899) );
  ADDFHX1 U2 ( .A(n647), .B(n646), .CI(n645), .CO(n641), .S(n673) );
  ADDFHX1 U3 ( .A(n763), .B(n762), .CI(n761), .CO(n754), .S(n796) );
  OAI2BB1X1 U4 ( .A0N(n81), .A1N(n792), .B0(n80), .Y(n762) );
  ADDFHX1 U5 ( .A(n607), .B(n606), .CI(n605), .CO(n581), .S(n613) );
  ADDFHX1 U6 ( .A(n640), .B(n639), .CI(n638), .CO(n614), .S(n645) );
  ADDFHX1 U7 ( .A(n495), .B(n494), .CI(n493), .CO(n497), .S(n507) );
  ADDFHX2 U8 ( .A(n671), .B(n670), .CI(n669), .CO(n646), .S(n686) );
  ADDFHX1 U9 ( .A(n628), .B(n627), .CI(n626), .CO(n640), .S(n670) );
  ADDFX2 U10 ( .A(n780), .B(n779), .CI(n778), .CO(n794), .S(n836) );
  CMPR32X1 U11 ( .A(n634), .B(n633), .C(n632), .CO(n626), .S(n690) );
  ADDFX2 U12 ( .A(n659), .B(n658), .CI(n657), .CO(n671), .S(n713) );
  ADDFHX1 U13 ( .A(n970), .B(n969), .CI(n968), .CO(n991), .S(n993) );
  NAND2X1 U14 ( .A(n16), .B(n99), .Y(n15) );
  ADDFX2 U15 ( .A(n747), .B(n746), .CI(n745), .CO(n737), .S(n805) );
  ADDFHX1 U16 ( .A(n1035), .B(n1034), .CI(n1033), .CO(n1043), .S(n386) );
  ADDFX2 U17 ( .A(n373), .B(n372), .CI(n371), .CO(n377), .S(n379) );
  XNOR2X2 U18 ( .A(B[10]), .B(n518), .Y(n351) );
  BUFX3 U19 ( .A(A[3]), .Y(n469) );
  BUFX3 U20 ( .A(A[1]), .Y(n518) );
  XNOR2X2 U21 ( .A(n612), .B(n611), .Y(PRODUCT[28]) );
  NAND2BX1 U22 ( .AN(n210), .B(n79), .Y(n501) );
  XNOR2X1 U23 ( .A(n760), .B(n759), .Y(PRODUCT[24]) );
  XOR2X2 U24 ( .A(n51), .B(n901), .Y(PRODUCT[20]) );
  XOR2X1 U25 ( .A(n937), .B(n1280), .Y(PRODUCT[16]) );
  XNOR2XL U26 ( .A(n438), .B(n437), .Y(PRODUCT[33]) );
  INVX1 U27 ( .A(n518), .Y(n8) );
  XOR2XL U28 ( .A(B[9]), .B(n8), .Y(n352) );
  XNOR2XL U29 ( .A(n1128), .B(n1127), .Y(PRODUCT[38]) );
  XNOR2XL U30 ( .A(n1091), .B(B[14]), .Y(n630) );
  XNOR2XL U31 ( .A(B[14]), .B(n469), .Y(n169) );
  XNOR2XL U32 ( .A(A[5]), .B(B[13]), .Y(n241) );
  XNOR2XL U33 ( .A(A[15]), .B(n781), .Y(n468) );
  XNOR2XL U34 ( .A(B[17]), .B(n1091), .Y(n75) );
  XNOR2XL U35 ( .A(A[2]), .B(n518), .Y(n556) );
  XNOR2XL U36 ( .A(A[10]), .B(A[9]), .Y(n1138) );
  OAI21XL U37 ( .A0(n19), .A1(n20), .B0(n18), .Y(n385) );
  XOR2XL U38 ( .A(n909), .B(n910), .Y(n34) );
  ADDFX2 U39 ( .A(n595), .B(n594), .CI(n593), .CO(n607), .S(n639) );
  XOR2XL U40 ( .A(n994), .B(n995), .Y(n112) );
  ADDFX2 U41 ( .A(n1085), .B(n1084), .CI(n1083), .CO(n1101), .S(n430) );
  XNOR2XL U42 ( .A(n1198), .B(n1197), .Y(n1310) );
  AND2X1 U43 ( .A(n800), .B(n1265), .Y(n5) );
  NOR2X1 U44 ( .A(n755), .B(n754), .Y(mult_x_1_n241) );
  XNOR2X1 U45 ( .A(n1076), .B(n1075), .Y(n1307) );
  NAND2XL U46 ( .A(n68), .B(n686), .Y(n67) );
  XOR2X1 U47 ( .A(n1188), .B(n1187), .Y(n1308) );
  NAND2X1 U48 ( .A(n997), .B(n996), .Y(mult_x_1_n313) );
  NOR2X1 U49 ( .A(n1049), .B(n1048), .Y(n1050) );
  INVX1 U50 ( .A(n1045), .Y(n30) );
  ADDFHX2 U51 ( .A(n533), .B(n532), .CI(n531), .CO(n508), .S(n544) );
  NOR2X1 U52 ( .A(n1044), .B(n1043), .Y(n1036) );
  NAND2X1 U53 ( .A(n384), .B(n383), .Y(n1068) );
  NAND2X1 U54 ( .A(n377), .B(n378), .Y(n18) );
  NOR2X1 U55 ( .A(n377), .B(n378), .Y(n19) );
  INVX1 U56 ( .A(n738), .Y(n62) );
  XNOR2X1 U57 ( .A(n553), .B(n552), .Y(n594) );
  XNOR2X1 U58 ( .A(n774), .B(B[24]), .Y(n407) );
  OAI22XL U59 ( .A0(n1161), .A1(n515), .B0(n1162), .B1(n513), .Y(n560) );
  OAI22X1 U60 ( .A0(n562), .A1(n1137), .B0(n75), .B1(n1110), .Y(n568) );
  INVX1 U61 ( .A(n378), .Y(n21) );
  XNOR2X1 U62 ( .A(n518), .B(n1174), .Y(n550) );
  ADDFHX1 U63 ( .A(n370), .B(n369), .CI(n368), .CO(n1025), .S(n378) );
  XNOR2X1 U64 ( .A(n1226), .B(n1231), .Y(PRODUCT[40]) );
  BUFX1 U65 ( .A(n1078), .Y(n1216) );
  INVX1 U66 ( .A(n501), .Y(n502) );
  CLKINVX3 U67 ( .A(n8), .Y(n769) );
  CLKINVX3 U68 ( .A(n399), .Y(n782) );
  INVXL U69 ( .A(n774), .Y(n7) );
  INVX1 U70 ( .A(n503), .Y(n6) );
  NAND2X1 U71 ( .A(n758), .B(n1263), .Y(n759) );
  INVX1 U72 ( .A(n841), .Y(n876) );
  INVX1 U73 ( .A(n1287), .Y(n12) );
  INVX1 U74 ( .A(n1248), .Y(n504) );
  NOR2X1 U75 ( .A(n1256), .B(n1254), .Y(n536) );
  AOI21X1 U76 ( .A0(n1056), .A1(n1060), .B0(n1047), .Y(n1053) );
  XNOR2X1 U77 ( .A(n1070), .B(n1069), .Y(n1306) );
  NAND2BX1 U78 ( .AN(n1046), .B(n30), .Y(n1056) );
  NAND2X1 U79 ( .A(n1049), .B(n1048), .Y(n1051) );
  OAI21X1 U80 ( .A0(n244), .A1(n245), .B0(n15), .Y(n13) );
  ADDFHX1 U81 ( .A(n509), .B(n508), .CI(n507), .CO(n500), .S(n535) );
  NOR2X1 U82 ( .A(n997), .B(n996), .Y(mult_x_1_n312) );
  NAND2XL U83 ( .A(n111), .B(n993), .Y(n110) );
  NAND2X1 U84 ( .A(n386), .B(n385), .Y(n1064) );
  NAND2X1 U85 ( .A(n1044), .B(n1043), .Y(n1057) );
  ADDFHX1 U86 ( .A(n1042), .B(n1041), .CI(n1040), .CO(n1048), .S(n1046) );
  NAND2BXL U87 ( .AN(n909), .B(n115), .Y(n114) );
  INVX1 U88 ( .A(n385), .Y(n24) );
  INVX1 U89 ( .A(n244), .Y(n14) );
  NAND2XL U90 ( .A(n1028), .B(n1029), .Y(n27) );
  NAND2X1 U91 ( .A(n23), .B(n22), .Y(n1034) );
  NAND2BXL U92 ( .AN(n1028), .B(n29), .Y(n28) );
  OR2X2 U93 ( .A(n384), .B(n383), .Y(n382) );
  INVXL U94 ( .A(n336), .Y(n95) );
  INVXL U95 ( .A(n1029), .Y(n29) );
  NAND2X1 U96 ( .A(n342), .B(n341), .Y(n1185) );
  OR2XL U97 ( .A(n553), .B(n552), .Y(n559) );
  NOR2X1 U98 ( .A(n342), .B(n341), .Y(n1184) );
  OAI22XL U99 ( .A0(n1141), .A1(n818), .B0(n1162), .B1(n777), .Y(n829) );
  NAND2X1 U100 ( .A(n675), .B(n206), .Y(n207) );
  NAND2X1 U101 ( .A(n643), .B(n1257), .Y(n644) );
  NAND2X1 U102 ( .A(n53), .B(n1273), .Y(n916) );
  INVX1 U103 ( .A(n46), .Y(n11) );
  NAND2X1 U104 ( .A(n926), .B(n1276), .Y(n927) );
  NAND2X1 U105 ( .A(n211), .B(n536), .Y(n503) );
  NAND2X1 U106 ( .A(n504), .B(n1249), .Y(n505) );
  NAND2X1 U107 ( .A(n541), .B(n1251), .Y(n542) );
  NAND2X1 U108 ( .A(n577), .B(n1253), .Y(n578) );
  NAND2X1 U109 ( .A(n465), .B(n1247), .Y(n466) );
  NAND2X1 U110 ( .A(n436), .B(n1245), .Y(n437) );
  INVX1 U111 ( .A(n1240), .Y(n232) );
  INVX1 U112 ( .A(n1242), .Y(n395) );
  INVX1 U113 ( .A(n1236), .Y(n1120) );
  INVX1 U114 ( .A(n1273), .Y(n52) );
  BUFX3 U115 ( .A(A[13]), .Y(n1129) );
  INVXL U116 ( .A(A[5]), .Y(n399) );
  NOR2X1 U117 ( .A(n1248), .B(n1246), .Y(n223) );
  NOR2X1 U118 ( .A(n930), .B(n929), .Y(mult_x_1_n299) );
  NAND2XL U119 ( .A(n899), .B(n898), .Y(mult_x_1_n278) );
  OAI2BB1X2 U120 ( .A0N(n244), .A1N(n245), .B0(n13), .Y(n922) );
  NAND2X1 U121 ( .A(n25), .B(n24), .Y(n1065) );
  NAND2XL U122 ( .A(n881), .B(n882), .Y(n89) );
  XNOR3X2 U123 ( .A(n245), .B(n14), .C(n15), .Y(n258) );
  NAND2XL U124 ( .A(n903), .B(n904), .Y(n116) );
  NAND2XL U125 ( .A(n105), .B(n850), .Y(n106) );
  INVX1 U126 ( .A(n386), .Y(n25) );
  NAND2XL U127 ( .A(n724), .B(n725), .Y(n35) );
  NAND2BXL U128 ( .AN(n724), .B(n37), .Y(n36) );
  INVXL U129 ( .A(n571), .Y(n58) );
  NAND2XL U130 ( .A(n571), .B(n572), .Y(n124) );
  NAND2XL U131 ( .A(n687), .B(n688), .Y(n66) );
  NAND2XL U132 ( .A(n994), .B(n995), .Y(n109) );
  NOR2X1 U133 ( .A(n1072), .B(n1184), .Y(n346) );
  OAI2BB1X1 U134 ( .A0N(n28), .A1N(n1027), .B0(n27), .Y(n1041) );
  INVXL U135 ( .A(n725), .Y(n37) );
  ADDFHX2 U136 ( .A(n753), .B(n752), .CI(n751), .CO(n724), .S(n761) );
  OR2XL U137 ( .A(n1181), .B(n1180), .Y(n1183) );
  NAND2XL U138 ( .A(n794), .B(n793), .Y(n80) );
  INVXL U139 ( .A(n793), .Y(n82) );
  INVXL U140 ( .A(n904), .Y(n119) );
  INVXL U141 ( .A(n910), .Y(n115) );
  XOR3X2 U142 ( .A(n1029), .B(n1028), .C(n1027), .Y(n1030) );
  ADDFHX2 U143 ( .A(n204), .B(n203), .CI(n202), .CO(n259), .S(n990) );
  ADDFHX2 U144 ( .A(n837), .B(n836), .CI(n835), .CO(n802), .S(n848) );
  NOR2X1 U145 ( .A(n344), .B(n343), .Y(n1072) );
  ADDFHX1 U146 ( .A(n527), .B(n526), .CI(n525), .CO(n520), .S(n584) );
  ADDFHX1 U147 ( .A(n861), .B(n860), .CI(n859), .CO(n873), .S(n896) );
  ADDFHX1 U148 ( .A(n569), .B(n568), .CI(n567), .CO(n585), .S(n616) );
  OAI2BB1XL U149 ( .A0N(n1077), .A1N(n953), .B0(n519), .Y(n564) );
  XOR3X2 U150 ( .A(n21), .B(n377), .C(n20), .Y(n384) );
  NAND2X1 U151 ( .A(n375), .B(n376), .Y(n22) );
  OAI22X1 U152 ( .A0(n963), .A1(n523), .B0(n961), .B1(n470), .Y(n488) );
  ADDFHX1 U153 ( .A(n831), .B(n830), .CI(n829), .CO(n820), .S(n884) );
  ADDFHX1 U154 ( .A(n867), .B(n866), .CI(n865), .CO(n859), .S(n906) );
  INVXL U155 ( .A(n87), .Y(n86) );
  XNOR3X2 U156 ( .A(n376), .B(n375), .C(n374), .Y(n20) );
  NAND2XL U157 ( .A(n73), .B(n70), .Y(n69) );
  OAI22X1 U158 ( .A0(n953), .A1(n26), .B0(n952), .B1(n1077), .Y(n985) );
  NAND2XL U159 ( .A(n73), .B(n72), .Y(n71) );
  OAI22X1 U160 ( .A0(n563), .A1(n959), .B0(n514), .B1(n957), .Y(n553) );
  OAI22X1 U161 ( .A0(n1077), .A1(n352), .B0(n266), .B1(n953), .Y(n350) );
  NAND2BXL U162 ( .AN(n775), .B(n40), .Y(n39) );
  INVXL U163 ( .A(n94), .Y(n93) );
  OR2X2 U164 ( .A(n315), .B(n314), .Y(n313) );
  XNOR2X1 U165 ( .A(n1168), .B(n1167), .Y(PRODUCT[39]) );
  AND2XL U166 ( .A(n1214), .B(n1213), .Y(n1315) );
  OR2XL U167 ( .A(n1212), .B(n1211), .Y(n1214) );
  OAI22XL U168 ( .A0(n1112), .A1(n955), .B0(n1110), .B1(n954), .Y(n984) );
  XOR2X2 U169 ( .A(n54), .B(n5), .Y(PRODUCT[23]) );
  NAND2BXL U170 ( .AN(n218), .B(n501), .Y(n78) );
  BUFX4 U171 ( .A(n674), .Y(n41) );
  INVXL U172 ( .A(n963), .Y(n70) );
  INVXL U173 ( .A(n798), .Y(n799) );
  AND2XL U174 ( .A(n1215), .B(n1218), .Y(n1222) );
  INVXL U175 ( .A(n1089), .Y(n40) );
  INVXL U176 ( .A(n961), .Y(n72) );
  NOR2BXL U177 ( .AN(B[0]), .B(n1162), .Y(n986) );
  NAND2X1 U178 ( .A(n900), .B(n1271), .Y(n901) );
  AND2X2 U179 ( .A(n878), .B(n1269), .Y(n879) );
  NAND2X1 U180 ( .A(n126), .B(n127), .Y(n347) );
  NAND2X1 U181 ( .A(n131), .B(n132), .Y(n697) );
  INVX1 U182 ( .A(n1129), .Y(n159) );
  INVXL U183 ( .A(n1091), .Y(n77) );
  INVX1 U184 ( .A(n1238), .Y(n1118) );
  XNOR2X1 U185 ( .A(A[8]), .B(A[7]), .Y(n132) );
  INVXL U186 ( .A(n942), .Y(n9) );
  INVX1 U187 ( .A(A[0]), .Y(n140) );
  INVX1 U188 ( .A(n1268), .Y(n878) );
  INVXL U189 ( .A(n1246), .Y(n465) );
  NOR2BX1 U190 ( .AN(n1267), .B(n97), .Y(n96) );
  NAND2BX1 U191 ( .AN(n207), .B(n798), .Y(n123) );
  OAI22X1 U192 ( .A0(n697), .A1(n733), .B0(n1090), .B1(n696), .Y(n747) );
  XNOR2X2 U193 ( .A(n722), .B(n721), .Y(PRODUCT[25]) );
  CLKINVX3 U194 ( .A(n41), .Y(n917) );
  ADDFX2 U195 ( .A(n897), .B(n896), .CI(n895), .CO(n881), .S(n902) );
  XNOR2X1 U196 ( .A(n774), .B(B[10]), .Y(n815) );
  OAI22X2 U197 ( .A0(n963), .A1(n960), .B0(n961), .B1(n197), .Y(n978) );
  NOR2X1 U198 ( .A(n999), .B(n998), .Y(n1000) );
  OAI21XL U199 ( .A0(n1072), .A1(n1185), .B0(n1073), .Y(n345) );
  XOR2X1 U200 ( .A(n1067), .B(n1066), .Y(n1305) );
  XNOR2X1 U201 ( .A(B[19]), .B(n469), .Y(n734) );
  NAND2X2 U202 ( .A(n10), .B(n42), .Y(n674) );
  NAND2X1 U203 ( .A(n1005), .B(n11), .Y(n10) );
  OAI2BB1X2 U204 ( .A0N(n1283), .A1N(n1290), .B0(n12), .Y(n1005) );
  NOR2X1 U205 ( .A(mult_x_1_n299), .B(mult_x_1_n302), .Y(mult_x_1_n297) );
  NOR2X1 U206 ( .A(n186), .B(n185), .Y(n17) );
  NAND2BX1 U207 ( .AN(n17), .B(n184), .Y(n16) );
  XOR2X1 U208 ( .A(B[8]), .B(n7), .Y(n167) );
  OAI21XL U209 ( .A0(n375), .A1(n376), .B0(n374), .Y(n23) );
  OAI22X1 U210 ( .A0(n351), .A1(n953), .B0(n1077), .B1(n26), .Y(n983) );
  XNOR2X1 U211 ( .A(n773), .B(n518), .Y(n26) );
  BUFX3 U212 ( .A(n33), .Y(n31) );
  AOI21X4 U213 ( .A0(n209), .A1(n41), .B0(n208), .Y(n33) );
  OAI21XL U214 ( .A0(n33), .A1(n576), .B0(n575), .Y(n579) );
  OAI21X1 U215 ( .A0(n33), .A1(n1256), .B0(n1257), .Y(n612) );
  OAI21XL U216 ( .A0(n33), .A1(n540), .B0(n539), .Y(n543) );
  XOR2X2 U217 ( .A(n33), .B(n644), .Y(PRODUCT[27]) );
  OAI2BB1X1 U218 ( .A0N(n6), .A1N(n32), .B0(n502), .Y(n506) );
  INVX1 U219 ( .A(n33), .Y(n32) );
  OAI21XL U220 ( .A0(n33), .A1(n464), .B0(n463), .Y(n467) );
  OAI21XL U221 ( .A0(n31), .A1(n231), .B0(n230), .Y(n234) );
  OAI21XL U222 ( .A0(n31), .A1(n394), .B0(n393), .Y(n397) );
  OAI21XL U223 ( .A0(n33), .A1(n435), .B0(n434), .Y(n438) );
  OAI21XL U224 ( .A0(n31), .A1(n220), .B0(n219), .Y(n222) );
  OAI21XL U225 ( .A0(n31), .A1(n1080), .B0(n1079), .Y(n1082) );
  OAI21XL U226 ( .A0(n31), .A1(n1125), .B0(n1124), .Y(n1128) );
  OAI21XL U227 ( .A0(n31), .A1(n1166), .B0(n1165), .Y(n1168) );
  OAI21XL U228 ( .A0(n31), .A1(n1225), .B0(n1224), .Y(n1226) );
  NAND2XL U229 ( .A(n930), .B(n929), .Y(mult_x_1_n300) );
  XOR2X1 U230 ( .A(n908), .B(n34), .Y(n921) );
  XNOR2X1 U231 ( .A(B[17]), .B(n769), .Y(n249) );
  OAI2BB1X1 U232 ( .A0N(n36), .A1N(n723), .B0(n35), .Y(n715) );
  XOR2X1 U233 ( .A(n723), .B(n38), .Y(n755) );
  XOR2X1 U234 ( .A(n724), .B(n725), .Y(n38) );
  OAI21XL U235 ( .A0(n1090), .A1(n733), .B0(n39), .Y(n788) );
  XNOR2X1 U236 ( .A(B[13]), .B(n774), .Y(n733) );
  XNOR2X1 U237 ( .A(B[18]), .B(n782), .Y(n703) );
  NAND3X1 U238 ( .A(n674), .B(n797), .C(n800), .Y(n45) );
  INVX1 U239 ( .A(n677), .Y(n797) );
  NAND2X1 U240 ( .A(n840), .B(n205), .Y(n677) );
  NOR2X2 U241 ( .A(n44), .B(n43), .Y(n42) );
  INVX1 U242 ( .A(n50), .Y(n43) );
  OAI21X2 U243 ( .A0(n1275), .A1(n1278), .B0(n1276), .Y(n44) );
  NAND2X1 U244 ( .A(n757), .B(n45), .Y(n760) );
  XOR2X2 U245 ( .A(n916), .B(n917), .Y(PRODUCT[19]) );
  NAND2X1 U246 ( .A(n1279), .B(n1274), .Y(n46) );
  XOR2X2 U247 ( .A(n47), .B(n879), .Y(PRODUCT[21]) );
  NAND2X1 U248 ( .A(n48), .B(n876), .Y(n47) );
  NAND2BX1 U249 ( .AN(n877), .B(n41), .Y(n48) );
  NAND2X1 U250 ( .A(n49), .B(n843), .Y(n847) );
  NAND2BX1 U251 ( .AN(n844), .B(n41), .Y(n49) );
  NAND2X1 U252 ( .A(n1286), .B(n1274), .Y(n50) );
  NOR2X1 U253 ( .A(n1268), .B(n1266), .Y(n205) );
  NOR2X1 U254 ( .A(n1272), .B(n1270), .Y(n840) );
  AOI21X1 U255 ( .A0(n41), .A1(n53), .B0(n52), .Y(n51) );
  INVX1 U256 ( .A(n1272), .Y(n53) );
  NAND2X1 U257 ( .A(n799), .B(n55), .Y(n54) );
  NAND2BXL U258 ( .AN(n677), .B(n674), .Y(n55) );
  NOR2X1 U259 ( .A(n1264), .B(n1262), .Y(n675) );
  XOR2X1 U260 ( .A(n881), .B(n882), .Y(n56) );
  OAI22X1 U261 ( .A0(n963), .A1(n172), .B0(n169), .B1(n961), .Y(n179) );
  XNOR2X1 U262 ( .A(B[13]), .B(n469), .Y(n172) );
  XNOR2X1 U263 ( .A(B[20]), .B(n769), .Y(n770) );
  OAI2BB1X1 U264 ( .A0N(n57), .A1N(n570), .B0(n124), .Y(n545) );
  NAND2BXL U265 ( .AN(n572), .B(n58), .Y(n57) );
  XOR2X1 U266 ( .A(B[21]), .B(n9), .Y(n514) );
  XNOR2X1 U267 ( .A(B[20]), .B(n942), .Y(n563) );
  XNOR2X1 U268 ( .A(n774), .B(B[17]), .Y(n591) );
  AOI2BB1X2 U269 ( .A0N(n239), .A1N(n961), .B0(n104), .Y(n103) );
  OAI21XL U270 ( .A0(n103), .A1(n102), .B0(n100), .Y(n886) );
  OAI22X1 U271 ( .A0(n967), .A1(n824), .B0(n965), .B1(n823), .Y(n870) );
  OAI22X1 U272 ( .A0(n953), .A1(n809), .B0(n770), .B1(n1077), .Y(n808) );
  NAND2XL U273 ( .A(n1118), .B(n1239), .Y(n221) );
  INVXL U274 ( .A(n1078), .Y(n220) );
  XNOR2XL U275 ( .A(n774), .B(n740), .Y(n623) );
  XNOR2XL U276 ( .A(n469), .B(B[22]), .Y(n624) );
  ADDFX2 U277 ( .A(n299), .B(n59), .CI(n297), .CO(n336), .S(n335) );
  OAI22XL U278 ( .A0(n963), .A1(n300), .B0(n961), .B1(n291), .Y(n299) );
  AOI21XL U279 ( .A0(n501), .A1(n392), .B0(n391), .Y(n393) );
  AOI21XL U280 ( .A0(n798), .A1(n800), .B0(n756), .Y(n757) );
  INVXL U281 ( .A(n1265), .Y(n756) );
  XNOR2X1 U282 ( .A(n234), .B(n233), .Y(PRODUCT[35]) );
  NAND2XL U283 ( .A(n232), .B(n1241), .Y(n233) );
  XNOR2X2 U284 ( .A(n579), .B(n578), .Y(PRODUCT[29]) );
  INVXL U285 ( .A(n1256), .Y(n643) );
  XNOR2X1 U286 ( .A(n685), .B(n684), .Y(PRODUCT[26]) );
  NAND2XL U287 ( .A(n683), .B(n1259), .Y(n684) );
  OAI21XL U288 ( .A0(n917), .A1(n682), .B0(n681), .Y(n685) );
  INVXL U289 ( .A(n1258), .Y(n683) );
  NAND2XL U290 ( .A(n676), .B(n1261), .Y(n721) );
  OAI21XL U291 ( .A0(n917), .A1(n720), .B0(n719), .Y(n722) );
  INVXL U292 ( .A(n1260), .Y(n676) );
  XNOR2XL U293 ( .A(n1129), .B(B[12]), .Y(n625) );
  XNOR2XL U294 ( .A(n1091), .B(B[8]), .Y(n826) );
  XNOR2XL U295 ( .A(n942), .B(B[12]), .Y(n828) );
  XNOR2XL U296 ( .A(n774), .B(B[9]), .Y(n238) );
  XNOR2XL U297 ( .A(n1091), .B(B[7]), .Y(n242) );
  XNOR2XL U298 ( .A(n942), .B(n773), .Y(n243) );
  XNOR2XL U299 ( .A(n942), .B(n1174), .Y(n403) );
  XNOR2XL U300 ( .A(B[25]), .B(n774), .Y(n419) );
  XNOR2XL U301 ( .A(n1129), .B(B[20]), .Y(n405) );
  XNOR2XL U302 ( .A(B[25]), .B(n942), .Y(n408) );
  XNOR2XL U303 ( .A(n1129), .B(B[18]), .Y(n443) );
  XNOR2X1 U304 ( .A(B[25]), .B(n469), .Y(n523) );
  XNOR2XL U305 ( .A(n942), .B(B[18]), .Y(n631) );
  NAND2XL U306 ( .A(n1126), .B(n1235), .Y(n1127) );
  INVXL U307 ( .A(n1234), .Y(n1126) );
  OAI22XL U308 ( .A0(n1141), .A1(n699), .B0(n1162), .B1(n656), .Y(n706) );
  OAI22XL U309 ( .A0(n1141), .A1(n736), .B0(n1162), .B1(n699), .Y(n745) );
  XNOR2XL U310 ( .A(n942), .B(B[8]), .Y(n177) );
  XNOR2XL U311 ( .A(n469), .B(B[12]), .Y(n173) );
  XNOR2XL U312 ( .A(n1091), .B(B[4]), .Y(n175) );
  XOR2XL U313 ( .A(B[18]), .B(n77), .Y(n76) );
  XNOR2XL U314 ( .A(n774), .B(B[21]), .Y(n481) );
  XNOR2XL U315 ( .A(n1129), .B(B[22]), .Y(n1093) );
  XNOR2XL U316 ( .A(B[25]), .B(n1091), .Y(n1111) );
  XNOR2XL U317 ( .A(n1129), .B(B[23]), .Y(n1108) );
  XNOR2XL U318 ( .A(n1091), .B(B[23]), .Y(n420) );
  XNOR2XL U319 ( .A(n774), .B(n1174), .Y(n1087) );
  XNOR2XL U320 ( .A(n774), .B(B[22]), .Y(n444) );
  XNOR2XL U321 ( .A(n1091), .B(B[22]), .Y(n406) );
  NAND2XL U322 ( .A(n1218), .B(n1233), .Y(n1167) );
  XNOR2XL U323 ( .A(n1129), .B(n1174), .Y(n1159) );
  XNOR2XL U324 ( .A(B[25]), .B(A[15]), .Y(n1177) );
  XNOR2XL U325 ( .A(B[25]), .B(n1129), .Y(n1140) );
  XNOR2XL U326 ( .A(n1129), .B(B[24]), .Y(n1130) );
  ADDFX2 U327 ( .A(n248), .B(n247), .CI(n246), .CO(n910), .S(n244) );
  OAI21XL U328 ( .A0(n340), .A1(n1189), .B0(n339), .Y(n1071) );
  NAND2XL U329 ( .A(n1192), .B(n1196), .Y(n340) );
  AOI21XL U330 ( .A0(n1192), .A1(n1190), .B0(n338), .Y(n339) );
  NAND2XL U331 ( .A(n1212), .B(n1211), .Y(n1213) );
  INVXL U332 ( .A(n1163), .Y(n1123) );
  INVXL U333 ( .A(n1239), .Y(n1121) );
  NAND2XL U334 ( .A(n1216), .B(n1118), .Y(n1080) );
  AOI21XL U335 ( .A0(n501), .A1(n229), .B0(n228), .Y(n230) );
  INVXL U336 ( .A(n1245), .Y(n225) );
  AOI21XL U337 ( .A0(n501), .A1(n504), .B0(n462), .Y(n463) );
  INVXL U338 ( .A(n1249), .Y(n462) );
  INVXL U339 ( .A(n1253), .Y(n538) );
  INVXL U340 ( .A(n1252), .Y(n577) );
  XNOR2X1 U341 ( .A(n942), .B(n771), .Y(n958) );
  XNOR2XL U342 ( .A(n469), .B(B[9]), .Y(n962) );
  XNOR2XL U343 ( .A(n1091), .B(B[1]), .Y(n955) );
  XNOR2XL U344 ( .A(n1091), .B(B[0]), .Y(n366) );
  NAND2BXL U345 ( .AN(B[0]), .B(n774), .Y(n265) );
  NAND2X1 U346 ( .A(n841), .B(n205), .Y(n98) );
  NAND2XL U347 ( .A(n395), .B(n1243), .Y(n396) );
  XNOR2XL U348 ( .A(n469), .B(B[21]), .Y(n655) );
  XNOR2XL U349 ( .A(n1129), .B(n773), .Y(n656) );
  XNOR2X1 U350 ( .A(n782), .B(B[19]), .Y(n660) );
  XNOR2XL U351 ( .A(n1091), .B(B[13]), .Y(n661) );
  XNOR2XL U352 ( .A(n942), .B(B[17]), .Y(n662) );
  XNOR2XL U353 ( .A(n942), .B(B[14]), .Y(n785) );
  XNOR2XL U354 ( .A(n942), .B(B[13]), .Y(n827) );
  XNOR2XL U355 ( .A(n1129), .B(B[7]), .Y(n818) );
  XNOR2XL U356 ( .A(n469), .B(n740), .Y(n817) );
  XNOR2XL U357 ( .A(n1129), .B(n941), .Y(n819) );
  XNOR2X1 U358 ( .A(n1129), .B(n771), .Y(n240) );
  INVXL U359 ( .A(A[15]), .Y(n144) );
  XNOR2XL U360 ( .A(n942), .B(B[7]), .Y(n943) );
  XNOR2XL U361 ( .A(n942), .B(n941), .Y(n956) );
  XNOR2XL U362 ( .A(n1091), .B(B[3]), .Y(n946) );
  XNOR2X1 U363 ( .A(n774), .B(n771), .Y(n196) );
  NAND2BXL U364 ( .AN(B[0]), .B(n1129), .Y(n158) );
  XNOR2XL U365 ( .A(n774), .B(B[3]), .Y(n981) );
  NAND2BXL U366 ( .AN(B[0]), .B(n1091), .Y(n348) );
  XNOR2XL U367 ( .A(n942), .B(B[3]), .Y(n361) );
  XNOR2XL U368 ( .A(n942), .B(B[4]), .Y(n365) );
  XNOR2XL U369 ( .A(n469), .B(B[8]), .Y(n367) );
  XNOR2XL U370 ( .A(n469), .B(B[7]), .Y(n364) );
  XNOR2X1 U371 ( .A(n1129), .B(B[19]), .Y(n409) );
  OAI22X1 U372 ( .A0(n652), .A1(n953), .B0(n621), .B1(n1077), .Y(n74) );
  NAND2BXL U373 ( .AN(B[0]), .B(n942), .Y(n263) );
  NOR2XL U374 ( .A(n1163), .B(n1234), .Y(n1215) );
  INVXL U375 ( .A(n1232), .Y(n1218) );
  OAI22XL U376 ( .A0(n1141), .A1(n625), .B0(n1162), .B1(n592), .Y(n632) );
  OAI21X1 U377 ( .A0(n624), .A1(n963), .B0(n71), .Y(n633) );
  CMPR32X1 U378 ( .A(n711), .B(n710), .C(n709), .CO(n728), .S(n764) );
  OAI22XL U379 ( .A0(n744), .A1(n705), .B0(n957), .B1(n662), .Y(n709) );
  OAI22XL U380 ( .A0(n1112), .A1(n704), .B0(n1110), .B1(n661), .Y(n710) );
  OAI22XL U381 ( .A0(n967), .A1(n703), .B0(n965), .B1(n660), .Y(n711) );
  OAI22XL U382 ( .A0(n1141), .A1(n777), .B0(n1162), .B1(n736), .Y(n786) );
  CMPR32X1 U383 ( .A(n791), .B(n790), .C(n789), .CO(n806), .S(n851) );
  OAI22XL U384 ( .A0(n744), .A1(n785), .B0(n957), .B1(n743), .Y(n789) );
  OAI22XL U385 ( .A0(n1112), .A1(n784), .B0(n1110), .B1(n742), .Y(n790) );
  OAI22XL U386 ( .A0(n967), .A1(n783), .B0(n965), .B1(n741), .Y(n791) );
  OAI22XL U387 ( .A0(n959), .A1(n243), .B0(n957), .B1(n828), .Y(n862) );
  OAI22XL U388 ( .A0(n1112), .A1(n242), .B0(n1110), .B1(n826), .Y(n863) );
  OAI22XL U389 ( .A0(n1141), .A1(n151), .B0(n1162), .B1(n171), .Y(n153) );
  OAI22XL U390 ( .A0(n1178), .A1(n150), .B0(n1176), .B1(n149), .Y(n154) );
  XNOR2XL U391 ( .A(n774), .B(B[20]), .Y(n486) );
  XNOR2X1 U392 ( .A(n1091), .B(B[19]), .Y(n482) );
  XNOR2XL U393 ( .A(n1091), .B(B[24]), .Y(n1092) );
  XNOR2XL U394 ( .A(n774), .B(B[23]), .Y(n439) );
  OAI22XL U395 ( .A0(n1089), .A1(n481), .B0(n1090), .B1(n444), .Y(n472) );
  XNOR2XL U396 ( .A(n1091), .B(B[21]), .Y(n410) );
  OAI2BB1XL U397 ( .A0N(n965), .A1N(n967), .B0(n401), .Y(n448) );
  OAI22XL U398 ( .A0(n1178), .A1(n442), .B0(n1176), .B1(n398), .Y(n450) );
  INVXL U399 ( .A(n400), .Y(n401) );
  OAI2BB1XL U400 ( .A0N(n957), .A1N(n744), .B0(n404), .Y(n421) );
  OAI22XL U401 ( .A0(n1178), .A1(n402), .B0(n1176), .B1(n418), .Y(n423) );
  INVXL U402 ( .A(n403), .Y(n404) );
  OAI22XL U403 ( .A0(n1141), .A1(n405), .B0(n1162), .B1(n417), .Y(n426) );
  OAI22XL U404 ( .A0(n1089), .A1(n407), .B0(n1090), .B1(n419), .Y(n424) );
  OAI22X1 U405 ( .A0(n76), .A1(n1110), .B0(n1112), .B1(n75), .Y(n527) );
  OAI22XL U406 ( .A0(n1141), .A1(n592), .B0(n1162), .B1(n557), .Y(n599) );
  OAI22XL U407 ( .A0(n1089), .A1(n591), .B0(n1090), .B1(n554), .Y(n601) );
  OAI21X1 U408 ( .A0(n555), .A1(n556), .B0(n69), .Y(n600) );
  OAI22XL U409 ( .A0(n959), .A1(n631), .B0(n957), .B1(n598), .Y(n635) );
  OAI22XL U410 ( .A0(n967), .A1(n629), .B0(n965), .B1(n596), .Y(n637) );
  OAI22XL U411 ( .A0(n959), .A1(n598), .B0(n957), .B1(n563), .Y(n602) );
  OAI21XL U412 ( .A0(n285), .A1(n94), .B0(n284), .Y(n91) );
  NAND2X1 U413 ( .A(n78), .B(n217), .Y(n1223) );
  INVXL U414 ( .A(n1220), .Y(n1221) );
  AOI21XL U415 ( .A0(n1219), .A1(n1218), .B0(n1217), .Y(n1220) );
  INVXL U416 ( .A(n1233), .Y(n1217) );
  OAI2BB1XL U417 ( .A0N(n1138), .A1N(n1137), .B0(n1136), .Y(n1142) );
  OAI22XL U418 ( .A0(n1178), .A1(n1134), .B0(n1176), .B1(n1139), .Y(n1143) );
  INVXL U419 ( .A(n1135), .Y(n1136) );
  OAI22XL U420 ( .A0(n1178), .A1(n1109), .B0(n1176), .B1(n1134), .Y(n1132) );
  OAI22XL U421 ( .A0(n1141), .A1(n1108), .B0(n1162), .B1(n1130), .Y(n1133) );
  INVXL U422 ( .A(n1144), .Y(n1131) );
  OAI21XL U423 ( .A0(n61), .A1(n62), .B0(n60), .Y(n753) );
  INVXL U424 ( .A(n739), .Y(n61) );
  INVXL U425 ( .A(n254), .Y(n102) );
  OAI22XL U426 ( .A0(n959), .A1(n177), .B0(n957), .B1(n176), .Y(n187) );
  OAI22XL U427 ( .A0(n1141), .A1(n171), .B0(n1162), .B1(n170), .Y(n178) );
  OAI22XL U428 ( .A0(n959), .A1(n176), .B0(n957), .B1(n138), .Y(n181) );
  OAI22XL U429 ( .A0(n1112), .A1(n174), .B0(n1110), .B1(n137), .Y(n182) );
  OAI22XL U430 ( .A0(n1141), .A1(n417), .B0(n1162), .B1(n1093), .Y(n1096) );
  OAI22XL U431 ( .A0(n1178), .A1(n418), .B0(n1176), .B1(n1086), .Y(n1095) );
  INVXL U432 ( .A(n1106), .Y(n1094) );
  NOR2BXL U433 ( .AN(B[0]), .B(n965), .Y(n330) );
  OAI22XL U434 ( .A0(n963), .A1(n320), .B0(n961), .B1(n319), .Y(n328) );
  OAI22XL U435 ( .A0(n953), .A1(n318), .B0(n317), .B1(n1077), .Y(n329) );
  OAI22XL U436 ( .A0(n347), .A1(n302), .B0(n965), .B1(n301), .Y(n326) );
  OAI22XL U437 ( .A0(n963), .A1(n319), .B0(n961), .B1(n300), .Y(n327) );
  AOI21XL U438 ( .A0(n1229), .A1(n1228), .B0(n333), .Y(n1189) );
  INVXL U439 ( .A(n1227), .Y(n333) );
  ADDFX2 U440 ( .A(n281), .B(n280), .CI(n279), .CO(n343), .S(n342) );
  OAI21XL U441 ( .A0(n93), .A1(n92), .B0(n91), .Y(n280) );
  INVXL U442 ( .A(n285), .Y(n92) );
  OAI22XL U443 ( .A0(n1178), .A1(n1177), .B0(n1176), .B1(n1175), .Y(n1179) );
  OAI2BB1XL U444 ( .A0N(n1162), .A1N(n1161), .B0(n1160), .Y(n1171) );
  OAI22XL U445 ( .A0(n1178), .A1(n1158), .B0(n1176), .B1(n1177), .Y(n1172) );
  INVXL U446 ( .A(n1159), .Y(n1160) );
  OAI22XL U447 ( .A0(n953), .A1(B[0]), .B0(n305), .B1(n1077), .Y(n1212) );
  NAND2XL U448 ( .A(n306), .B(n953), .Y(n1211) );
  NAND2BXL U449 ( .AN(B[0]), .B(n518), .Y(n306) );
  INVXL U450 ( .A(n1204), .Y(n316) );
  NOR2XL U451 ( .A(n324), .B(n323), .Y(n1199) );
  NAND2XL U452 ( .A(n324), .B(n323), .Y(n1200) );
  NAND2XL U453 ( .A(n332), .B(n331), .Y(n1227) );
  INVXL U454 ( .A(n1189), .Y(n1197) );
  INVXL U455 ( .A(n433), .Y(n390) );
  NAND2XL U456 ( .A(n680), .B(n797), .Y(n682) );
  AOI21XL U457 ( .A0(n798), .A1(n680), .B0(n679), .Y(n681) );
  NAND2BXL U458 ( .AN(B[0]), .B(A[15]), .Y(n143) );
  XOR2XL U459 ( .A(B[23]), .B(n469), .Y(n73) );
  NAND2XL U460 ( .A(n1216), .B(n1123), .Y(n1125) );
  INVXL U461 ( .A(n1164), .Y(n1122) );
  AOI21XL U462 ( .A0(n1121), .A1(n1120), .B0(n1119), .Y(n1164) );
  INVXL U463 ( .A(n1237), .Y(n1119) );
  NAND2XL U464 ( .A(n1118), .B(n1120), .Y(n1163) );
  XNOR2X1 U465 ( .A(n1082), .B(n1081), .Y(PRODUCT[37]) );
  NAND2XL U466 ( .A(n1120), .B(n1237), .Y(n1081) );
  INVXL U467 ( .A(n1262), .Y(n758) );
  NAND2XL U468 ( .A(n1003), .B(n1282), .Y(n1004) );
  XNOR2XL U469 ( .A(n774), .B(B[14]), .Y(n696) );
  XNOR2XL U470 ( .A(n1129), .B(B[10]), .Y(n699) );
  XNOR2XL U471 ( .A(n1091), .B(B[12]), .Y(n704) );
  XNOR2XL U472 ( .A(n942), .B(n740), .Y(n705) );
  XNOR2XL U473 ( .A(n1129), .B(B[9]), .Y(n736) );
  XNOR2XL U474 ( .A(n942), .B(n781), .Y(n743) );
  XNOR2XL U475 ( .A(n774), .B(B[12]), .Y(n775) );
  XNOR2XL U476 ( .A(n1129), .B(B[8]), .Y(n777) );
  XNOR2XL U477 ( .A(n469), .B(n781), .Y(n239) );
  OAI22XL U478 ( .A0(n959), .A1(n958), .B0(n957), .B1(n956), .Y(n1017) );
  OAI22XL U479 ( .A0(n963), .A1(n367), .B0(n961), .B1(n962), .Y(n1009) );
  NOR2BXL U480 ( .AN(B[0]), .B(n1110), .Y(n360) );
  OAI22XL U481 ( .A0(n697), .A1(n354), .B0(n1090), .B1(n353), .Y(n358) );
  XNOR2XL U482 ( .A(B[25]), .B(n782), .Y(n478) );
  XNOR2XL U483 ( .A(n942), .B(B[23]), .Y(n480) );
  XNOR2XL U484 ( .A(n942), .B(B[22]), .Y(n484) );
  INVXL U485 ( .A(n550), .Y(n519) );
  XNOR2XL U486 ( .A(n782), .B(B[23]), .Y(n524) );
  XNOR2X1 U487 ( .A(n774), .B(B[18]), .Y(n554) );
  XNOR2XL U488 ( .A(n1129), .B(B[14]), .Y(n557) );
  XNOR2XL U489 ( .A(n1129), .B(B[13]), .Y(n592) );
  XNOR2XL U490 ( .A(n782), .B(B[21]), .Y(n596) );
  XNOR2X1 U491 ( .A(n942), .B(B[19]), .Y(n598) );
  XNOR2XL U492 ( .A(n782), .B(B[22]), .Y(n561) );
  XNOR2X1 U493 ( .A(n469), .B(n771), .Y(n272) );
  NAND2XL U494 ( .A(n1216), .B(n1215), .Y(n1166) );
  NAND2XL U495 ( .A(n537), .B(n211), .Y(n79) );
  INVXL U496 ( .A(n1241), .Y(n212) );
  OAI21XL U497 ( .A0(n1261), .A1(n1258), .B0(n1259), .Y(n122) );
  XNOR2XL U498 ( .A(n1091), .B(n1174), .Y(n1135) );
  OAI22XL U499 ( .A0(n1141), .A1(n656), .B0(n1162), .B1(n625), .Y(n663) );
  OAI22X1 U500 ( .A0(n963), .A1(n655), .B0(n961), .B1(n624), .Y(n664) );
  CMPR32X1 U501 ( .A(n668), .B(n667), .C(n666), .CO(n691), .S(n726) );
  OAI22XL U502 ( .A0(n1112), .A1(n661), .B0(n1110), .B1(n630), .Y(n667) );
  OAI22XL U503 ( .A0(n967), .A1(n660), .B0(n965), .B1(n629), .Y(n668) );
  CMPR32X1 U504 ( .A(n750), .B(n749), .C(n748), .CO(n766), .S(n804) );
  OAI22XL U505 ( .A0(n959), .A1(n743), .B0(n957), .B1(n705), .Y(n748) );
  OAI22X1 U506 ( .A0(n967), .A1(n741), .B0(n965), .B1(n703), .Y(n750) );
  OAI22XL U507 ( .A0(n1112), .A1(n742), .B0(n1110), .B1(n704), .Y(n749) );
  ADDFX2 U508 ( .A(n822), .B(n821), .CI(n820), .CO(n837), .S(n872) );
  OAI22XL U509 ( .A0(n959), .A1(n827), .B0(n957), .B1(n785), .Y(n832) );
  OAI22XL U510 ( .A0(n959), .A1(n828), .B0(n957), .B1(n827), .Y(n868) );
  OAI22XL U511 ( .A0(n1141), .A1(n819), .B0(n1162), .B1(n818), .Y(n865) );
  OAI2BB1XL U512 ( .A0N(n858), .A1N(n86), .B0(n84), .Y(n889) );
  AND2X1 U513 ( .A(n120), .B(n856), .Y(n890) );
  NAND2XL U514 ( .A(n85), .B(n857), .Y(n84) );
  AOI2BB1X2 U515 ( .A0N(n239), .A1N(n963), .B0(n88), .Y(n87) );
  NOR2X1 U516 ( .A(n817), .B(n961), .Y(n88) );
  OAI22X1 U517 ( .A0(n1089), .A1(n238), .B0(n1090), .B1(n815), .Y(n858) );
  NAND2XL U518 ( .A(n101), .B(n253), .Y(n100) );
  NAND2BXL U519 ( .AN(n254), .B(n103), .Y(n101) );
  NOR2X1 U520 ( .A(n169), .B(n963), .Y(n104) );
  OAI22XL U521 ( .A0(n959), .A1(n138), .B0(n957), .B1(n243), .Y(n235) );
  OAI22XL U522 ( .A0(n1112), .A1(n137), .B0(n1110), .B1(n242), .Y(n236) );
  XNOR2XL U523 ( .A(n774), .B(B[7]), .Y(n168) );
  XNOR2XL U524 ( .A(n1129), .B(B[3]), .Y(n171) );
  XNOR2XL U525 ( .A(n1091), .B(n941), .Y(n137) );
  XNOR2X1 U526 ( .A(n1091), .B(n771), .Y(n174) );
  XNOR2XL U527 ( .A(n942), .B(B[10]), .Y(n138) );
  XNOR2XL U528 ( .A(n942), .B(B[9]), .Y(n176) );
  CMPR32X1 U529 ( .A(n949), .B(n948), .C(n947), .CO(n938), .S(n988) );
  NOR2BXL U530 ( .AN(B[0]), .B(n1176), .Y(n195) );
  OAI22XL U531 ( .A0(n1141), .A1(n944), .B0(n1162), .B1(n151), .Y(n193) );
  CMPR32X1 U532 ( .A(n201), .B(n200), .C(n199), .CO(n940), .S(n971) );
  OAI22XL U533 ( .A0(n1112), .A1(n946), .B0(n1110), .B1(n175), .Y(n200) );
  OAI22XL U534 ( .A0(n1112), .A1(n954), .B0(n1110), .B1(n946), .Y(n974) );
  OAI22XL U535 ( .A0(n959), .A1(n956), .B0(n957), .B1(n943), .Y(n976) );
  OAI22XL U536 ( .A0(n1141), .A1(n945), .B0(n1162), .B1(n944), .Y(n975) );
  OAI22XL U537 ( .A0(n1089), .A1(n981), .B0(n1090), .B1(n980), .Y(n1023) );
  CMPR32X1 U538 ( .A(n357), .B(n356), .C(n355), .CO(n374), .S(n381) );
  OAI22XL U539 ( .A0(n967), .A1(n262), .B0(n965), .B1(n363), .Y(n355) );
  OAI22X1 U540 ( .A0(n1089), .A1(n261), .B0(n1090), .B1(n354), .Y(n356) );
  OAI22XL U541 ( .A0(n959), .A1(n268), .B0(n957), .B1(n361), .Y(n357) );
  OAI22XL U542 ( .A0(n963), .A1(n364), .B0(n961), .B1(n367), .Y(n368) );
  XNOR2X1 U543 ( .A(n1129), .B(n740), .Y(n513) );
  ADDFX2 U544 ( .A(n489), .B(n488), .CI(n487), .CO(n512), .S(n548) );
  OAI2BB1XL U545 ( .A0N(n556), .A1N(n735), .B0(n471), .Y(n487) );
  XNOR2XL U546 ( .A(n1129), .B(B[21]), .Y(n417) );
  OAI22XL U547 ( .A0(n1161), .A1(n409), .B0(n1162), .B1(n405), .Y(n413) );
  OAI22XL U548 ( .A0(n1161), .A1(n443), .B0(n1162), .B1(n409), .Y(n446) );
  CMPR32X1 U549 ( .A(n530), .B(n529), .C(n528), .CO(n549), .S(n583) );
  OAI22XL U550 ( .A0(n1089), .A1(n516), .B0(n1090), .B1(n486), .Y(n528) );
  OAI22X1 U551 ( .A0(n959), .A1(n514), .B0(n957), .B1(n484), .Y(n530) );
  OAI22XL U552 ( .A0(n1178), .A1(n517), .B0(n1176), .B1(n485), .Y(n529) );
  ADDFX2 U553 ( .A(n702), .B(n701), .CI(n700), .CO(n714), .S(n752) );
  XNOR2XL U554 ( .A(n518), .B(B[3]), .Y(n318) );
  OAI22XL U555 ( .A0(n967), .A1(n399), .B0(n965), .B1(n293), .Y(n303) );
  NAND2BXL U556 ( .AN(B[0]), .B(A[5]), .Y(n293) );
  XNOR2XL U557 ( .A(n469), .B(B[3]), .Y(n300) );
  NOR2BXL U558 ( .AN(B[0]), .B(n1090), .Y(n271) );
  OAI22XL U559 ( .A0(n959), .A1(n273), .B0(n957), .B1(n268), .Y(n269) );
  OAI22X1 U560 ( .A0(n953), .A1(n267), .B0(n266), .B1(n1077), .Y(n270) );
  NOR2BXL U561 ( .AN(B[0]), .B(n957), .Y(n296) );
  OAI22XL U562 ( .A0(n967), .A1(n301), .B0(n965), .B1(n287), .Y(n294) );
  XNOR2XL U563 ( .A(n942), .B(B[0]), .Y(n274) );
  OAI22XL U564 ( .A0(n959), .A1(n9), .B0(n957), .B1(n263), .Y(n282) );
  ADDFX2 U565 ( .A(n691), .B(n690), .CI(n689), .CO(n669), .S(n725) );
  ADDFX2 U566 ( .A(n885), .B(n884), .CI(n883), .CO(n871), .S(n904) );
  ADDFX2 U567 ( .A(n907), .B(n906), .CI(n905), .CO(n895), .S(n920) );
  NAND2X1 U568 ( .A(n185), .B(n186), .Y(n99) );
  NAND2X1 U569 ( .A(n110), .B(n109), .Y(n998) );
  OR2X2 U570 ( .A(n994), .B(n995), .Y(n111) );
  OAI22XL U571 ( .A0(n482), .A1(n1110), .B0(n1137), .B1(n76), .Y(n521) );
  OAI22XL U572 ( .A0(n1141), .A1(n1093), .B0(n1162), .B1(n1108), .Y(n1114) );
  OAI22XL U573 ( .A0(n1112), .A1(n1092), .B0(n1138), .B1(n1111), .Y(n1115) );
  OAI22XL U574 ( .A0(n1112), .A1(n420), .B0(n1138), .B1(n1092), .Y(n1099) );
  OAI2BB1XL U575 ( .A0N(n1090), .A1N(n1089), .B0(n1088), .Y(n1105) );
  OAI22XL U576 ( .A0(n1178), .A1(n1086), .B0(n1176), .B1(n1109), .Y(n1107) );
  INVXL U577 ( .A(n1087), .Y(n1088) );
  OAI22XL U578 ( .A0(n1089), .A1(n444), .B0(n1090), .B1(n439), .Y(n453) );
  OAI22XL U579 ( .A0(n1112), .A1(n410), .B0(n1110), .B1(n406), .Y(n416) );
  OAI22XL U580 ( .A0(n1178), .A1(n398), .B0(n1176), .B1(n402), .Y(n415) );
  CMPR32X1 U581 ( .A(n456), .B(n455), .C(n454), .CO(n457), .S(n496) );
  NAND2X1 U582 ( .A(n64), .B(n63), .Y(n638) );
  NAND2XL U583 ( .A(n650), .B(n649), .Y(n63) );
  NAND2X1 U584 ( .A(n65), .B(n648), .Y(n64) );
  OAI22XL U585 ( .A0(n953), .A1(n305), .B0(n309), .B1(n1077), .Y(n308) );
  NOR2BXL U586 ( .AN(B[0]), .B(n961), .Y(n307) );
  OAI22XL U587 ( .A0(n963), .A1(n312), .B0(n556), .B1(n311), .Y(n314) );
  NAND2BXL U588 ( .AN(B[0]), .B(n469), .Y(n311) );
  NAND2XL U589 ( .A(n1216), .B(n1222), .Y(n1225) );
  INVXL U590 ( .A(n1036), .Y(n1059) );
  OAI22XL U591 ( .A0(n1178), .A1(n1139), .B0(n1176), .B1(n1158), .Y(n1157) );
  INVXL U592 ( .A(n1173), .Y(n1156) );
  OAI22XL U593 ( .A0(n1141), .A1(n1130), .B0(n1162), .B1(n1140), .Y(n1152) );
  XOR3X2 U594 ( .A(n688), .B(n686), .C(n687), .Y(n716) );
  NAND2BXL U595 ( .AN(n794), .B(n82), .Y(n81) );
  NAND2X1 U596 ( .A(n107), .B(n106), .Y(n838) );
  OAI21XL U597 ( .A0(n105), .A1(n850), .B0(n848), .Y(n107) );
  BUFX1 U598 ( .A(n849), .Y(n105) );
  XOR2X1 U599 ( .A(n108), .B(n848), .Y(n875) );
  XOR2X1 U600 ( .A(n849), .B(n850), .Y(n108) );
  NAND2X1 U601 ( .A(n90), .B(n89), .Y(n874) );
  OAI21XL U602 ( .A0(n881), .A1(n882), .B0(n880), .Y(n90) );
  NAND2X1 U603 ( .A(n117), .B(n116), .Y(n898) );
  OAI21XL U604 ( .A0(n903), .A1(n904), .B0(n902), .Y(n117) );
  XOR2X1 U605 ( .A(n118), .B(n903), .Y(n915) );
  XNOR2X1 U606 ( .A(n902), .B(n119), .Y(n118) );
  OAI2BB1X1 U607 ( .A0N(n114), .A1N(n908), .B0(n113), .Y(n919) );
  NAND2XL U608 ( .A(n909), .B(n910), .Y(n113) );
  ADDFX2 U609 ( .A(n923), .B(n922), .CI(n921), .CO(n924), .S(n930) );
  XOR3X2 U610 ( .A(n184), .B(n186), .C(n185), .Y(n992) );
  XOR2X1 U611 ( .A(n112), .B(n993), .Y(n997) );
  ADDFX2 U612 ( .A(n1039), .B(n1038), .CI(n1037), .CO(n996), .S(n1049) );
  CMPR32X1 U613 ( .A(n1104), .B(n1103), .C(n1102), .CO(n1117), .S(n1100) );
  NAND2X1 U614 ( .A(n67), .B(n66), .Y(n672) );
  OR2X2 U615 ( .A(n687), .B(n688), .Y(n68) );
  NOR2XL U616 ( .A(n308), .B(n307), .Y(n1207) );
  NAND2XL U617 ( .A(n308), .B(n307), .Y(n1208) );
  NAND2XL U618 ( .A(n315), .B(n314), .Y(n1204) );
  NAND2XL U619 ( .A(n1154), .B(n1153), .Y(mult_x_1_n126) );
  NAND2XL U620 ( .A(n1074), .B(n1073), .Y(n1075) );
  NAND2XL U621 ( .A(n1065), .B(n1064), .Y(n1066) );
  OAI21XL U622 ( .A0(n1000), .A1(mult_x_1_n313), .B0(n1001), .Y(mult_x_1_n306)
         );
  NAND2XL U623 ( .A(n1183), .B(n1182), .Y(mult_x_1_n54) );
  NAND2XL U624 ( .A(n1181), .B(n1180), .Y(n1182) );
  INVXL U625 ( .A(n1179), .Y(n1180) );
  NOR2XL U626 ( .A(n1170), .B(n1169), .Y(mult_x_1_n105) );
  NAND2XL U627 ( .A(n1170), .B(n1169), .Y(mult_x_1_n106) );
  NOR2XL U628 ( .A(n1146), .B(n1145), .Y(mult_x_1_n114) );
  NAND2XL U629 ( .A(n1146), .B(n1145), .Y(mult_x_1_n115) );
  NOR2XL U630 ( .A(n1154), .B(n1153), .Y(mult_x_1_n125) );
  NOR2XL U631 ( .A(n1117), .B(n1116), .Y(mult_x_1_n134) );
  NAND2XL U632 ( .A(n1117), .B(n1116), .Y(mult_x_1_n135) );
  NAND2XL U633 ( .A(n1101), .B(n1100), .Y(mult_x_1_n150) );
  NOR2XL U634 ( .A(n1101), .B(n1100), .Y(mult_x_1_n149) );
  NOR2BXL U635 ( .AN(B[0]), .B(n1077), .Y(n1316) );
  XOR2XL U636 ( .A(n1210), .B(n1213), .Y(n1314) );
  NAND2XL U637 ( .A(n1209), .B(n1208), .Y(n1210) );
  INVXL U638 ( .A(n1207), .Y(n1209) );
  XNOR2XL U639 ( .A(n1206), .B(n1205), .Y(n1313) );
  NAND2XL U640 ( .A(n313), .B(n1204), .Y(n1206) );
  XOR2XL U641 ( .A(n1203), .B(n1202), .Y(n1312) );
  NAND2XL U642 ( .A(n1201), .B(n1200), .Y(n1203) );
  INVXL U643 ( .A(n1199), .Y(n1201) );
  NAND2XL U644 ( .A(n1228), .B(n1227), .Y(n1230) );
  NAND2XL U645 ( .A(n1196), .B(n1195), .Y(n1198) );
  XOR2XL U646 ( .A(n1194), .B(n1193), .Y(n1309) );
  NAND2XL U647 ( .A(n1192), .B(n1191), .Y(n1193) );
  NAND2XL U648 ( .A(n1186), .B(n1185), .Y(n1187) );
  INVXL U649 ( .A(n1184), .Y(n1186) );
  BUFX3 U650 ( .A(A[9]), .Y(n774) );
  BUFX3 U651 ( .A(A[7]), .Y(n942) );
  OAI21XL U652 ( .A0(n1265), .A1(n1262), .B0(n1263), .Y(n678) );
  NAND2X1 U653 ( .A(n98), .B(n96), .Y(n798) );
  BUFX3 U654 ( .A(A[11]), .Y(n1091) );
  OAI22X1 U655 ( .A0(n967), .A1(n478), .B0(n965), .B1(n400), .Y(n449) );
  OAI22X1 U656 ( .A0(n589), .A1(n146), .B0(n163), .B1(n1077), .Y(n166) );
  XNOR2X1 U657 ( .A(n769), .B(n740), .Y(n163) );
  OAI22X1 U658 ( .A0(n813), .A1(n622), .B0(n1176), .B1(n590), .Y(n619) );
  OAI22X1 U659 ( .A0(n1178), .A1(n695), .B0(n1176), .B1(n653), .Y(n692) );
  OAI22X1 U660 ( .A0(n959), .A1(n361), .B0(n957), .B1(n365), .Y(n370) );
  OAI22X1 U661 ( .A0(n1089), .A1(n815), .B0(n1090), .B1(n814), .Y(n867) );
  ADDFX2 U662 ( .A(n566), .B(n565), .CI(n564), .CO(n558), .S(n617) );
  OAI22X1 U663 ( .A0(n1178), .A1(n551), .B0(n1176), .B1(n517), .Y(n565) );
  NAND2BX1 U664 ( .AN(n858), .B(n87), .Y(n85) );
  OAI22X1 U665 ( .A0(n744), .A1(n408), .B0(n957), .B1(n403), .Y(n422) );
  BUFX1 U666 ( .A(n298), .Y(n59) );
  OAI22X1 U667 ( .A0(n1178), .A1(n590), .B0(n1176), .B1(n551), .Y(n586) );
  OAI22X1 U668 ( .A0(n1089), .A1(n814), .B0(n1090), .B1(n775), .Y(n831) );
  OAI22X1 U669 ( .A0(n963), .A1(n264), .B0(n961), .B1(n364), .Y(n373) );
  CMPR22X1 U670 ( .A(n252), .B(n251), .CO(n887), .S(n248) );
  XNOR2X1 U671 ( .A(n222), .B(n221), .Y(PRODUCT[36]) );
  AND2X1 U672 ( .A(n74), .B(n651), .Y(n658) );
  XOR2X1 U673 ( .A(n651), .B(n74), .Y(n702) );
  CMPR22X1 U674 ( .A(n166), .B(n165), .CO(n247), .S(n162) );
  XNOR3X2 U675 ( .A(n253), .B(n103), .C(n254), .Y(n256) );
  XNOR2X1 U676 ( .A(n782), .B(B[17]), .Y(n741) );
  OAI21XL U677 ( .A0(n739), .A1(n738), .B0(n737), .Y(n60) );
  XNOR3X2 U678 ( .A(n62), .B(n739), .C(n737), .Y(n793) );
  OR2X2 U679 ( .A(n650), .B(n649), .Y(n65) );
  XOR3X2 U680 ( .A(n649), .B(n650), .C(n648), .Y(n688) );
  XNOR2X1 U681 ( .A(B[20]), .B(n469), .Y(n698) );
  XOR2X1 U682 ( .A(n792), .B(n83), .Y(n801) );
  XOR2X1 U683 ( .A(n793), .B(n794), .Y(n83) );
  XNOR3X2 U684 ( .A(n857), .B(n87), .C(n858), .Y(n893) );
  XOR3X2 U685 ( .A(n285), .B(n94), .C(n284), .Y(n289) );
  OAI22X2 U686 ( .A0(n272), .A1(n961), .B0(n963), .B1(n291), .Y(n94) );
  NAND2BX1 U687 ( .AN(n337), .B(n95), .Y(n1192) );
  NOR2X1 U688 ( .A(n1266), .B(n1269), .Y(n97) );
  OAI21X2 U689 ( .A0(n1273), .A1(n1270), .B0(n1271), .Y(n841) );
  XOR2X1 U690 ( .A(n120), .B(n856), .Y(n888) );
  OAI22X1 U691 ( .A0(n810), .A1(n1077), .B0(n249), .B1(n953), .Y(n120) );
  OAI22X1 U692 ( .A0(n735), .A1(n698), .B0(n961), .B1(n655), .Y(n707) );
  NAND2X2 U693 ( .A(n123), .B(n121), .Y(n208) );
  AOI21X1 U694 ( .A0(n206), .A1(n678), .B0(n122), .Y(n121) );
  XOR2X1 U695 ( .A(n570), .B(n125), .Y(n580) );
  XOR2X1 U696 ( .A(n571), .B(n572), .Y(n125) );
  NAND2X1 U697 ( .A(n999), .B(n998), .Y(n1001) );
  OAI22X1 U698 ( .A0(n953), .A1(n731), .B0(n694), .B1(n1077), .Y(n730) );
  OAI22X1 U699 ( .A0(n735), .A1(n734), .B0(n961), .B1(n698), .Y(n746) );
  CMPR22X1 U700 ( .A(n587), .B(n586), .CO(n595), .S(n628) );
  OAI22X1 U701 ( .A0(n589), .A1(n588), .B0(n550), .B1(n1077), .Y(n587) );
  OAI22X1 U702 ( .A0(n953), .A1(n157), .B0(n145), .B1(n1077), .Y(n194) );
  OAI22X1 U703 ( .A0(n953), .A1(n145), .B0(n146), .B1(n1077), .Y(n148) );
  OAI22X1 U704 ( .A0(n1089), .A1(n696), .B0(n1090), .B1(n654), .Y(n708) );
  CMPR22X1 U705 ( .A(n951), .B(n950), .CO(n947), .S(n1008) );
  OAI22X1 U706 ( .A0(n953), .A1(n952), .B0(n157), .B1(n1077), .Y(n951) );
  OAI22X1 U707 ( .A0(n959), .A1(n480), .B0(n957), .B1(n441), .Y(n476) );
  OAI21X1 U708 ( .A0(n1254), .A1(n1257), .B0(n1255), .Y(n537) );
  AOI21XL U709 ( .A0(n1223), .A1(n1118), .B0(n1121), .Y(n1079) );
  XNOR2XL U710 ( .A(A[15]), .B(B[0]), .Y(n150) );
  OAI22X1 U711 ( .A0(n1089), .A1(n554), .B0(n1090), .B1(n516), .Y(n566) );
  AOI21XL U712 ( .A0(n1205), .A1(n313), .B0(n316), .Y(n1202) );
  XOR2XL U713 ( .A(A[4]), .B(A[5]), .Y(n126) );
  XNOR2XL U714 ( .A(A[4]), .B(A[3]), .Y(n127) );
  BUFX3 U715 ( .A(n347), .Y(n967) );
  BUFX3 U716 ( .A(B[11]), .Y(n773) );
  XNOR2X1 U717 ( .A(A[5]), .B(n773), .Y(n139) );
  BUFX3 U718 ( .A(n127), .Y(n965) );
  XNOR2X1 U719 ( .A(A[5]), .B(B[12]), .Y(n136) );
  OAI22XL U720 ( .A0(n967), .A1(n139), .B0(n965), .B1(n136), .Y(n183) );
  XOR2XL U721 ( .A(A[10]), .B(A[11]), .Y(n128) );
  NAND2X1 U722 ( .A(n128), .B(n1138), .Y(n1137) );
  BUFX3 U723 ( .A(n1137), .Y(n1112) );
  BUFX3 U724 ( .A(B[5]), .Y(n771) );
  BUFX3 U725 ( .A(n1138), .Y(n1110) );
  BUFX3 U726 ( .A(B[6]), .Y(n941) );
  XOR2XL U727 ( .A(A[6]), .B(A[7]), .Y(n129) );
  XNOR2XL U728 ( .A(A[6]), .B(A[5]), .Y(n130) );
  NAND2X1 U729 ( .A(n129), .B(n130), .Y(n744) );
  BUFX3 U730 ( .A(n744), .Y(n959) );
  BUFX3 U731 ( .A(n130), .Y(n957) );
  XOR2XL U732 ( .A(A[8]), .B(A[9]), .Y(n131) );
  BUFX3 U733 ( .A(n697), .Y(n1089) );
  BUFX3 U734 ( .A(n132), .Y(n1090) );
  OAI22X1 U735 ( .A0(n1089), .A1(n167), .B0(n1090), .B1(n238), .Y(n254) );
  XOR2XL U736 ( .A(A[2]), .B(A[3]), .Y(n133) );
  NAND2X1 U737 ( .A(n133), .B(n556), .Y(n735) );
  BUFX3 U738 ( .A(n735), .Y(n963) );
  BUFX3 U739 ( .A(n556), .Y(n961) );
  INVXL U740 ( .A(n469), .Y(n312) );
  BUFX3 U741 ( .A(B[15]), .Y(n781) );
  XOR2XL U742 ( .A(A[12]), .B(A[13]), .Y(n134) );
  XNOR2XL U743 ( .A(A[12]), .B(A[11]), .Y(n135) );
  NAND2X1 U744 ( .A(n134), .B(n135), .Y(n1161) );
  BUFX3 U745 ( .A(n1161), .Y(n1141) );
  XNOR2XL U746 ( .A(n1129), .B(B[4]), .Y(n170) );
  BUFX3 U747 ( .A(n135), .Y(n1162) );
  OAI22X1 U748 ( .A0(n1141), .A1(n170), .B0(n1162), .B1(n240), .Y(n253) );
  OAI22XL U749 ( .A0(n967), .A1(n136), .B0(n965), .B1(n241), .Y(n237) );
  XNOR2X1 U750 ( .A(A[5]), .B(B[10]), .Y(n156) );
  OAI22XL U751 ( .A0(n967), .A1(n156), .B0(n965), .B1(n139), .Y(n192) );
  NAND2X1 U752 ( .A(A[1]), .B(n140), .Y(n589) );
  BUFX3 U753 ( .A(n589), .Y(n953) );
  XNOR2X1 U754 ( .A(n518), .B(B[14]), .Y(n145) );
  XNOR2X1 U755 ( .A(n769), .B(B[15]), .Y(n146) );
  BUFX3 U756 ( .A(n140), .Y(n1077) );
  XOR2XL U757 ( .A(A[14]), .B(A[15]), .Y(n141) );
  XNOR2XL U758 ( .A(A[14]), .B(A[13]), .Y(n142) );
  NAND2X1 U759 ( .A(n141), .B(n142), .Y(n813) );
  BUFX3 U760 ( .A(n813), .Y(n1178) );
  BUFX3 U761 ( .A(n142), .Y(n1176) );
  OAI22X1 U762 ( .A0(n1178), .A1(n144), .B0(n1176), .B1(n143), .Y(n147) );
  XNOR2X1 U763 ( .A(n518), .B(B[13]), .Y(n157) );
  XNOR2XL U764 ( .A(n1129), .B(B[1]), .Y(n944) );
  XNOR2XL U765 ( .A(n1129), .B(B[2]), .Y(n151) );
  BUFX3 U766 ( .A(B[16]), .Y(n740) );
  XNOR2XL U767 ( .A(A[15]), .B(B[1]), .Y(n149) );
  XNOR2XL U768 ( .A(A[15]), .B(B[2]), .Y(n164) );
  OAI22X1 U769 ( .A0(n1178), .A1(n149), .B0(n1176), .B1(n164), .Y(n165) );
  CMPR22X1 U770 ( .A(n148), .B(n147), .CO(n161), .S(n191) );
  XNOR2X1 U771 ( .A(n774), .B(n941), .Y(n152) );
  OAI22XL U772 ( .A0(n697), .A1(n152), .B0(n1090), .B1(n168), .Y(n155) );
  OAI22XL U773 ( .A0(n697), .A1(n196), .B0(n1090), .B1(n152), .Y(n201) );
  XNOR2X2 U774 ( .A(n469), .B(n773), .Y(n197) );
  OAI22XL U775 ( .A0(n963), .A1(n197), .B0(n961), .B1(n173), .Y(n199) );
  CMPR32X1 U776 ( .A(n155), .B(n154), .C(n153), .CO(n160), .S(n939) );
  XNOR2X1 U777 ( .A(A[5]), .B(B[9]), .Y(n198) );
  OAI22XL U778 ( .A0(n967), .A1(n198), .B0(n965), .B1(n156), .Y(n949) );
  OAI22XL U779 ( .A0(n959), .A1(n943), .B0(n957), .B1(n177), .Y(n948) );
  XNOR2X1 U780 ( .A(n518), .B(B[12]), .Y(n952) );
  OAI22X1 U781 ( .A0(n1141), .A1(n159), .B0(n1162), .B1(n158), .Y(n950) );
  CMPR32X1 U782 ( .A(n162), .B(n161), .C(n160), .CO(n245), .S(n203) );
  OAI22X1 U783 ( .A0(n589), .A1(n163), .B0(n249), .B1(n1077), .Y(n252) );
  XNOR2X1 U784 ( .A(A[15]), .B(B[3]), .Y(n250) );
  OAI22X1 U785 ( .A0(n1178), .A1(n164), .B0(n1176), .B1(n250), .Y(n251) );
  OAI22XL U786 ( .A0(n1089), .A1(n168), .B0(n1090), .B1(n167), .Y(n180) );
  OAI22XL U787 ( .A0(n963), .A1(n173), .B0(n961), .B1(n172), .Y(n189) );
  OAI22X1 U788 ( .A0(n1112), .A1(n175), .B0(n1110), .B1(n174), .Y(n188) );
  CMPR32X1 U789 ( .A(n180), .B(n179), .C(n178), .CO(n246), .S(n185) );
  CMPR32X1 U790 ( .A(n183), .B(n182), .C(n181), .CO(n257), .S(n184) );
  CMPR32X1 U791 ( .A(n189), .B(n188), .C(n187), .CO(n186), .S(n970) );
  CMPR32X1 U792 ( .A(n192), .B(n191), .C(n190), .CO(n204), .S(n969) );
  ADDFHX1 U793 ( .A(n195), .B(n194), .CI(n193), .CO(n190), .S(n973) );
  XNOR2XL U794 ( .A(n774), .B(B[4]), .Y(n980) );
  OAI22XL U795 ( .A0(n1089), .A1(n980), .B0(n1090), .B1(n196), .Y(n979) );
  XNOR2X1 U796 ( .A(n469), .B(B[10]), .Y(n960) );
  XNOR2X1 U797 ( .A(A[5]), .B(B[8]), .Y(n964) );
  OAI22XL U798 ( .A0(n347), .A1(n964), .B0(n965), .B1(n198), .Y(n977) );
  NOR2X1 U799 ( .A(n935), .B(n934), .Y(mult_x_1_n302) );
  NOR2X1 U800 ( .A(n1260), .B(n1258), .Y(n206) );
  NOR2X1 U801 ( .A(n677), .B(n207), .Y(n209) );
  NOR2XL U802 ( .A(n1252), .B(n1250), .Y(n211) );
  NAND2XL U803 ( .A(n395), .B(n232), .Y(n214) );
  NOR2XL U804 ( .A(n1244), .B(n214), .Y(n216) );
  NAND2XL U805 ( .A(n223), .B(n216), .Y(n218) );
  NOR2XL U806 ( .A(n503), .B(n218), .Y(n1078) );
  OAI21XL U807 ( .A0(n1250), .A1(n1253), .B0(n1251), .Y(n210) );
  OAI21XL U808 ( .A0(n1246), .A1(n1249), .B0(n1247), .Y(n433) );
  INVXL U809 ( .A(n1243), .Y(n224) );
  AOI21XL U810 ( .A0(n232), .A1(n224), .B0(n212), .Y(n213) );
  OAI21XL U811 ( .A0(n214), .A1(n1245), .B0(n213), .Y(n215) );
  AOI21XL U812 ( .A0(n433), .A1(n216), .B0(n215), .Y(n217) );
  INVXL U813 ( .A(n1223), .Y(n219) );
  INVXL U814 ( .A(n223), .Y(n432) );
  INVXL U815 ( .A(n1244), .Y(n436) );
  NAND2XL U816 ( .A(n436), .B(n395), .Y(n227) );
  NOR2XL U817 ( .A(n432), .B(n227), .Y(n229) );
  NAND2XL U818 ( .A(n6), .B(n229), .Y(n231) );
  AOI21XL U819 ( .A0(n225), .A1(n395), .B0(n224), .Y(n226) );
  OAI21XL U820 ( .A0(n390), .A1(n227), .B0(n226), .Y(n228) );
  CMPR32X1 U821 ( .A(n237), .B(n236), .C(n235), .CO(n894), .S(n255) );
  OAI22X1 U822 ( .A0(n1141), .A1(n240), .B0(n1162), .B1(n819), .Y(n857) );
  XNOR2X1 U823 ( .A(A[5]), .B(B[14]), .Y(n824) );
  OAI22XL U824 ( .A0(n967), .A1(n241), .B0(n965), .B1(n824), .Y(n864) );
  XNOR2X1 U825 ( .A(n769), .B(B[18]), .Y(n810) );
  XNOR2XL U826 ( .A(A[15]), .B(B[4]), .Y(n812) );
  OAI22X1 U827 ( .A0(n1178), .A1(n250), .B0(n1176), .B1(n812), .Y(n856) );
  CMPR32X1 U828 ( .A(n257), .B(n256), .C(n255), .CO(n908), .S(n260) );
  CMPR32X1 U829 ( .A(n260), .B(n259), .C(n258), .CO(n929), .S(n935) );
  XNOR2XL U830 ( .A(n942), .B(B[2]), .Y(n268) );
  XNOR2XL U831 ( .A(n774), .B(B[0]), .Y(n261) );
  XNOR2XL U832 ( .A(n774), .B(B[1]), .Y(n354) );
  XNOR2X1 U833 ( .A(A[5]), .B(B[4]), .Y(n262) );
  XNOR2X1 U834 ( .A(A[5]), .B(n771), .Y(n363) );
  XNOR2X1 U835 ( .A(n469), .B(n941), .Y(n264) );
  OAI22XL U836 ( .A0(n963), .A1(n272), .B0(n961), .B1(n264), .Y(n278) );
  XNOR2X1 U837 ( .A(A[5]), .B(B[3]), .Y(n275) );
  OAI22XL U838 ( .A0(n347), .A1(n275), .B0(n965), .B1(n262), .Y(n277) );
  XNOR2X1 U839 ( .A(n518), .B(B[6]), .Y(n286) );
  XNOR2X1 U840 ( .A(n518), .B(B[7]), .Y(n267) );
  OAI22XL U841 ( .A0(n953), .A1(n286), .B0(n267), .B1(n1077), .Y(n283) );
  XNOR2X1 U842 ( .A(n518), .B(B[8]), .Y(n266) );
  OAI22X1 U843 ( .A0(n1089), .A1(n7), .B0(n1090), .B1(n265), .Y(n349) );
  XNOR2XL U844 ( .A(n942), .B(B[1]), .Y(n273) );
  CMPR32X1 U845 ( .A(n271), .B(n270), .C(n269), .CO(n371), .S(n281) );
  XNOR2XL U846 ( .A(n469), .B(B[4]), .Y(n291) );
  OAI22X1 U847 ( .A0(n959), .A1(n274), .B0(n957), .B1(n273), .Y(n285) );
  XNOR2XL U848 ( .A(A[5]), .B(B[2]), .Y(n287) );
  OAI22X1 U849 ( .A0(n967), .A1(n287), .B0(n965), .B1(n275), .Y(n284) );
  CMPR32X1 U850 ( .A(n278), .B(n277), .C(n276), .CO(n380), .S(n279) );
  ADDHXL U851 ( .A(n283), .B(n282), .CO(n276), .S(n290) );
  XNOR2X1 U852 ( .A(n518), .B(n771), .Y(n292) );
  OAI22XL U853 ( .A0(n953), .A1(n292), .B0(n286), .B1(n1077), .Y(n295) );
  XNOR2XL U854 ( .A(A[5]), .B(B[1]), .Y(n301) );
  CMPR32X1 U855 ( .A(n288), .B(n289), .C(n290), .CO(n341), .S(n337) );
  XNOR2XL U856 ( .A(n518), .B(B[4]), .Y(n317) );
  OAI22XL U857 ( .A0(n953), .A1(n317), .B0(n292), .B1(n1077), .Y(n304) );
  CMPR32X1 U858 ( .A(n296), .B(n295), .C(n294), .CO(n288), .S(n297) );
  XNOR2XL U859 ( .A(n469), .B(B[2]), .Y(n319) );
  XNOR2XL U860 ( .A(A[5]), .B(B[0]), .Y(n302) );
  ADDHXL U861 ( .A(n304), .B(n303), .CO(n298), .S(n325) );
  OR2X2 U862 ( .A(n335), .B(n334), .Y(n1196) );
  XNOR2XL U863 ( .A(n518), .B(B[1]), .Y(n305) );
  XNOR2XL U864 ( .A(n518), .B(B[2]), .Y(n309) );
  OAI21XL U865 ( .A0(n1207), .A1(n1213), .B0(n1208), .Y(n1205) );
  OAI22X1 U866 ( .A0(n953), .A1(n309), .B0(n318), .B1(n1077), .Y(n322) );
  XNOR2XL U867 ( .A(n469), .B(B[0]), .Y(n310) );
  XNOR2XL U868 ( .A(n469), .B(B[1]), .Y(n320) );
  OAI22X1 U869 ( .A0(n963), .A1(n310), .B0(n961), .B1(n320), .Y(n321) );
  CMPR22X1 U870 ( .A(n322), .B(n321), .CO(n323), .S(n315) );
  OAI21XL U871 ( .A0(n1202), .A1(n1199), .B0(n1200), .Y(n1229) );
  CMPR32X1 U872 ( .A(n327), .B(n326), .C(n325), .CO(n334), .S(n332) );
  CMPR32X1 U873 ( .A(n330), .B(n329), .C(n328), .CO(n331), .S(n324) );
  OR2X2 U874 ( .A(n332), .B(n331), .Y(n1228) );
  NAND2XL U875 ( .A(n335), .B(n334), .Y(n1195) );
  INVXL U876 ( .A(n1195), .Y(n1190) );
  NAND2XL U877 ( .A(n337), .B(n336), .Y(n1191) );
  INVXL U878 ( .A(n1191), .Y(n338) );
  NAND2XL U879 ( .A(n344), .B(n343), .Y(n1073) );
  AOI21X1 U880 ( .A0(n346), .A1(n1071), .B0(n345), .Y(n1062) );
  XNOR2X1 U881 ( .A(A[5]), .B(n941), .Y(n362) );
  XNOR2X1 U882 ( .A(A[5]), .B(B[7]), .Y(n966) );
  OAI22XL U883 ( .A0(n347), .A1(n362), .B0(n965), .B1(n966), .Y(n1014) );
  XNOR2XL U884 ( .A(n774), .B(B[2]), .Y(n353) );
  OAI22XL U885 ( .A0(n1089), .A1(n353), .B0(n1090), .B1(n981), .Y(n1013) );
  OAI22X1 U886 ( .A0(n1112), .A1(n77), .B0(n1110), .B1(n348), .Y(n982) );
  CMPR22X1 U887 ( .A(n350), .B(n349), .CO(n376), .S(n372) );
  OAI22X1 U888 ( .A0(n953), .A1(n352), .B0(n351), .B1(n1077), .Y(n359) );
  ADDFHX1 U889 ( .A(n360), .B(n359), .CI(n358), .CO(n1026), .S(n375) );
  OAI22X1 U890 ( .A0(n967), .A1(n363), .B0(n965), .B1(n362), .Y(n369) );
  OAI22XL U891 ( .A0(n959), .A1(n365), .B0(n957), .B1(n958), .Y(n1011) );
  OAI22XL U892 ( .A0(n1112), .A1(n366), .B0(n1110), .B1(n955), .Y(n1010) );
  CMPR32X1 U893 ( .A(n381), .B(n380), .C(n379), .CO(n383), .S(n344) );
  NAND2XL U894 ( .A(n1065), .B(n382), .Y(n389) );
  INVXL U895 ( .A(n1068), .Y(n1063) );
  INVXL U896 ( .A(n1064), .Y(n387) );
  AOI21XL U897 ( .A0(n1065), .A1(n1063), .B0(n387), .Y(n388) );
  OAI21XL U898 ( .A0(n1062), .A1(n389), .B0(n388), .Y(mult_x_1_n335) );
  NOR2XL U899 ( .A(n432), .B(n1244), .Y(n392) );
  NAND2XL U900 ( .A(n6), .B(n392), .Y(n394) );
  OAI21XL U901 ( .A0(n390), .A1(n1244), .B0(n1245), .Y(n391) );
  XNOR2X1 U902 ( .A(n397), .B(n396), .Y(PRODUCT[34]) );
  XNOR2X1 U903 ( .A(A[15]), .B(B[17]), .Y(n398) );
  XNOR2X1 U904 ( .A(A[15]), .B(B[18]), .Y(n402) );
  XNOR2X1 U905 ( .A(A[15]), .B(n740), .Y(n442) );
  BUFX3 U906 ( .A(B[26]), .Y(n1174) );
  XNOR2X1 U907 ( .A(A[5]), .B(n1174), .Y(n400) );
  OAI22XL U908 ( .A0(n1089), .A1(n439), .B0(n1090), .B1(n407), .Y(n412) );
  INVXL U909 ( .A(n422), .Y(n411) );
  XNOR2X1 U910 ( .A(A[15]), .B(B[19]), .Y(n418) );
  OAI22XL U911 ( .A0(n1137), .A1(n406), .B0(n1110), .B1(n420), .Y(n425) );
  XNOR2X1 U912 ( .A(n942), .B(B[24]), .Y(n441) );
  OAI22XL U913 ( .A0(n959), .A1(n441), .B0(n957), .B1(n408), .Y(n447) );
  XNOR2X1 U914 ( .A(n1091), .B(B[20]), .Y(n440) );
  OAI22XL U915 ( .A0(n1112), .A1(n440), .B0(n1110), .B1(n410), .Y(n445) );
  CMPR32X1 U916 ( .A(n413), .B(n412), .C(n411), .CO(n429), .S(n455) );
  CMPR32X1 U917 ( .A(n416), .B(n415), .C(n414), .CO(n459), .S(n454) );
  XNOR2X1 U918 ( .A(A[15]), .B(B[20]), .Y(n1086) );
  OAI22X1 U919 ( .A0(n1089), .A1(n419), .B0(n1090), .B1(n1087), .Y(n1106) );
  CMPR32X1 U920 ( .A(n423), .B(n422), .C(n421), .CO(n1098), .S(n428) );
  CMPR32X1 U921 ( .A(n426), .B(n425), .C(n424), .CO(n1097), .S(n427) );
  CMPR32X1 U922 ( .A(n429), .B(n428), .C(n427), .CO(n1083), .S(n458) );
  NOR2XL U923 ( .A(n431), .B(n430), .Y(mult_x_1_n162) );
  NAND2XL U924 ( .A(n431), .B(n430), .Y(mult_x_1_n163) );
  NAND2XL U925 ( .A(n6), .B(n223), .Y(n435) );
  AOI21XL U926 ( .A0(n501), .A1(n223), .B0(n433), .Y(n434) );
  OAI22XL U927 ( .A0(n1137), .A1(n482), .B0(n1110), .B1(n440), .Y(n477) );
  INVXL U928 ( .A(n449), .Y(n475) );
  OAI22XL U929 ( .A0(n1178), .A1(n468), .B0(n1176), .B1(n442), .Y(n474) );
  XNOR2X1 U930 ( .A(n1129), .B(B[17]), .Y(n479) );
  OAI22XL U931 ( .A0(n1161), .A1(n479), .B0(n1162), .B1(n443), .Y(n473) );
  CMPR32X1 U932 ( .A(n447), .B(n446), .C(n445), .CO(n456), .S(n495) );
  CMPR32X1 U933 ( .A(n450), .B(n449), .C(n448), .CO(n414), .S(n494) );
  ADDFHX1 U934 ( .A(n453), .B(n452), .CI(n451), .CO(n498), .S(n493) );
  CMPR32X1 U935 ( .A(n459), .B(n458), .C(n457), .CO(n431), .S(n460) );
  NOR2XL U936 ( .A(n461), .B(n460), .Y(mult_x_1_n173) );
  NAND2XL U937 ( .A(n461), .B(n460), .Y(mult_x_1_n174) );
  NAND2XL U938 ( .A(n6), .B(n504), .Y(n464) );
  XNOR2X2 U939 ( .A(n467), .B(n466), .Y(PRODUCT[32]) );
  XNOR2X1 U940 ( .A(A[15]), .B(B[14]), .Y(n485) );
  OAI22XL U941 ( .A0(n1178), .A1(n485), .B0(n1176), .B1(n468), .Y(n489) );
  XNOR2X1 U942 ( .A(n469), .B(n1174), .Y(n470) );
  INVXL U943 ( .A(n470), .Y(n471) );
  CMPR32X1 U944 ( .A(n474), .B(n473), .C(n472), .CO(n451), .S(n511) );
  CMPR32X1 U945 ( .A(n477), .B(n476), .C(n475), .CO(n452), .S(n510) );
  XNOR2X1 U946 ( .A(n782), .B(B[24]), .Y(n483) );
  OAI22XL U947 ( .A0(n967), .A1(n483), .B0(n965), .B1(n478), .Y(n492) );
  OAI22XL U948 ( .A0(n1141), .A1(n513), .B0(n1162), .B1(n479), .Y(n491) );
  OAI22XL U949 ( .A0(n959), .A1(n484), .B0(n957), .B1(n480), .Y(n490) );
  OAI22XL U950 ( .A0(n1089), .A1(n486), .B0(n1090), .B1(n481), .Y(n522) );
  OAI22X2 U951 ( .A0(n967), .A1(n524), .B0(n965), .B1(n483), .Y(n526) );
  INVXL U952 ( .A(n488), .Y(n525) );
  XNOR2X1 U953 ( .A(A[15]), .B(B[13]), .Y(n517) );
  XNOR2X1 U954 ( .A(n774), .B(B[19]), .Y(n516) );
  CMPR32X1 U955 ( .A(n492), .B(n491), .C(n490), .CO(n533), .S(n547) );
  CMPR32X1 U956 ( .A(n498), .B(n497), .C(n496), .CO(n461), .S(n499) );
  NOR2XL U957 ( .A(n500), .B(n499), .Y(mult_x_1_n184) );
  NAND2XL U958 ( .A(n500), .B(n499), .Y(mult_x_1_n185) );
  XNOR2X2 U959 ( .A(n506), .B(n505), .Y(PRODUCT[31]) );
  CMPR32X1 U960 ( .A(n512), .B(n511), .C(n510), .CO(n509), .S(n546) );
  XNOR2X1 U961 ( .A(n1129), .B(n781), .Y(n515) );
  OAI22XL U962 ( .A0(n1141), .A1(n557), .B0(n1162), .B1(n515), .Y(n552) );
  XNOR2X1 U963 ( .A(A[15]), .B(B[12]), .Y(n551) );
  CMPR32X1 U964 ( .A(n522), .B(n521), .C(n520), .CO(n532), .S(n571) );
  XNOR2X1 U965 ( .A(n469), .B(B[24]), .Y(n555) );
  OAI22X1 U966 ( .A0(n963), .A1(n555), .B0(n556), .B1(n523), .Y(n569) );
  XNOR2X1 U967 ( .A(n1091), .B(n740), .Y(n562) );
  OAI22XL U968 ( .A0(n967), .A1(n561), .B0(n965), .B1(n524), .Y(n567) );
  NOR2XL U969 ( .A(n535), .B(n534), .Y(mult_x_1_n191) );
  NAND2XL U970 ( .A(n535), .B(n534), .Y(mult_x_1_n192) );
  INVXL U971 ( .A(n536), .Y(n576) );
  NAND2XL U972 ( .A(n536), .B(n577), .Y(n540) );
  AOI21XL U973 ( .A0(n537), .A1(n577), .B0(n538), .Y(n539) );
  INVXL U974 ( .A(n1250), .Y(n541) );
  XNOR2X2 U975 ( .A(n543), .B(n542), .Y(PRODUCT[30]) );
  CMPR32X1 U976 ( .A(n546), .B(n545), .C(n544), .CO(n534), .S(n574) );
  CMPR32X1 U977 ( .A(n549), .B(n548), .C(n547), .CO(n531), .S(n582) );
  XNOR2X1 U978 ( .A(n769), .B(B[25]), .Y(n588) );
  XNOR2X1 U979 ( .A(A[15]), .B(n773), .Y(n590) );
  CMPR32X1 U980 ( .A(n560), .B(n559), .C(n558), .CO(n572), .S(n606) );
  OAI22X1 U981 ( .A0(n967), .A1(n596), .B0(n965), .B1(n561), .Y(n604) );
  XNOR2X1 U982 ( .A(n1091), .B(n781), .Y(n597) );
  OAI22XL U983 ( .A0(n1112), .A1(n597), .B0(n1110), .B1(n562), .Y(n603) );
  NOR2XL U984 ( .A(n574), .B(n573), .Y(mult_x_1_n202) );
  NAND2XL U985 ( .A(n574), .B(n573), .Y(mult_x_1_n203) );
  INVXL U986 ( .A(n537), .Y(n575) );
  CMPR32X1 U987 ( .A(n582), .B(n581), .C(n580), .CO(n573), .S(n609) );
  CMPR32X1 U988 ( .A(n585), .B(n584), .C(n583), .CO(n570), .S(n615) );
  XNOR2X1 U989 ( .A(n769), .B(B[24]), .Y(n621) );
  OAI22X1 U990 ( .A0(n589), .A1(n621), .B0(n588), .B1(n1077), .Y(n620) );
  XNOR2X1 U991 ( .A(A[15]), .B(B[10]), .Y(n622) );
  OAI22XL U992 ( .A0(n1089), .A1(n623), .B0(n1090), .B1(n591), .Y(n634) );
  XNOR2X1 U993 ( .A(n782), .B(B[20]), .Y(n629) );
  OAI22XL U994 ( .A0(n1112), .A1(n630), .B0(n1110), .B1(n597), .Y(n636) );
  ADDFHX1 U995 ( .A(n601), .B(n600), .CI(n599), .CO(n593), .S(n649) );
  CMPR32X1 U996 ( .A(n604), .B(n603), .C(n602), .CO(n618), .S(n648) );
  NOR2XL U997 ( .A(n609), .B(n608), .Y(mult_x_1_n209) );
  NAND2XL U998 ( .A(n609), .B(n608), .Y(mult_x_1_n210) );
  INVXL U999 ( .A(n1254), .Y(n610) );
  NAND2X1 U1000 ( .A(n610), .B(n1255), .Y(n611) );
  CMPR32X1 U1001 ( .A(n615), .B(n614), .C(n613), .CO(n608), .S(n642) );
  CMPR32X1 U1002 ( .A(n618), .B(n617), .C(n616), .CO(n605), .S(n647) );
  CMPR22X1 U1003 ( .A(n620), .B(n619), .CO(n627), .S(n659) );
  XNOR2X1 U1004 ( .A(n769), .B(B[23]), .Y(n652) );
  XNOR2X1 U1005 ( .A(A[15]), .B(B[9]), .Y(n653) );
  OAI22XL U1006 ( .A0(n813), .A1(n653), .B0(n1176), .B1(n622), .Y(n651) );
  XNOR2X1 U1007 ( .A(n774), .B(n781), .Y(n654) );
  OAI22XL U1008 ( .A0(n1089), .A1(n654), .B0(n1090), .B1(n623), .Y(n665) );
  OAI22XL U1009 ( .A0(n744), .A1(n662), .B0(n957), .B1(n631), .Y(n666) );
  CMPR32X1 U1010 ( .A(n637), .B(n636), .C(n635), .CO(n650), .S(n689) );
  NOR2XL U1011 ( .A(n642), .B(n641), .Y(mult_x_1_n220) );
  NAND2XL U1012 ( .A(n642), .B(n641), .Y(mult_x_1_n221) );
  XNOR2X1 U1013 ( .A(n769), .B(B[22]), .Y(n694) );
  OAI22X1 U1014 ( .A0(n953), .A1(n694), .B0(n652), .B1(n1077), .Y(n693) );
  XNOR2X1 U1015 ( .A(A[15]), .B(B[8]), .Y(n695) );
  ADDFHX1 U1016 ( .A(n665), .B(n664), .CI(n663), .CO(n657), .S(n727) );
  NOR2XL U1017 ( .A(n673), .B(n672), .Y(mult_x_1_n223) );
  NAND2XL U1018 ( .A(n673), .B(n672), .Y(mult_x_1_n224) );
  INVXL U1019 ( .A(n675), .Y(n717) );
  NOR2XL U1020 ( .A(n717), .B(n1260), .Y(n680) );
  INVXL U1021 ( .A(n678), .Y(n718) );
  OAI21XL U1022 ( .A0(n718), .A1(n1260), .B0(n1261), .Y(n679) );
  CMPR22X1 U1023 ( .A(n693), .B(n692), .CO(n701), .S(n739) );
  XNOR2X1 U1024 ( .A(n769), .B(B[21]), .Y(n731) );
  XNOR2X1 U1025 ( .A(A[15]), .B(B[7]), .Y(n732) );
  OAI22X1 U1026 ( .A0(n813), .A1(n732), .B0(n1176), .B1(n695), .Y(n729) );
  XNOR2X1 U1027 ( .A(n1091), .B(n773), .Y(n742) );
  ADDFHX1 U1028 ( .A(n708), .B(n707), .CI(n706), .CO(n700), .S(n765) );
  CMPR32X1 U1029 ( .A(n714), .B(n713), .C(n712), .CO(n687), .S(n723) );
  NOR2XL U1030 ( .A(n716), .B(n715), .Y(mult_x_1_n232) );
  NAND2XL U1031 ( .A(n716), .B(n715), .Y(mult_x_1_n233) );
  NAND2XL U1032 ( .A(n797), .B(n675), .Y(n720) );
  AOI21XL U1033 ( .A0(n798), .A1(n675), .B0(n678), .Y(n719) );
  CMPR32X1 U1034 ( .A(n728), .B(n727), .C(n726), .CO(n712), .S(n763) );
  CMPR22X1 U1035 ( .A(n730), .B(n729), .CO(n738), .S(n780) );
  OAI22X1 U1036 ( .A0(n953), .A1(n770), .B0(n731), .B1(n1077), .Y(n768) );
  XNOR2X1 U1037 ( .A(A[15]), .B(n941), .Y(n772) );
  OAI22X1 U1038 ( .A0(n1178), .A1(n772), .B0(n1176), .B1(n732), .Y(n767) );
  XNOR2X1 U1039 ( .A(n469), .B(B[18]), .Y(n776) );
  OAI22X1 U1040 ( .A0(n735), .A1(n776), .B0(n961), .B1(n734), .Y(n787) );
  XNOR2X1 U1041 ( .A(n782), .B(n740), .Y(n783) );
  XNOR2X1 U1042 ( .A(n1091), .B(B[10]), .Y(n784) );
  NAND2XL U1043 ( .A(n755), .B(n754), .Y(mult_x_1_n242) );
  INVX1 U1044 ( .A(n1264), .Y(n800) );
  CMPR32X1 U1045 ( .A(n766), .B(n765), .C(n764), .CO(n751), .S(n803) );
  CMPR22X1 U1046 ( .A(n768), .B(n767), .CO(n779), .S(n822) );
  XNOR2X1 U1047 ( .A(n769), .B(B[19]), .Y(n809) );
  XNOR2X1 U1048 ( .A(A[15]), .B(n771), .Y(n811) );
  OAI22X1 U1049 ( .A0(n1178), .A1(n811), .B0(n1176), .B1(n772), .Y(n807) );
  XNOR2X1 U1050 ( .A(n774), .B(n773), .Y(n814) );
  XNOR2X1 U1051 ( .A(n469), .B(B[17]), .Y(n816) );
  OAI22X1 U1052 ( .A0(n963), .A1(n816), .B0(n961), .B1(n776), .Y(n830) );
  XNOR2X1 U1053 ( .A(n782), .B(n781), .Y(n823) );
  OAI22XL U1054 ( .A0(n967), .A1(n823), .B0(n965), .B1(n783), .Y(n834) );
  XNOR2X1 U1055 ( .A(n1091), .B(B[9]), .Y(n825) );
  OAI22XL U1056 ( .A0(n1112), .A1(n825), .B0(n1110), .B1(n784), .Y(n833) );
  CMPR32X1 U1057 ( .A(n788), .B(n787), .C(n786), .CO(n778), .S(n852) );
  NOR2XL U1058 ( .A(n796), .B(n795), .Y(mult_x_1_n252) );
  NAND2XL U1059 ( .A(n796), .B(n795), .Y(mult_x_1_n253) );
  CMPR32X1 U1060 ( .A(n803), .B(n802), .C(n801), .CO(n795), .S(n839) );
  CMPR32X1 U1061 ( .A(n806), .B(n805), .C(n804), .CO(n792), .S(n850) );
  CMPR22X1 U1062 ( .A(n808), .B(n807), .CO(n821), .S(n861) );
  OAI22X1 U1063 ( .A0(n953), .A1(n810), .B0(n809), .B1(n1077), .Y(n855) );
  OAI22X1 U1064 ( .A0(n813), .A1(n812), .B0(n1176), .B1(n811), .Y(n854) );
  OAI22X2 U1065 ( .A0(n963), .A1(n817), .B0(n961), .B1(n816), .Y(n866) );
  OAI22XL U1066 ( .A0(n1112), .A1(n826), .B0(n1110), .B1(n825), .Y(n869) );
  CMPR32X1 U1067 ( .A(n834), .B(n833), .C(n832), .CO(n853), .S(n883) );
  NOR2XL U1068 ( .A(n839), .B(n838), .Y(mult_x_1_n259) );
  NAND2XL U1069 ( .A(n839), .B(n838), .Y(mult_x_1_n260) );
  INVXL U1070 ( .A(n840), .Y(n877) );
  NAND2XL U1071 ( .A(n840), .B(n878), .Y(n844) );
  INVXL U1072 ( .A(n1269), .Y(n842) );
  AOI21XL U1073 ( .A0(n841), .A1(n878), .B0(n842), .Y(n843) );
  INVXL U1074 ( .A(n1266), .Y(n845) );
  NAND2XL U1075 ( .A(n845), .B(n1267), .Y(n846) );
  XNOR2X1 U1076 ( .A(n847), .B(n846), .Y(PRODUCT[22]) );
  CMPR32X1 U1077 ( .A(n853), .B(n852), .C(n851), .CO(n835), .S(n882) );
  CMPR22X1 U1078 ( .A(n855), .B(n854), .CO(n860), .S(n891) );
  CMPR32X1 U1079 ( .A(n864), .B(n863), .C(n862), .CO(n907), .S(n892) );
  CMPR32X1 U1080 ( .A(n870), .B(n869), .C(n868), .CO(n885), .S(n905) );
  CMPR32X1 U1081 ( .A(n873), .B(n872), .C(n871), .CO(n849), .S(n880) );
  NOR2XL U1082 ( .A(n875), .B(n874), .Y(mult_x_1_n270) );
  NAND2XL U1083 ( .A(n875), .B(n874), .Y(mult_x_1_n271) );
  CMPR32X1 U1084 ( .A(n888), .B(n887), .C(n886), .CO(n913), .S(n909) );
  CMPR32X1 U1085 ( .A(n891), .B(n890), .C(n889), .CO(n897), .S(n912) );
  CMPR32X1 U1086 ( .A(n894), .B(n893), .C(n892), .CO(n911), .S(n923) );
  NOR2XL U1087 ( .A(n899), .B(n898), .Y(mult_x_1_n277) );
  INVXL U1088 ( .A(n1270), .Y(n900) );
  CMPR32X1 U1089 ( .A(n913), .B(n912), .C(n911), .CO(n903), .S(n918) );
  NOR2XL U1090 ( .A(n915), .B(n914), .Y(mult_x_1_n288) );
  NAND2XL U1091 ( .A(n915), .B(n914), .Y(mult_x_1_n289) );
  CMPR32X1 U1092 ( .A(n920), .B(n919), .C(n918), .CO(n914), .S(n925) );
  NOR2XL U1093 ( .A(n925), .B(n924), .Y(mult_x_1_n291) );
  NAND2XL U1094 ( .A(n925), .B(n924), .Y(mult_x_1_n292) );
  AOI21X1 U1095 ( .A0(n1005), .A1(n1279), .B0(n1286), .Y(n933) );
  OAI21XL U1096 ( .A0(n933), .A1(n1277), .B0(n1278), .Y(n928) );
  INVXL U1097 ( .A(n1275), .Y(n926) );
  XNOR2X2 U1098 ( .A(n928), .B(n927), .Y(PRODUCT[18]) );
  INVXL U1099 ( .A(n1277), .Y(n931) );
  NAND2XL U1100 ( .A(n931), .B(n1278), .Y(n932) );
  XOR2X1 U1101 ( .A(n933), .B(n932), .Y(PRODUCT[17]) );
  NAND2XL U1102 ( .A(n935), .B(n934), .Y(mult_x_1_n303) );
  INVX1 U1103 ( .A(n1281), .Y(n1003) );
  INVXL U1104 ( .A(n1282), .Y(n936) );
  AOI21X1 U1105 ( .A0(n1005), .A1(n1003), .B0(n936), .Y(n937) );
  CMPR32X1 U1106 ( .A(n940), .B(n939), .C(n938), .CO(n202), .S(n995) );
  XNOR2XL U1107 ( .A(n1129), .B(B[0]), .Y(n945) );
  XNOR2XL U1108 ( .A(n1091), .B(B[2]), .Y(n954) );
  OAI22XL U1109 ( .A0(n963), .A1(n962), .B0(n961), .B1(n960), .Y(n1016) );
  OAI22XL U1110 ( .A0(n967), .A1(n966), .B0(n965), .B1(n964), .Y(n1015) );
  CMPR32X1 U1111 ( .A(n973), .B(n972), .C(n971), .CO(n968), .S(n1039) );
  CMPR32X1 U1112 ( .A(n976), .B(n975), .C(n974), .CO(n989), .S(n1020) );
  ADDFHX1 U1113 ( .A(n979), .B(n978), .CI(n977), .CO(n972), .S(n1019) );
  CMPR22X1 U1114 ( .A(n983), .B(n982), .CO(n1022), .S(n1012) );
  ADDFHX1 U1115 ( .A(n986), .B(n985), .CI(n984), .CO(n1007), .S(n1021) );
  CMPR32X1 U1116 ( .A(n989), .B(n988), .C(n987), .CO(n994), .S(n1037) );
  CMPR32X1 U1117 ( .A(n992), .B(n991), .C(n990), .CO(n934), .S(n999) );
  NOR2XL U1118 ( .A(n1000), .B(mult_x_1_n312), .Y(mult_x_1_n305) );
  INVXL U1119 ( .A(n1000), .Y(n1002) );
  NAND2XL U1120 ( .A(n1002), .B(n1001), .Y(mult_x_1_n78) );
  XNOR2X1 U1121 ( .A(n1005), .B(n1004), .Y(PRODUCT[15]) );
  XNOR2X1 U1122 ( .A(n1288), .B(n1284), .Y(PRODUCT[14]) );
  CMPR32X1 U1123 ( .A(n1008), .B(n1007), .C(n1006), .CO(n987), .S(n1042) );
  CMPR32X1 U1124 ( .A(n1011), .B(n1010), .C(n1009), .CO(n1029), .S(n1024) );
  CMPR32X1 U1125 ( .A(n1014), .B(n1013), .C(n1012), .CO(n1028), .S(n1035) );
  CMPR32X1 U1126 ( .A(n1017), .B(n1016), .C(n1015), .CO(n1006), .S(n1027) );
  CMPR32X1 U1127 ( .A(n1020), .B(n1019), .C(n1018), .CO(n1038), .S(n1040) );
  CMPR32X1 U1128 ( .A(n1023), .B(n1022), .C(n1021), .CO(n1018), .S(n1032) );
  CMPR32X1 U1129 ( .A(n1026), .B(n1025), .C(n1024), .CO(n1031), .S(n1033) );
  CMPR32X1 U1130 ( .A(n1032), .B(n1031), .C(n1030), .CO(n1045), .S(n1044) );
  NAND2XL U1131 ( .A(n1056), .B(n1059), .Y(n1054) );
  NOR2XL U1132 ( .A(n1054), .B(n1050), .Y(mult_x_1_n316) );
  INVXL U1133 ( .A(n1057), .Y(n1060) );
  NAND2XL U1134 ( .A(n1046), .B(n1045), .Y(n1055) );
  INVXL U1135 ( .A(n1055), .Y(n1047) );
  OAI21XL U1136 ( .A0(n1053), .A1(n1050), .B0(n1051), .Y(mult_x_1_n317) );
  INVXL U1137 ( .A(n1050), .Y(n1052) );
  NAND2XL U1138 ( .A(n1052), .B(n1051), .Y(mult_x_1_n80) );
  XNOR2X1 U1139 ( .A(n1289), .B(n1285), .Y(PRODUCT[13]) );
  INVX1 U1140 ( .A(mult_x_1_n335), .Y(n1061) );
  OAI21XL U1141 ( .A0(n1061), .A1(n1054), .B0(n1053), .Y(mult_x_1_n320) );
  NAND2XL U1142 ( .A(n1056), .B(n1055), .Y(mult_x_1_n81) );
  NAND2XL U1143 ( .A(n1059), .B(n1057), .Y(n1058) );
  XOR2X1 U1144 ( .A(n1061), .B(n1058), .Y(n1304) );
  OAI21XL U1145 ( .A0(n1061), .A1(n1036), .B0(n1057), .Y(mult_x_1_n327) );
  INVXL U1146 ( .A(n1062), .Y(n1070) );
  AOI21XL U1147 ( .A0(n1070), .A1(n382), .B0(n1063), .Y(n1067) );
  NAND2XL U1148 ( .A(n382), .B(n1068), .Y(n1069) );
  INVXL U1149 ( .A(n1071), .Y(n1188) );
  OAI21XL U1150 ( .A0(n1188), .A1(n1184), .B0(n1185), .Y(n1076) );
  INVXL U1151 ( .A(n1072), .Y(n1074) );
  XNOR2X1 U1152 ( .A(A[15]), .B(B[21]), .Y(n1109) );
  CMPR32X1 U1153 ( .A(n1096), .B(n1095), .C(n1094), .CO(n1113), .S(n1085) );
  CMPR32X1 U1154 ( .A(n1099), .B(n1098), .C(n1097), .CO(n1102), .S(n1084) );
  CMPR32X1 U1155 ( .A(n1107), .B(n1106), .C(n1105), .CO(n1149), .S(n1104) );
  XNOR2X1 U1156 ( .A(A[15]), .B(B[22]), .Y(n1134) );
  OAI22X1 U1157 ( .A0(n1112), .A1(n1111), .B0(n1110), .B1(n1135), .Y(n1144) );
  CMPR32X1 U1158 ( .A(n1115), .B(n1114), .C(n1113), .CO(n1147), .S(n1103) );
  AOI21XL U1159 ( .A0(n1223), .A1(n1123), .B0(n1122), .Y(n1124) );
  CMPR32X1 U1160 ( .A(n1133), .B(n1132), .C(n1131), .CO(n1151), .S(n1148) );
  XNOR2X1 U1161 ( .A(A[15]), .B(B[23]), .Y(n1139) );
  XNOR2X1 U1162 ( .A(A[15]), .B(B[24]), .Y(n1158) );
  OAI22X1 U1163 ( .A0(n1141), .A1(n1140), .B0(n1162), .B1(n1159), .Y(n1173) );
  CMPR32X1 U1164 ( .A(n1144), .B(n1143), .C(n1142), .CO(n1155), .S(n1150) );
  CMPR32X1 U1165 ( .A(n1149), .B(n1148), .C(n1147), .CO(n1154), .S(n1116) );
  CMPR32X1 U1166 ( .A(n1152), .B(n1151), .C(n1150), .CO(n1146), .S(n1153) );
  CMPR32X1 U1167 ( .A(n1157), .B(n1156), .C(n1155), .CO(n1170), .S(n1145) );
  OAI21XL U1168 ( .A0(n1164), .A1(n1234), .B0(n1235), .Y(n1219) );
  AOI21XL U1169 ( .A0(n1223), .A1(n1215), .B0(n1219), .Y(n1165) );
  CMPR32X1 U1170 ( .A(n1173), .B(n1172), .C(n1171), .CO(n1181), .S(n1169) );
  XNOR2XL U1171 ( .A(A[15]), .B(n1174), .Y(n1175) );
  AOI21XL U1172 ( .A0(n1197), .A1(n1196), .B0(n1190), .Y(n1194) );
  AOI21XL U1173 ( .A0(n1223), .A1(n1222), .B0(n1221), .Y(n1224) );
  XNOR2XL U1174 ( .A(n1230), .B(n1229), .Y(n1311) );
endmodule


module FFT2048_DW02_mult_2_stage_J1_13 ( A, B, TC, CLK, PRODUCT );
  input [15:0] A;
  input [26:0] B;
  output [42:0] PRODUCT;
  input TC, CLK;
  wire   n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, mult_x_1_n335, mult_x_1_n327, mult_x_1_n320,
         mult_x_1_n317, mult_x_1_n316, mult_x_1_n313, mult_x_1_n312,
         mult_x_1_n306, mult_x_1_n305, mult_x_1_n303, mult_x_1_n302,
         mult_x_1_n300, mult_x_1_n299, mult_x_1_n297, mult_x_1_n292,
         mult_x_1_n291, mult_x_1_n289, mult_x_1_n288, mult_x_1_n278,
         mult_x_1_n277, mult_x_1_n271, mult_x_1_n270, mult_x_1_n260,
         mult_x_1_n259, mult_x_1_n253, mult_x_1_n252, mult_x_1_n242,
         mult_x_1_n241, mult_x_1_n233, mult_x_1_n232, mult_x_1_n224,
         mult_x_1_n223, mult_x_1_n221, mult_x_1_n220, mult_x_1_n210,
         mult_x_1_n209, mult_x_1_n203, mult_x_1_n202, mult_x_1_n192,
         mult_x_1_n191, mult_x_1_n185, mult_x_1_n184, mult_x_1_n174,
         mult_x_1_n173, mult_x_1_n163, mult_x_1_n162, mult_x_1_n150,
         mult_x_1_n149, mult_x_1_n135, mult_x_1_n134, mult_x_1_n126,
         mult_x_1_n125, mult_x_1_n115, mult_x_1_n114, mult_x_1_n106,
         mult_x_1_n105, mult_x_1_n81, mult_x_1_n80, mult_x_1_n78, mult_x_1_n54,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233;

  DFFHQXL mult_x_1_clk_r_REG20_S1 ( .D(mult_x_1_n223), .CK(CLK), .Q(n1199) );
  DFFHQXL mult_x_1_clk_r_REG22_S1 ( .D(mult_x_1_n220), .CK(CLK), .Q(n1197) );
  DFFHQXL mult_x_1_clk_r_REG19_S1 ( .D(mult_x_1_n224), .CK(CLK), .Q(n1200) );
  DFFHQXL mult_x_1_clk_r_REG40_S1 ( .D(mult_x_1_n173), .CK(CLK), .Q(n1187) );
  DFFHQXL mult_x_1_clk_r_REG24_S1 ( .D(mult_x_1_n209), .CK(CLK), .Q(n1195) );
  DFFHQX4 mult_x_1_clk_r_REG61_S1 ( .D(mult_x_1_n335), .CK(CLK), .Q(n1233) );
  DFFHQX4 mult_x_1_clk_r_REG57_S1 ( .D(mult_x_1_n320), .CK(CLK), .Q(n1231) );
  DFFHQX4 mult_x_1_clk_r_REG54_S1 ( .D(mult_x_1_n317), .CK(CLK), .Q(n1230) );
  DFFHQX4 mult_x_1_clk_r_REG1_S1 ( .D(mult_x_1_n306), .CK(CLK), .Q(n1229) );
  DFFHQX4 mult_x_1_clk_r_REG55_S1 ( .D(mult_x_1_n316), .CK(CLK), .Q(n1226) );
  DFFHQX1 mult_x_1_clk_r_REG0_S1 ( .D(mult_x_1_n313), .CK(CLK), .Q(n1225) );
  DFFHQX4 mult_x_1_clk_r_REG7_S1 ( .D(mult_x_1_n297), .CK(CLK), .Q(n1217) );
  DFFHQX4 mult_x_1_clk_r_REG10_S1 ( .D(mult_x_1_n292), .CK(CLK), .Q(n1216) );
  DFFHQX4 mult_x_1_clk_r_REG32_S1 ( .D(mult_x_1_n288), .CK(CLK), .Q(n1213) );
  DFFHQX4 mult_x_1_clk_r_REG29_S1 ( .D(mult_x_1_n278), .CK(CLK), .Q(n1212) );
  DFFHQX4 mult_x_1_clk_r_REG30_S1 ( .D(mult_x_1_n277), .CK(CLK), .Q(n1211) );
  DFFHQX4 mult_x_1_clk_r_REG28_S1 ( .D(mult_x_1_n270), .CK(CLK), .Q(n1209) );
  DFFHQX4 mult_x_1_clk_r_REG26_S1 ( .D(mult_x_1_n259), .CK(CLK), .Q(n1207) );
  DFFHQX4 mult_x_1_clk_r_REG14_S1 ( .D(mult_x_1_n252), .CK(CLK), .Q(n1205) );
  DFFHQX1 mult_x_1_clk_r_REG17_S1 ( .D(mult_x_1_n233), .CK(CLK), .Q(n1202) );
  DFFHQXL clk_r_REG58_S1 ( .D(n1247), .CK(CLK), .Q(PRODUCT[12]) );
  DFFHQXL clk_r_REG60_S1 ( .D(n1248), .CK(CLK), .Q(PRODUCT[11]) );
  DFFHQXL mult_x_1_clk_r_REG37_S1 ( .D(mult_x_1_n185), .CK(CLK), .Q(n1190) );
  DFFHQXL mult_x_1_clk_r_REG34_S1 ( .D(mult_x_1_n202), .CK(CLK), .Q(n1193) );
  DFFHQXL mult_x_1_clk_r_REG4_S1 ( .D(mult_x_1_n78), .CK(CLK), .Q(n1223) );
  DFFHQXL mult_x_1_clk_r_REG36_S1 ( .D(mult_x_1_n191), .CK(CLK), .Q(n1191) );
  DFFHQXL mult_x_1_clk_r_REG44_S1 ( .D(mult_x_1_n149), .CK(CLK), .Q(n1183) );
  DFFHQXL clk_r_REG62_S1 ( .D(n1249), .CK(CLK), .Q(PRODUCT[10]) );
  DFFHQXL clk_r_REG63_S1 ( .D(n1250), .CK(CLK), .Q(PRODUCT[9]) );
  DFFHQXL mult_x_1_clk_r_REG23_S1 ( .D(mult_x_1_n210), .CK(CLK), .Q(n1196) );
  DFFHQXL mult_x_1_clk_r_REG42_S1 ( .D(mult_x_1_n162), .CK(CLK), .Q(n1185) );
  DFFHQXL mult_x_1_clk_r_REG41_S1 ( .D(mult_x_1_n163), .CK(CLK), .Q(n1186) );
  DFFHQXL mult_x_1_clk_r_REG35_S1 ( .D(mult_x_1_n192), .CK(CLK), .Q(n1192) );
  DFFHQXL mult_x_1_clk_r_REG33_S1 ( .D(mult_x_1_n203), .CK(CLK), .Q(n1194) );
  DFFHQXL clk_r_REG68_S1 ( .D(n1255), .CK(CLK), .Q(PRODUCT[4]) );
  DFFHQXL mult_x_1_clk_r_REG49_S1 ( .D(mult_x_1_n115), .CK(CLK), .Q(n1178) );
  DFFHQXL mult_x_1_clk_r_REG39_S1 ( .D(mult_x_1_n174), .CK(CLK), .Q(n1188) );
  DFFHQXL clk_r_REG64_S1 ( .D(n1251), .CK(CLK), .Q(PRODUCT[8]) );
  DFFHQXL clk_r_REG72_S1 ( .D(n1259), .CK(CLK), .Q(PRODUCT[0]) );
  DFFHQXL clk_r_REG65_S1 ( .D(n1252), .CK(CLK), .Q(PRODUCT[7]) );
  DFFHQXL clk_r_REG66_S1 ( .D(n1253), .CK(CLK), .Q(PRODUCT[6]) );
  DFFHQXL clk_r_REG67_S1 ( .D(n1254), .CK(CLK), .Q(PRODUCT[5]) );
  DFFHQXL clk_r_REG69_S1 ( .D(n1256), .CK(CLK), .Q(PRODUCT[3]) );
  DFFHQXL clk_r_REG70_S1 ( .D(n1257), .CK(CLK), .Q(PRODUCT[2]) );
  DFFHQXL clk_r_REG71_S1 ( .D(n1258), .CK(CLK), .Q(PRODUCT[1]) );
  DFFHQX1 mult_x_1_clk_r_REG2_S1 ( .D(mult_x_1_n312), .CK(CLK), .Q(n1224) );
  DFFHQXL mult_x_1_clk_r_REG59_S1 ( .D(mult_x_1_n327), .CK(CLK), .Q(n1232) );
  DFFHQXL mult_x_1_clk_r_REG56_S1 ( .D(mult_x_1_n81), .CK(CLK), .Q(n1228) );
  DFFHQX1 mult_x_1_clk_r_REG53_S1 ( .D(mult_x_1_n80), .CK(CLK), .Q(n1227) );
  DFFHQXL mult_x_1_clk_r_REG6_S1 ( .D(mult_x_1_n302), .CK(CLK), .Q(n1220) );
  DFFHQXL mult_x_1_clk_r_REG21_S1 ( .D(mult_x_1_n221), .CK(CLK), .Q(n1198) );
  DFFHQXL mult_x_1_clk_r_REG38_S1 ( .D(mult_x_1_n184), .CK(CLK), .Q(n1189) );
  DFFHQXL mult_x_1_clk_r_REG43_S1 ( .D(mult_x_1_n150), .CK(CLK), .Q(n1184) );
  DFFHQXL mult_x_1_clk_r_REG45_S1 ( .D(mult_x_1_n135), .CK(CLK), .Q(n1182) );
  DFFHQXL mult_x_1_clk_r_REG46_S1 ( .D(mult_x_1_n134), .CK(CLK), .Q(n1181) );
  DFFHQXL mult_x_1_clk_r_REG47_S1 ( .D(mult_x_1_n126), .CK(CLK), .Q(n1180) );
  DFFHQXL mult_x_1_clk_r_REG48_S1 ( .D(mult_x_1_n125), .CK(CLK), .Q(n1179) );
  DFFHQXL mult_x_1_clk_r_REG50_S1 ( .D(mult_x_1_n114), .CK(CLK), .Q(n1177) );
  DFFHQXL mult_x_1_clk_r_REG51_S1 ( .D(mult_x_1_n106), .CK(CLK), .Q(n1176) );
  DFFHQXL mult_x_1_clk_r_REG52_S1 ( .D(mult_x_1_n105), .CK(CLK), .Q(n1175) );
  DFFHQXL mult_x_1_clk_r_REG12_S1 ( .D(mult_x_1_n54), .CK(CLK), .Q(n1174) );
  DFFHQX2 mult_x_1_clk_r_REG27_S1 ( .D(mult_x_1_n271), .CK(CLK), .Q(n1210) );
  DFFHQX1 mult_x_1_clk_r_REG15_S1 ( .D(mult_x_1_n242), .CK(CLK), .Q(n1204) );
  DFFHQX2 mult_x_1_clk_r_REG25_S1 ( .D(mult_x_1_n260), .CK(CLK), .Q(n1208) );
  DFFHQX2 mult_x_1_clk_r_REG31_S1 ( .D(mult_x_1_n289), .CK(CLK), .Q(n1214) );
  DFFHQX1 mult_x_1_clk_r_REG11_S1 ( .D(mult_x_1_n291), .CK(CLK), .Q(n1215) );
  DFFHQX1 mult_x_1_clk_r_REG9_S1 ( .D(mult_x_1_n299), .CK(CLK), .Q(n1218) );
  DFFHQX1 mult_x_1_clk_r_REG8_S1 ( .D(mult_x_1_n300), .CK(CLK), .Q(n1219) );
  DFFHQX2 mult_x_1_clk_r_REG5_S1 ( .D(mult_x_1_n303), .CK(CLK), .Q(n1221) );
  DFFHQX2 mult_x_1_clk_r_REG16_S1 ( .D(mult_x_1_n241), .CK(CLK), .Q(n1203) );
  DFFHQX2 mult_x_1_clk_r_REG13_S1 ( .D(mult_x_1_n253), .CK(CLK), .Q(n1206) );
  DFFHQX2 mult_x_1_clk_r_REG18_S1 ( .D(mult_x_1_n232), .CK(CLK), .Q(n1201) );
  DFFHQX1 mult_x_1_clk_r_REG3_S1 ( .D(mult_x_1_n305), .CK(CLK), .Q(n1222) );
  CMPR32X1 U1 ( .A(n1025), .B(n1024), .C(n1023), .CO(n1040), .S(n398) );
  ADDFHX1 U2 ( .A(n514), .B(n513), .CI(n512), .CO(n501), .S(n542) );
  ADDFHX1 U3 ( .A(n476), .B(n475), .CI(n474), .CO(n469), .S(n502) );
  ADDFHX2 U4 ( .A(n500), .B(n499), .CI(n498), .CO(n475), .S(n512) );
  ADDFHX1 U5 ( .A(n576), .B(n575), .CI(n574), .CO(n549), .S(n582) );
  ADDFHX1 U6 ( .A(n540), .B(n539), .CI(n538), .CO(n513), .S(n548) );
  ADDFHX1 U7 ( .A(n904), .B(n903), .CI(n902), .CO(n905), .S(n917) );
  ADDFHX2 U8 ( .A(n752), .B(n751), .CI(n750), .CO(n767), .S(n815) );
  CMPR32X1 U9 ( .A(n966), .B(n965), .C(n964), .CO(n925), .S(n976) );
  ADDFHX1 U10 ( .A(n270), .B(n269), .CI(n268), .CO(n903), .S(n910) );
  ADDFHX1 U11 ( .A(n609), .B(n608), .CI(n607), .CO(n583), .S(n614) );
  ADDFX2 U12 ( .A(n764), .B(n763), .CI(n762), .CO(n779), .S(n830) );
  ADDFHX1 U13 ( .A(n325), .B(n324), .CI(n323), .CO(n336), .S(n964) );
  ADDFHX1 U14 ( .A(n842), .B(n841), .CI(n840), .CO(n854), .S(n878) );
  CMPR32X1 U15 ( .A(n797), .B(n796), .C(n795), .CO(n816), .S(n853) );
  ADDFX2 U16 ( .A(n570), .B(n569), .CI(n568), .CO(n562), .S(n618) );
  ADDFX2 U17 ( .A(n603), .B(n602), .CI(n601), .CO(n595), .S(n659) );
  ADDFX2 U18 ( .A(n712), .B(n711), .CI(n710), .CO(n725), .S(n766) );
  ADDFX2 U19 ( .A(n719), .B(n718), .CI(n717), .CO(n710), .S(n778) );
  BUFX3 U20 ( .A(A[11]), .Y(n1049) );
  BUFX3 U21 ( .A(A[3]), .Y(n437) );
  BUFX3 U22 ( .A(A[1]), .Y(n485) );
  XNOR2X1 U23 ( .A(n24), .B(n1157), .Y(PRODUCT[36]) );
  OAI21X1 U24 ( .A0(n1018), .A1(n1017), .B0(n1016), .Y(n1169) );
  OAI21XL U25 ( .A0(n432), .A1(n1172), .B0(n23), .Y(n435) );
  XOR2X1 U26 ( .A(n1172), .B(n613), .Y(PRODUCT[27]) );
  XNOR2X1 U27 ( .A(n654), .B(n653), .Y(PRODUCT[26]) );
  XNOR2X1 U28 ( .A(n733), .B(n732), .Y(PRODUCT[24]) );
  XNOR2X1 U29 ( .A(n826), .B(n825), .Y(PRODUCT[22]) );
  XNOR2X2 U30 ( .A(n861), .B(n860), .Y(PRODUCT[21]) );
  XOR2X1 U31 ( .A(n920), .B(n919), .Y(PRODUCT[17]) );
  NAND2X2 U32 ( .A(n16), .B(n15), .Y(n932) );
  NOR2X1 U33 ( .A(n1209), .B(n1211), .Y(n340) );
  OAI21XL U34 ( .A0(n1209), .A1(n1212), .B0(n1210), .Y(n30) );
  CLKINVX2 U35 ( .A(n1230), .Y(n15) );
  OAI21XL U36 ( .A0(n1172), .A1(n1006), .B0(n1018), .Y(n473) );
  XNOR2XL U37 ( .A(n1022), .B(n1021), .Y(PRODUCT[37]) );
  XOR2X2 U38 ( .A(n581), .B(n580), .Y(PRODUCT[28]) );
  XNOR2X1 U39 ( .A(n909), .B(n908), .Y(PRODUCT[18]) );
  XNOR2XL U40 ( .A(n757), .B(n708), .Y(n264) );
  XNOR2XL U41 ( .A(n1049), .B(n257), .Y(n277) );
  XNOR2XL U42 ( .A(n1067), .B(B[18]), .Y(n411) );
  XNOR2XL U43 ( .A(n1114), .B(B[14]), .Y(n454) );
  XNOR2XL U44 ( .A(n1096), .B(B[20]), .Y(n1026) );
  ADDFX2 U45 ( .A(n695), .B(n694), .CI(n693), .CO(n684), .S(n727) );
  XNOR2XL U46 ( .A(n1138), .B(n1137), .Y(n1253) );
  XNOR2XL U47 ( .A(n993), .B(n992), .Y(n1249) );
  OAI21XL U48 ( .A0(n986), .A1(n197), .B0(n196), .Y(mult_x_1_n335) );
  OR2X2 U49 ( .A(n192), .B(n191), .Y(n5) );
  NOR2X1 U50 ( .A(n502), .B(n501), .Y(mult_x_1_n191) );
  XOR2X1 U51 ( .A(n1134), .B(n1133), .Y(n1252) );
  NAND2X1 U52 ( .A(n971), .B(n970), .Y(n981) );
  XNOR2X1 U53 ( .A(n521), .B(n520), .Y(n563) );
  OR2X1 U54 ( .A(n521), .B(n520), .Y(n527) );
  ADDFHX1 U55 ( .A(n810), .B(n809), .CI(n808), .CO(n795), .S(n866) );
  XNOR2X1 U56 ( .A(n1096), .B(n753), .Y(n436) );
  XNOR2X1 U57 ( .A(n757), .B(n753), .Y(n715) );
  XNOR2X1 U58 ( .A(n485), .B(n1113), .Y(n518) );
  OAI2BB1X1 U59 ( .A0N(n1007), .A1N(n25), .B0(n1155), .Y(n24) );
  XNOR2X1 U60 ( .A(n1114), .B(n257), .Y(n228) );
  XNOR2X1 U61 ( .A(n485), .B(n257), .Y(n125) );
  INVXL U62 ( .A(n1172), .Y(n25) );
  BUFX3 U63 ( .A(B[3]), .Y(n257) );
  INVX1 U64 ( .A(n1018), .Y(n470) );
  NOR2XL U65 ( .A(n1012), .B(n1187), .Y(n1014) );
  OAI21X1 U66 ( .A0(n1208), .A1(n1205), .B0(n1206), .Y(n647) );
  INVXL U67 ( .A(n1205), .Y(n731) );
  INVX1 U68 ( .A(n1191), .Y(n471) );
  XNOR2X1 U69 ( .A(A[8]), .B(A[7]), .Y(n62) );
  XNOR2X1 U70 ( .A(n999), .B(n998), .Y(n1250) );
  XOR2X1 U71 ( .A(n1128), .B(n1127), .Y(n1251) );
  INVX1 U72 ( .A(n986), .Y(n993) );
  NAND2X1 U73 ( .A(n50), .B(n49), .Y(n610) );
  NAND2X1 U74 ( .A(n976), .B(n975), .Y(n1002) );
  INVXL U75 ( .A(n972), .Y(n53) );
  NOR2X1 U76 ( .A(n971), .B(n970), .Y(n963) );
  XNOR2X1 U77 ( .A(n724), .B(n34), .Y(n33) );
  INVX1 U78 ( .A(n104), .Y(n1132) );
  INVX1 U79 ( .A(n991), .Y(n987) );
  NOR2X1 U80 ( .A(n149), .B(n148), .Y(n1124) );
  ADDFHX1 U81 ( .A(n867), .B(n866), .CI(n865), .CO(n852), .S(n887) );
  NAND2X1 U82 ( .A(n149), .B(n148), .Y(n1125) );
  NOR2X1 U83 ( .A(n151), .B(n150), .Y(n995) );
  OAI22X1 U84 ( .A0(n259), .A1(n791), .B0(n792), .B1(n22), .Y(n304) );
  XNOR2X1 U85 ( .A(n365), .B(n1113), .Y(n366) );
  BUFX3 U86 ( .A(B[15]), .Y(n753) );
  NAND2X1 U87 ( .A(n1005), .B(n1014), .Y(n1017) );
  INVX1 U88 ( .A(n1006), .Y(n430) );
  NAND2X1 U89 ( .A(n690), .B(n1204), .Y(n691) );
  INVX2 U90 ( .A(n646), .Y(n6) );
  NAND2X1 U91 ( .A(n652), .B(n1202), .Y(n653) );
  NAND2X1 U92 ( .A(n907), .B(n1219), .Y(n908) );
  NAND2X1 U93 ( .A(n824), .B(n1210), .Y(n825) );
  INVX1 U94 ( .A(n819), .Y(n858) );
  NAND2X1 U95 ( .A(n1156), .B(n1182), .Y(n1157) );
  NAND2X1 U96 ( .A(n433), .B(n1190), .Y(n434) );
  NAND2X1 U97 ( .A(n404), .B(n1188), .Y(n405) );
  NAND2X1 U98 ( .A(n471), .B(n1192), .Y(n472) );
  XOR2X1 U99 ( .A(A[10]), .B(A[11]), .Y(n154) );
  BUFX3 U100 ( .A(A[5]), .Y(n365) );
  NAND2X1 U101 ( .A(n1229), .B(n1217), .Y(n13) );
  NOR2X1 U102 ( .A(n1191), .B(n1189), .Y(n1005) );
  INVX1 U103 ( .A(n1179), .Y(n1058) );
  INVXL U104 ( .A(n1224), .Y(n930) );
  OAI21XL U105 ( .A0(n1204), .A1(n1201), .B0(n1202), .Y(n17) );
  AOI21X1 U106 ( .A0(n980), .A1(n984), .B0(n974), .Y(n977) );
  NAND2XL U107 ( .A(n727), .B(n726), .Y(mult_x_1_n242) );
  NAND2BX2 U108 ( .AN(n973), .B(n53), .Y(n980) );
  NOR2X1 U109 ( .A(n976), .B(n975), .Y(n1001) );
  NOR2X1 U110 ( .A(n922), .B(n921), .Y(mult_x_1_n302) );
  NAND2XL U111 ( .A(n615), .B(n616), .Y(n49) );
  NOR2X1 U112 ( .A(n926), .B(n925), .Y(mult_x_1_n312) );
  NAND2XL U113 ( .A(n863), .B(n864), .Y(n38) );
  XOR2X1 U114 ( .A(n723), .B(n33), .Y(n734) );
  NAND2BXL U115 ( .AN(n892), .B(n57), .Y(n56) );
  NAND2XL U116 ( .A(n892), .B(n893), .Y(n55) );
  ADDFHX2 U117 ( .A(n334), .B(n333), .CI(n332), .CO(n911), .S(n913) );
  OR2XL U118 ( .A(n1121), .B(n1120), .Y(n1123) );
  ADDFHX2 U119 ( .A(n816), .B(n815), .CI(n814), .CO(n775), .S(n827) );
  NAND2BXL U120 ( .AN(n724), .B(n34), .Y(n32) );
  NAND2XL U121 ( .A(n724), .B(n725), .Y(n31) );
  ADDFHX2 U122 ( .A(n767), .B(n766), .CI(n765), .CO(n735), .S(n774) );
  INVXL U123 ( .A(n893), .Y(n57) );
  NAND2XL U124 ( .A(n184), .B(n182), .Y(n47) );
  OR2XL U125 ( .A(n494), .B(n44), .Y(n42) );
  ADDFHX2 U126 ( .A(n181), .B(n180), .CI(n179), .CO(n186), .S(n188) );
  INVXL U127 ( .A(n956), .Y(n52) );
  OR2X2 U128 ( .A(n122), .B(n121), .Y(n120) );
  ADDFHX1 U129 ( .A(n178), .B(n177), .CI(n176), .CO(n952), .S(n187) );
  OAI22XL U130 ( .A0(n807), .A1(n223), .B0(n805), .B1(n222), .Y(n236) );
  XNOR2X1 U131 ( .A(n1066), .B(n1065), .Y(PRODUCT[38]) );
  XNOR2X1 U132 ( .A(n1109), .B(n1108), .Y(PRODUCT[39]) );
  OR2XL U133 ( .A(n1152), .B(n1151), .Y(n1154) );
  NAND2BXL U134 ( .AN(n823), .B(n35), .Y(n29) );
  AND2XL U135 ( .A(n1162), .B(n1164), .Y(n1168) );
  NOR2X1 U136 ( .A(n18), .B(n17), .Y(n342) );
  NAND2X1 U137 ( .A(n61), .B(n62), .Y(n666) );
  BUFX3 U138 ( .A(n485), .Y(n205) );
  INVX2 U139 ( .A(n362), .Y(n1096) );
  AND2X2 U140 ( .A(n579), .B(n1198), .Y(n580) );
  NAND2X1 U141 ( .A(n345), .B(n503), .Y(n1006) );
  INVX1 U142 ( .A(n365), .Y(n364) );
  NAND2X1 U143 ( .A(n64), .B(n65), .Y(n303) );
  NAND2X1 U144 ( .A(n154), .B(n155), .Y(n1075) );
  NAND2X1 U145 ( .A(n13), .B(n1219), .Y(n12) );
  AND2X2 U146 ( .A(n341), .B(n647), .Y(n18) );
  NAND2X1 U147 ( .A(n198), .B(n199), .Y(n1100) );
  INVXL U148 ( .A(n1183), .Y(n1010) );
  INVX1 U149 ( .A(n1181), .Y(n1156) );
  XNOR2X1 U150 ( .A(A[10]), .B(A[9]), .Y(n155) );
  XNOR2X1 U151 ( .A(A[12]), .B(A[11]), .Y(n199) );
  INVXL U152 ( .A(n437), .Y(n7) );
  INVX1 U153 ( .A(A[15]), .Y(n362) );
  INVX1 U154 ( .A(A[0]), .Y(n68) );
  NAND2X2 U155 ( .A(n1233), .B(n1226), .Y(n16) );
  INVX1 U156 ( .A(n1211), .Y(n821) );
  INVXL U157 ( .A(n1213), .Y(n882) );
  INVX1 U158 ( .A(n1207), .Y(n771) );
  NOR2X1 U159 ( .A(n1203), .B(n1201), .Y(n341) );
  OAI22X1 U160 ( .A0(n1029), .A1(n232), .B0(n1030), .B1(n231), .Y(n241) );
  NAND2X1 U161 ( .A(n339), .B(n338), .Y(n928) );
  XNOR2X1 U162 ( .A(n757), .B(B[23]), .Y(n448) );
  XNOR2X1 U163 ( .A(B[19]), .B(n1049), .Y(n450) );
  OAI2BB1X2 U164 ( .A0N(n954), .A1N(n8), .B0(n51), .Y(n968) );
  NAND2BX1 U165 ( .AN(n955), .B(n52), .Y(n8) );
  OAI22X1 U166 ( .A0(n159), .A1(n784), .B0(n1000), .B1(n9), .Y(n319) );
  OAI22X1 U167 ( .A0(n283), .A1(n1000), .B0(n784), .B1(n9), .Y(n321) );
  XNOR2X1 U168 ( .A(n745), .B(n485), .Y(n9) );
  NAND2X4 U169 ( .A(n14), .B(n10), .Y(n35) );
  NOR2X2 U170 ( .A(n12), .B(n11), .Y(n10) );
  NOR2X1 U171 ( .A(n1218), .B(n1221), .Y(n11) );
  NAND3X2 U172 ( .A(n932), .B(n1217), .C(n1222), .Y(n14) );
  NOR2X2 U173 ( .A(n28), .B(n344), .Y(n1018) );
  NOR2X4 U174 ( .A(n20), .B(n19), .Y(n1172) );
  NOR3BX4 U175 ( .AN(n35), .B(n343), .C(n645), .Y(n19) );
  NAND2X2 U176 ( .A(n21), .B(n342), .Y(n20) );
  NAND2BX2 U177 ( .AN(n343), .B(n6), .Y(n21) );
  XNOR2X2 U178 ( .A(B[24]), .B(n757), .Y(n409) );
  NOR2X2 U179 ( .A(n339), .B(n338), .Y(n927) );
  OAI22X1 U180 ( .A0(n300), .A1(n792), .B0(n791), .B1(n22), .Y(n314) );
  XNOR2X4 U181 ( .A(n745), .B(n437), .Y(n22) );
  NOR2X1 U182 ( .A(n1195), .B(n1193), .Y(n345) );
  AOI21X1 U183 ( .A0(n470), .A1(n471), .B0(n431), .Y(n23) );
  NOR2X1 U184 ( .A(n1197), .B(n1199), .Y(n503) );
  INVXL U185 ( .A(n1185), .Y(n1004) );
  OR2X2 U186 ( .A(n1183), .B(n1185), .Y(n1012) );
  NOR2X1 U187 ( .A(n1017), .B(n1006), .Y(n1007) );
  CLKINVX3 U188 ( .A(n35), .Y(n26) );
  NAND2BX1 U189 ( .AN(n1215), .B(n1216), .Y(n27) );
  XOR2X2 U190 ( .A(n26), .B(n27), .Y(PRODUCT[19]) );
  OAI22X1 U191 ( .A0(n1076), .A1(n408), .B0(n450), .B1(n1075), .Y(n445) );
  XNOR2X1 U192 ( .A(B[20]), .B(n1049), .Y(n408) );
  XNOR2X2 U193 ( .A(B[17]), .B(n205), .Y(n227) );
  AND2X2 U194 ( .A(n504), .B(n345), .Y(n28) );
  NAND2X1 U195 ( .A(n29), .B(n822), .Y(n826) );
  AOI21X2 U196 ( .A0(n819), .A1(n340), .B0(n30), .Y(n646) );
  OAI21X2 U197 ( .A0(n1213), .A1(n1216), .B0(n1214), .Y(n819) );
  OAI2BB1X2 U198 ( .A0N(n32), .A1N(n723), .B0(n31), .Y(n694) );
  INVX1 U199 ( .A(n725), .Y(n34) );
  OAI21X1 U200 ( .A0(n1172), .A1(n544), .B0(n505), .Y(n547) );
  NOR2X1 U201 ( .A(n1207), .B(n1205), .Y(n644) );
  NAND2X2 U202 ( .A(n857), .B(n340), .Y(n645) );
  NOR2X2 U203 ( .A(n1215), .B(n1213), .Y(n857) );
  XNOR2X1 U204 ( .A(n746), .B(B[17]), .Y(n559) );
  OAI22X1 U205 ( .A0(n1118), .A1(n519), .B0(n1116), .B1(n484), .Y(n533) );
  XNOR2X1 U206 ( .A(n1114), .B(n756), .Y(n484) );
  OAI21X1 U207 ( .A0(n1172), .A1(n1199), .B0(n1200), .Y(n581) );
  OAI22X1 U208 ( .A0(n801), .A1(n672), .B0(n799), .B1(n630), .Y(n680) );
  XNOR2X1 U209 ( .A(n365), .B(B[18]), .Y(n672) );
  OAI22X1 U210 ( .A0(n1051), .A1(n755), .B0(n1076), .B1(n714), .Y(n763) );
  ADDFX2 U211 ( .A(n528), .B(n527), .CI(n526), .CO(n540), .S(n575) );
  OAI22X1 U212 ( .A0(n1029), .A1(n522), .B0(n1030), .B1(n483), .Y(n534) );
  OAI22X1 U213 ( .A0(n807), .A1(n448), .B0(n805), .B1(n409), .Y(n444) );
  OAI22X1 U214 ( .A0(n801), .A1(n754), .B0(n799), .B1(n713), .Y(n764) );
  XNOR2X1 U215 ( .A(n365), .B(B[17]), .Y(n713) );
  XNOR2X1 U216 ( .A(n354), .B(n353), .Y(PRODUCT[35]) );
  NAND2XL U217 ( .A(n1010), .B(n1184), .Y(n353) );
  XNOR2X1 U218 ( .A(n437), .B(B[23]), .Y(n560) );
  NAND2XL U219 ( .A(n1164), .B(n1176), .Y(n1108) );
  NAND2XL U220 ( .A(n1007), .B(n1162), .Y(n1107) );
  INVXL U221 ( .A(n1104), .Y(n1061) );
  XNOR2XL U222 ( .A(n757), .B(n756), .Y(n804) );
  XNOR2X1 U223 ( .A(n365), .B(B[14]), .Y(n800) );
  XNOR2XL U224 ( .A(n757), .B(n704), .Y(n806) );
  XNOR2XL U225 ( .A(n365), .B(n708), .Y(n302) );
  INVXL U226 ( .A(n1049), .Y(n361) );
  XNOR2XL U227 ( .A(n757), .B(n702), .Y(n286) );
  XNOR2XL U228 ( .A(n757), .B(n1113), .Y(n371) );
  XNOR2XL U229 ( .A(n746), .B(B[25]), .Y(n387) );
  XNOR2X1 U230 ( .A(n746), .B(B[24]), .Y(n375) );
  XNOR2XL U231 ( .A(n1067), .B(B[20]), .Y(n373) );
  XNOR2X1 U232 ( .A(n1067), .B(B[14]), .Y(n525) );
  XNOR2XL U233 ( .A(A[13]), .B(n756), .Y(n561) );
  XNOR2XL U234 ( .A(n1049), .B(B[23]), .Y(n388) );
  XNOR2XL U235 ( .A(n1067), .B(B[22]), .Y(n1032) );
  XNOR2XL U236 ( .A(n1049), .B(B[25]), .Y(n1050) );
  XNOR2XL U237 ( .A(n1067), .B(B[23]), .Y(n1047) );
  XNOR2XL U238 ( .A(n746), .B(n1113), .Y(n1027) );
  XNOR2XL U239 ( .A(n1096), .B(B[21]), .Y(n1048) );
  XNOR2XL U240 ( .A(n1096), .B(B[17]), .Y(n363) );
  XNOR2XL U241 ( .A(n1096), .B(B[18]), .Y(n370) );
  XNOR2XL U242 ( .A(n1049), .B(B[22]), .Y(n374) );
  OAI22XL U243 ( .A0(n801), .A1(n364), .B0(n799), .B1(n100), .Y(n111) );
  NAND2BXL U244 ( .AN(B[0]), .B(n365), .Y(n100) );
  XNOR2XL U245 ( .A(n437), .B(n257), .Y(n108) );
  NOR2BXL U246 ( .AN(B[0]), .B(n805), .Y(n103) );
  OAI22XL U247 ( .A0(n801), .A1(n109), .B0(n799), .B1(n94), .Y(n101) );
  XNOR2XL U248 ( .A(A[13]), .B(n1113), .Y(n1098) );
  XNOR2XL U249 ( .A(n1096), .B(B[25]), .Y(n1117) );
  XNOR2X1 U250 ( .A(n1096), .B(B[24]), .Y(n1097) );
  XNOR2XL U251 ( .A(n1096), .B(B[23]), .Y(n1077) );
  XNOR2XL U252 ( .A(n1067), .B(B[25]), .Y(n1078) );
  XNOR2X1 U253 ( .A(n1067), .B(B[24]), .Y(n1068) );
  XNOR2XL U254 ( .A(n1114), .B(B[7]), .Y(n703) );
  XNOR2XL U255 ( .A(n1114), .B(n708), .Y(n664) );
  NAND2XL U256 ( .A(n1004), .B(n1186), .Y(n359) );
  INVXL U257 ( .A(n1189), .Y(n433) );
  INVXL U258 ( .A(n1105), .Y(n1060) );
  NAND2XL U259 ( .A(n1007), .B(n1061), .Y(n1063) );
  NAND2XL U260 ( .A(n1058), .B(n1180), .Y(n1021) );
  NAND2XL U261 ( .A(n1007), .B(n1156), .Y(n1020) );
  OAI21X1 U262 ( .A0(n1172), .A1(n508), .B0(n507), .Y(n511) );
  INVXL U263 ( .A(n1193), .Y(n509) );
  INVXL U264 ( .A(n1203), .Y(n690) );
  XNOR2X1 U265 ( .A(n773), .B(n772), .Y(PRODUCT[23]) );
  NAND2XL U266 ( .A(n771), .B(n1208), .Y(n772) );
  OAI21XL U267 ( .A0(n26), .A1(n645), .B0(n646), .Y(n773) );
  AOI21XL U268 ( .A0(n932), .A1(n930), .B0(n923), .Y(n924) );
  XNOR2XL U269 ( .A(n746), .B(B[16]), .Y(n592) );
  XNOR2XL U270 ( .A(A[13]), .B(n704), .Y(n594) );
  XNOR2XL U271 ( .A(A[13]), .B(n745), .Y(n626) );
  XNOR2XL U272 ( .A(n757), .B(B[17]), .Y(n632) );
  XNOR2X1 U273 ( .A(n746), .B(B[14]), .Y(n665) );
  XNOR2X1 U274 ( .A(n1049), .B(n743), .Y(n221) );
  XNOR2XL U275 ( .A(n757), .B(B[9]), .Y(n223) );
  XNOR2XL U276 ( .A(n1067), .B(B[2]), .Y(n252) );
  XNOR2XL U277 ( .A(n365), .B(B[10]), .Y(n263) );
  NAND2BXL U278 ( .AN(B[0]), .B(A[13]), .Y(n266) );
  XNOR2XL U279 ( .A(n365), .B(B[9]), .Y(n301) );
  XNOR2XL U280 ( .A(n757), .B(B[7]), .Y(n274) );
  XNOR2XL U281 ( .A(n437), .B(n1113), .Y(n438) );
  XNOR2XL U282 ( .A(n1067), .B(B[17]), .Y(n447) );
  XNOR2XL U283 ( .A(n746), .B(B[21]), .Y(n449) );
  XNOR2X1 U284 ( .A(n1067), .B(B[19]), .Y(n377) );
  OAI22X1 U285 ( .A0(n792), .A1(n490), .B0(n791), .B1(n438), .Y(n457) );
  XNOR2XL U286 ( .A(n746), .B(B[20]), .Y(n455) );
  XNOR2XL U287 ( .A(n1067), .B(B[16]), .Y(n480) );
  XNOR2X1 U288 ( .A(n1049), .B(B[14]), .Y(n599) );
  XNOR2XL U289 ( .A(n757), .B(B[18]), .Y(n600) );
  XNOR2XL U290 ( .A(n1049), .B(B[16]), .Y(n530) );
  XNOR2XL U291 ( .A(n757), .B(B[19]), .Y(n567) );
  XNOR2XL U292 ( .A(n485), .B(B[6]), .Y(n93) );
  NAND2BXL U293 ( .AN(B[0]), .B(n757), .Y(n69) );
  NOR2XL U294 ( .A(n1104), .B(n1177), .Y(n1162) );
  INVXL U295 ( .A(n1175), .Y(n1164) );
  XNOR2X1 U296 ( .A(n1049), .B(B[24]), .Y(n1031) );
  OAI22XL U297 ( .A0(n807), .A1(n804), .B0(n805), .B1(n758), .Y(n811) );
  OAI22XL U298 ( .A0(n807), .A1(n201), .B0(n805), .B1(n806), .Y(n843) );
  OAI22X1 U299 ( .A0(n800), .A1(n799), .B0(n46), .B1(n801), .Y(n845) );
  OAI22XL U300 ( .A0(n1079), .A1(n235), .B0(n1101), .B1(n234), .Y(n239) );
  OAI22X1 U301 ( .A0(n791), .A1(n54), .B0(n233), .B1(n792), .Y(n240) );
  OAI22XL U302 ( .A0(n807), .A1(n222), .B0(n805), .B1(n201), .Y(n242) );
  OAI22XL U303 ( .A0(n1051), .A1(n220), .B0(n1076), .B1(n200), .Y(n243) );
  OAI22X1 U304 ( .A0(n219), .A1(n801), .B0(n799), .B1(n46), .Y(n244) );
  OAI22XL U305 ( .A0(n1079), .A1(n214), .B0(n1101), .B1(n235), .Y(n216) );
  OAI22XL U306 ( .A0(n1051), .A1(n174), .B0(n1076), .B1(n285), .Y(n937) );
  OAI22XL U307 ( .A0(n807), .A1(n287), .B0(n805), .B1(n286), .Y(n944) );
  INVXL U308 ( .A(n746), .Y(n368) );
  OAI22X1 U309 ( .A0(n1029), .A1(n63), .B0(n1030), .B1(n162), .Y(n164) );
  OAI22XL U310 ( .A0(n801), .A1(n67), .B0(n799), .B1(n171), .Y(n163) );
  NOR2BXL U311 ( .AN(B[0]), .B(n1076), .Y(n168) );
  OAI22XL U312 ( .A0(n666), .A1(n162), .B0(n1030), .B1(n161), .Y(n166) );
  OAI22XL U313 ( .A0(n1029), .A1(n317), .B0(n1030), .B1(n316), .Y(n950) );
  XNOR2XL U314 ( .A(n746), .B(B[22]), .Y(n412) );
  XNOR2XL U315 ( .A(n746), .B(B[23]), .Y(n407) );
  XNOR2XL U316 ( .A(n1049), .B(B[21]), .Y(n378) );
  OAI2BB1XL U317 ( .A0N(n799), .A1N(n801), .B0(n367), .Y(n416) );
  OAI22XL U318 ( .A0(n1118), .A1(n410), .B0(n1116), .B1(n363), .Y(n418) );
  INVXL U319 ( .A(n366), .Y(n367) );
  OAI2BB1XL U320 ( .A0N(n805), .A1N(n716), .B0(n372), .Y(n389) );
  OAI22XL U321 ( .A0(n1118), .A1(n370), .B0(n1116), .B1(n386), .Y(n391) );
  INVXL U322 ( .A(n371), .Y(n372) );
  OAI22XL U323 ( .A0(n1029), .A1(n375), .B0(n1030), .B1(n387), .Y(n392) );
  OAI22XL U324 ( .A0(n1079), .A1(n373), .B0(n1101), .B1(n385), .Y(n394) );
  OAI22XL U325 ( .A0(n1075), .A1(n374), .B0(n1076), .B1(n388), .Y(n393) );
  OAI22XL U326 ( .A0(n1079), .A1(n561), .B0(n1101), .B1(n525), .Y(n568) );
  NOR2BXL U327 ( .AN(B[0]), .B(n1030), .Y(n77) );
  OAI22XL U328 ( .A0(n807), .A1(n79), .B0(n805), .B1(n74), .Y(n75) );
  INVXL U329 ( .A(n1166), .Y(n1167) );
  AOI21XL U330 ( .A0(n1165), .A1(n1164), .B0(n1163), .Y(n1166) );
  INVXL U331 ( .A(n1176), .Y(n1163) );
  OAI2BB1XL U332 ( .A0N(n1076), .A1N(n1075), .B0(n1074), .Y(n1080) );
  OAI22XL U333 ( .A0(n1118), .A1(n1072), .B0(n1116), .B1(n1077), .Y(n1081) );
  INVXL U334 ( .A(n1073), .Y(n1074) );
  OAI22XL U335 ( .A0(n1079), .A1(n1047), .B0(n1101), .B1(n1068), .Y(n1071) );
  INVXL U336 ( .A(n1082), .Y(n1069) );
  OAI22XL U337 ( .A0(n1118), .A1(n1048), .B0(n1116), .B1(n1072), .Y(n1070) );
  OAI22XL U338 ( .A0(n1079), .A1(n385), .B0(n1101), .B1(n1032), .Y(n1035) );
  OAI22XL U339 ( .A0(n1118), .A1(n386), .B0(n1116), .B1(n1026), .Y(n1034) );
  INVXL U340 ( .A(n1045), .Y(n1033) );
  ADDFX2 U341 ( .A(n890), .B(n889), .CI(n888), .CO(n877), .S(n901) );
  ADDFX2 U342 ( .A(n226), .B(n225), .CI(n224), .CO(n893), .S(n269) );
  NOR2BXL U343 ( .AN(B[0]), .B(n799), .Y(n137) );
  OAI22XL U344 ( .A0(n792), .A1(n127), .B0(n791), .B1(n126), .Y(n135) );
  OAI22XL U345 ( .A0(n784), .A1(n125), .B0(n124), .B1(n1000), .Y(n136) );
  ADDFX2 U346 ( .A(n107), .B(n37), .CI(n105), .CO(n143), .S(n142) );
  OAI22XL U347 ( .A0(n792), .A1(n108), .B0(n791), .B1(n98), .Y(n107) );
  ADDFX2 U348 ( .A(n87), .B(n86), .CI(n85), .CO(n150), .S(n149) );
  ADDFX2 U349 ( .A(n97), .B(n96), .CI(n95), .CO(n148), .S(n144) );
  NOR2XL U350 ( .A(n131), .B(n130), .Y(n1139) );
  AOI21XL U351 ( .A0(n1145), .A1(n120), .B0(n123), .Y(n1142) );
  INVXL U352 ( .A(n1144), .Y(n123) );
  NAND2XL U353 ( .A(n131), .B(n130), .Y(n1140) );
  OAI22XL U354 ( .A0(n1118), .A1(n1117), .B0(n1116), .B1(n1115), .Y(n1119) );
  OAI2BB1XL U355 ( .A0N(n1101), .A1N(n1100), .B0(n1099), .Y(n1110) );
  OAI22XL U356 ( .A0(n1118), .A1(n1097), .B0(n1116), .B1(n1117), .Y(n1111) );
  INVXL U357 ( .A(n1098), .Y(n1099) );
  OAI22XL U358 ( .A0(n784), .A1(B[0]), .B0(n113), .B1(n1000), .Y(n1152) );
  NAND2XL U359 ( .A(n114), .B(n784), .Y(n1151) );
  NAND2BXL U360 ( .AN(B[0]), .B(n485), .Y(n114) );
  NAND2XL U361 ( .A(n1152), .B(n1151), .Y(n1153) );
  NAND2XL U362 ( .A(n139), .B(n138), .Y(n1158) );
  INVXL U363 ( .A(n1169), .Y(n1155) );
  INVXL U364 ( .A(n1188), .Y(n346) );
  INVXL U365 ( .A(n1187), .Y(n404) );
  INVXL U366 ( .A(n1192), .Y(n431) );
  INVXL U367 ( .A(n1182), .Y(n1059) );
  INVXL U368 ( .A(n1196), .Y(n506) );
  INVXL U369 ( .A(n1195), .Y(n545) );
  NAND2XL U370 ( .A(n770), .B(n644), .Y(n689) );
  AOI21XL U371 ( .A0(n6), .A1(n771), .B0(n728), .Y(n729) );
  INVXL U372 ( .A(n1208), .Y(n728) );
  NAND2XL U373 ( .A(n770), .B(n771), .Y(n730) );
  XNOR2XL U374 ( .A(n1114), .B(n702), .Y(n744) );
  XNOR2X1 U375 ( .A(n1114), .B(n743), .Y(n785) );
  INVXL U376 ( .A(n1067), .Y(n267) );
  NAND2BXL U377 ( .AN(B[0]), .B(n1049), .Y(n156) );
  XNOR2X1 U378 ( .A(n205), .B(B[23]), .Y(n622) );
  XNOR2XL U379 ( .A(n1114), .B(B[9]), .Y(n623) );
  XNOR2XL U380 ( .A(n1114), .B(B[10]), .Y(n591) );
  AOI21XL U381 ( .A0(n1059), .A1(n1058), .B0(n1057), .Y(n1105) );
  INVXL U382 ( .A(n1180), .Y(n1057) );
  NAND2XL U383 ( .A(n1156), .B(n1058), .Y(n1104) );
  INVXL U384 ( .A(n1201), .Y(n652) );
  OAI21X1 U385 ( .A0(n26), .A1(n859), .B0(n858), .Y(n861) );
  INVXL U386 ( .A(n857), .Y(n859) );
  XNOR2X1 U387 ( .A(n1049), .B(n704), .Y(n673) );
  XNOR2XL U388 ( .A(n757), .B(B[16]), .Y(n674) );
  OAI22X1 U389 ( .A0(n784), .A1(n701), .B0(n663), .B1(n1000), .Y(n700) );
  XNOR2X1 U390 ( .A(n1049), .B(n745), .Y(n714) );
  XNOR2XL U391 ( .A(n365), .B(B[16]), .Y(n754) );
  XNOR2XL U392 ( .A(n1049), .B(B[10]), .Y(n755) );
  XNOR2X1 U393 ( .A(n757), .B(B[14]), .Y(n758) );
  XNOR2X1 U394 ( .A(n205), .B(B[18]), .Y(n783) );
  XNOR2XL U395 ( .A(n746), .B(B[10]), .Y(n789) );
  XOR2XL U396 ( .A(B[16]), .B(n7), .Y(n45) );
  XNOR2XL U397 ( .A(n1067), .B(n702), .Y(n794) );
  XNOR2X1 U398 ( .A(n753), .B(n437), .Y(n54) );
  XNOR2XL U399 ( .A(n746), .B(B[9]), .Y(n231) );
  XNOR2XL U400 ( .A(n757), .B(n745), .Y(n201) );
  XNOR2XL U401 ( .A(n1049), .B(n702), .Y(n220) );
  XNOR2XL U402 ( .A(n757), .B(B[10]), .Y(n222) );
  XNOR2XL U403 ( .A(n437), .B(B[9]), .Y(n288) );
  NAND2BXL U404 ( .AN(B[0]), .B(n746), .Y(n71) );
  XNOR2XL U405 ( .A(n757), .B(B[4]), .Y(n173) );
  XNOR2X1 U406 ( .A(B[10]), .B(n485), .Y(n159) );
  XNOR2XL U407 ( .A(n437), .B(B[7]), .Y(n172) );
  NAND2BXL U408 ( .AN(B[0]), .B(n1114), .Y(n206) );
  NOR2BXL U409 ( .AN(B[0]), .B(n1101), .Y(n322) );
  OAI22XL U410 ( .A0(n1051), .A1(n285), .B0(n1076), .B1(n284), .Y(n320) );
  XNOR2XL U411 ( .A(n757), .B(B[22]), .Y(n453) );
  XNOR2XL U412 ( .A(n1114), .B(n704), .Y(n519) );
  XNOR2X1 U413 ( .A(n746), .B(B[19]), .Y(n483) );
  XNOR2X1 U414 ( .A(n746), .B(B[18]), .Y(n522) );
  XNOR2XL U415 ( .A(n365), .B(B[4]), .Y(n67) );
  XNOR2XL U416 ( .A(n485), .B(B[8]), .Y(n72) );
  INVXL U417 ( .A(n1186), .Y(n1009) );
  INVXL U418 ( .A(n1184), .Y(n1008) );
  NAND2XL U419 ( .A(n1064), .B(n1178), .Y(n1065) );
  INVXL U420 ( .A(n1177), .Y(n1064) );
  XNOR2XL U421 ( .A(n1049), .B(n1113), .Y(n1073) );
  XNOR2X1 U422 ( .A(n1096), .B(B[19]), .Y(n386) );
  XNOR2XL U423 ( .A(n1067), .B(B[21]), .Y(n385) );
  OAI22XL U424 ( .A0(n1079), .A1(n594), .B0(n1101), .B1(n561), .Y(n601) );
  OAI22XL U425 ( .A0(n1029), .A1(n592), .B0(n1030), .B1(n559), .Y(n603) );
  OAI22X1 U426 ( .A0(n792), .A1(n593), .B0(n791), .B1(n560), .Y(n602) );
  ADDFX2 U427 ( .A(n638), .B(n637), .CI(n636), .CO(n660), .S(n696) );
  OAI22X1 U428 ( .A0(n1051), .A1(n631), .B0(n1076), .B1(n599), .Y(n637) );
  OAI22XL U429 ( .A0(n801), .A1(n630), .B0(n799), .B1(n598), .Y(n638) );
  OAI22XL U430 ( .A0(n1079), .A1(n626), .B0(n1101), .B1(n594), .Y(n633) );
  OAI22X1 U431 ( .A0(n792), .A1(n625), .B0(n791), .B1(n593), .Y(n634) );
  OAI22XL U432 ( .A0(n1079), .A1(n668), .B0(n1101), .B1(n626), .Y(n675) );
  ADDFX2 U433 ( .A(n680), .B(n679), .CI(n678), .CO(n698), .S(n737) );
  OAI22XL U434 ( .A0(n716), .A1(n674), .B0(n805), .B1(n632), .Y(n678) );
  OAI22X1 U435 ( .A0(n1051), .A1(n673), .B0(n1076), .B1(n631), .Y(n679) );
  ADDFX2 U436 ( .A(n722), .B(n721), .CI(n720), .CO(n739), .S(n777) );
  OAI22XL U437 ( .A0(n807), .A1(n715), .B0(n805), .B1(n674), .Y(n720) );
  OAI22XL U438 ( .A0(n1051), .A1(n714), .B0(n1076), .B1(n673), .Y(n721) );
  OAI22X1 U439 ( .A0(n801), .A1(n713), .B0(n799), .B1(n672), .Y(n722) );
  OAI22XL U440 ( .A0(n1079), .A1(n709), .B0(n1101), .B1(n668), .Y(n717) );
  OAI22XL U441 ( .A0(n1079), .A1(n749), .B0(n1101), .B1(n709), .Y(n759) );
  OAI22XL U442 ( .A0(n716), .A1(n758), .B0(n805), .B1(n715), .Y(n762) );
  OAI22XL U443 ( .A0(n1079), .A1(n793), .B0(n1101), .B1(n749), .Y(n808) );
  OAI22XL U444 ( .A0(n807), .A1(n806), .B0(n805), .B1(n804), .Y(n849) );
  ADDFX2 U445 ( .A(n848), .B(n847), .CI(n846), .CO(n840), .S(n889) );
  OAI22XL U446 ( .A0(n1079), .A1(n794), .B0(n1101), .B1(n793), .Y(n846) );
  OAI22X1 U447 ( .A0(n790), .A1(n791), .B0(n792), .B1(n45), .Y(n847) );
  OAI22XL U448 ( .A0(n1029), .A1(n789), .B0(n1030), .B1(n788), .Y(n848) );
  CMPR32X1 U449 ( .A(n839), .B(n838), .C(n837), .CO(n871), .S(n875) );
  OAI22XL U450 ( .A0(n1079), .A1(n234), .B0(n1101), .B1(n794), .Y(n837) );
  OAI22XL U451 ( .A0(n1029), .A1(n231), .B0(n1030), .B1(n789), .Y(n839) );
  OAI22X1 U452 ( .A0(n54), .A1(n792), .B0(n45), .B1(n791), .Y(n838) );
  OAI22XL U453 ( .A0(n807), .A1(n264), .B0(n805), .B1(n223), .Y(n290) );
  OAI22XL U454 ( .A0(n1051), .A1(n258), .B0(n1076), .B1(n221), .Y(n291) );
  OAI22XL U455 ( .A0(n1079), .A1(n252), .B0(n1101), .B1(n214), .Y(n260) );
  OAI22XL U456 ( .A0(n1118), .A1(n204), .B0(n1116), .B1(n208), .Y(n261) );
  OAI22X1 U457 ( .A0(n666), .A1(n256), .B0(n1030), .B1(n213), .Y(n262) );
  ADDFX2 U458 ( .A(n306), .B(n305), .CI(n304), .CO(n273), .S(n307) );
  OAI22X1 U459 ( .A0(n1051), .A1(n277), .B0(n1076), .B1(n258), .Y(n305) );
  OAI22XL U460 ( .A0(n666), .A1(n299), .B0(n1030), .B1(n256), .Y(n306) );
  ADDFX2 U461 ( .A(n298), .B(n297), .CI(n296), .CO(n293), .S(n309) );
  NOR2BXL U462 ( .AN(B[0]), .B(n1116), .Y(n298) );
  OAI22XL U463 ( .A0(n1079), .A1(n275), .B0(n1101), .B1(n252), .Y(n296) );
  CMPR32X1 U464 ( .A(n280), .B(n279), .C(n278), .CO(n271), .S(n324) );
  OAI22XL U465 ( .A0(n1051), .A1(n284), .B0(n1076), .B1(n277), .Y(n310) );
  OAI22XL U466 ( .A0(n1079), .A1(n276), .B0(n1101), .B1(n275), .Y(n311) );
  OAI22XL U467 ( .A0(n807), .A1(n286), .B0(n805), .B1(n274), .Y(n312) );
  CMPR32X1 U468 ( .A(n458), .B(n457), .C(n456), .CO(n479), .S(n516) );
  OAI2BB1XL U469 ( .A0N(n524), .A1N(n707), .B0(n439), .Y(n456) );
  OAI2BB1XL U470 ( .A0N(n493), .A1N(n42), .B0(n41), .Y(n487) );
  OAI22XL U471 ( .A0(n1029), .A1(n449), .B0(n1030), .B1(n412), .Y(n440) );
  OAI22XL U472 ( .A0(n1100), .A1(n411), .B0(n1101), .B1(n377), .Y(n414) );
  OAI22XL U473 ( .A0(n1100), .A1(n377), .B0(n1101), .B1(n373), .Y(n381) );
  ADDFX2 U474 ( .A(n497), .B(n496), .CI(n495), .CO(n517), .S(n551) );
  OAI22XL U475 ( .A0(n1029), .A1(n483), .B0(n1030), .B1(n455), .Y(n495) );
  OAI22X1 U476 ( .A0(n1118), .A1(n484), .B0(n1116), .B1(n454), .Y(n496) );
  OAI22X1 U477 ( .A0(n807), .A1(n481), .B0(n805), .B1(n453), .Y(n497) );
  OAI22XL U478 ( .A0(n1100), .A1(n482), .B0(n1101), .B1(n480), .Y(n528) );
  OAI22XL U479 ( .A0(n807), .A1(n600), .B0(n805), .B1(n567), .Y(n604) );
  OAI22XL U480 ( .A0(n801), .A1(n598), .B0(n799), .B1(n565), .Y(n606) );
  CMPR32X1 U481 ( .A(n671), .B(n670), .C(n669), .CO(n683), .S(n724) );
  ADDFX2 U482 ( .A(n629), .B(n628), .CI(n627), .CO(n641), .S(n682) );
  OAI22XL U483 ( .A0(n792), .A1(n523), .B0(n524), .B1(n490), .Y(n537) );
  OAI22XL U484 ( .A0(n1075), .A1(n530), .B0(n1076), .B1(n491), .Y(n536) );
  CMPR32X1 U485 ( .A(n534), .B(n533), .C(n532), .CO(n526), .S(n586) );
  OAI2BB1XL U486 ( .A0N(n1000), .A1N(n784), .B0(n486), .Y(n532) );
  OAI22XL U487 ( .A0(n807), .A1(n567), .B0(n805), .B1(n531), .Y(n571) );
  OAI22XL U488 ( .A0(n801), .A1(n565), .B0(n799), .B1(n529), .Y(n573) );
  ADDFX2 U489 ( .A(n564), .B(n563), .CI(n562), .CO(n576), .S(n608) );
  INVXL U490 ( .A(n757), .Y(n369) );
  OAI22XL U491 ( .A0(n801), .A1(n94), .B0(n799), .B1(n81), .Y(n90) );
  OAI22XL U492 ( .A0(n807), .A1(n80), .B0(n805), .B1(n79), .Y(n91) );
  OAI22X1 U493 ( .A0(n792), .A1(n98), .B0(n791), .B1(n78), .Y(n92) );
  OAI22XL U494 ( .A0(n1051), .A1(n388), .B0(n1076), .B1(n1031), .Y(n1038) );
  OAI22XL U495 ( .A0(n1079), .A1(n1032), .B0(n1101), .B1(n1047), .Y(n1053) );
  OAI22XL U496 ( .A0(n1051), .A1(n1031), .B0(n1076), .B1(n1050), .Y(n1054) );
  OAI2BB1XL U497 ( .A0N(n1030), .A1N(n1029), .B0(n1028), .Y(n1044) );
  OAI22XL U498 ( .A0(n1118), .A1(n1026), .B0(n1116), .B1(n1048), .Y(n1046) );
  INVXL U499 ( .A(n1027), .Y(n1028) );
  ADDFX2 U500 ( .A(n969), .B(n968), .CI(n967), .CO(n975), .S(n973) );
  NAND2XL U501 ( .A(n955), .B(n956), .Y(n51) );
  XOR3X2 U502 ( .A(n956), .B(n955), .C(n954), .Y(n957) );
  ADDFX2 U503 ( .A(n962), .B(n961), .CI(n960), .CO(n970), .S(n194) );
  NAND2X1 U504 ( .A(n48), .B(n47), .Y(n961) );
  OAI21XL U505 ( .A0(n184), .A1(n182), .B0(n183), .Y(n48) );
  XOR3X2 U506 ( .A(n184), .B(n182), .C(n183), .Y(n185) );
  ADDFX2 U507 ( .A(n421), .B(n420), .CI(n419), .CO(n467), .S(n462) );
  OAI22XL U508 ( .A0(n1029), .A1(n412), .B0(n1030), .B1(n407), .Y(n421) );
  ADDFX2 U509 ( .A(n464), .B(n463), .CI(n462), .CO(n466), .S(n474) );
  OAI22XL U510 ( .A0(n1051), .A1(n378), .B0(n1076), .B1(n374), .Y(n384) );
  OAI22XL U511 ( .A0(n1118), .A1(n363), .B0(n1116), .B1(n370), .Y(n383) );
  ADDFX2 U512 ( .A(n424), .B(n423), .CI(n422), .CO(n425), .S(n465) );
  OAI22XL U513 ( .A0(n784), .A1(n113), .B0(n117), .B1(n1000), .Y(n116) );
  NOR2BXL U514 ( .AN(B[0]), .B(n791), .Y(n115) );
  OAI22XL U515 ( .A0(n792), .A1(n7), .B0(n524), .B1(n119), .Y(n121) );
  NAND2BXL U516 ( .AN(B[0]), .B(n437), .Y(n119) );
  OAI22XL U517 ( .A0(n303), .A1(n110), .B0(n799), .B1(n109), .Y(n133) );
  OAI22XL U518 ( .A0(n792), .A1(n126), .B0(n791), .B1(n108), .Y(n134) );
  AOI21XL U519 ( .A0(n1160), .A1(n1159), .B0(n140), .Y(n1129) );
  INVXL U520 ( .A(n1158), .Y(n140) );
  NAND2XL U521 ( .A(n1007), .B(n1168), .Y(n1171) );
  INVXL U522 ( .A(n963), .Y(n983) );
  OAI22XL U523 ( .A0(n1118), .A1(n1077), .B0(n1116), .B1(n1097), .Y(n1095) );
  INVXL U524 ( .A(n1112), .Y(n1094) );
  OAI22XL U525 ( .A0(n1079), .A1(n1068), .B0(n1101), .B1(n1078), .Y(n1090) );
  ADDFX2 U526 ( .A(n1043), .B(n1042), .CI(n1041), .CO(n1056), .S(n1039) );
  NAND2X1 U527 ( .A(n39), .B(n38), .Y(n855) );
  OAI21XL U528 ( .A0(n863), .A1(n864), .B0(n862), .Y(n39) );
  XOR2X1 U529 ( .A(n862), .B(n864), .Y(n40) );
  OAI2BB1X1 U530 ( .A0N(n56), .A1N(n891), .B0(n55), .Y(n900) );
  XOR2X1 U531 ( .A(n891), .B(n58), .Y(n902) );
  XOR2X1 U532 ( .A(n892), .B(n893), .Y(n58) );
  ADDFX2 U533 ( .A(n912), .B(n911), .CI(n910), .CO(n916), .S(n922) );
  OAI21XL U534 ( .A0(n615), .A1(n616), .B0(n614), .Y(n50) );
  XOR3X2 U535 ( .A(n616), .B(n614), .C(n615), .Y(n643) );
  NOR2XL U536 ( .A(n116), .B(n115), .Y(n1147) );
  NAND2XL U537 ( .A(n116), .B(n115), .Y(n1148) );
  NAND2XL U538 ( .A(n122), .B(n121), .Y(n1144) );
  INVXL U539 ( .A(n1129), .Y(n1137) );
  NAND2XL U540 ( .A(n1084), .B(n1083), .Y(mult_x_1_n115) );
  XOR2XL U541 ( .A(n1143), .B(n1142), .Y(n1255) );
  NAND2XL U542 ( .A(n1141), .B(n1140), .Y(n1143) );
  INVXL U543 ( .A(n1139), .Y(n1141) );
  NAND2XL U544 ( .A(n997), .B(n996), .Y(n998) );
  NOR2XL U545 ( .A(n1040), .B(n1039), .Y(mult_x_1_n149) );
  NAND2XL U546 ( .A(n1123), .B(n1122), .Y(mult_x_1_n54) );
  NAND2XL U547 ( .A(n1121), .B(n1120), .Y(n1122) );
  INVXL U548 ( .A(n1119), .Y(n1120) );
  NOR2XL U549 ( .A(n1103), .B(n1102), .Y(mult_x_1_n105) );
  NAND2XL U550 ( .A(n1103), .B(n1102), .Y(mult_x_1_n106) );
  NOR2XL U551 ( .A(n1084), .B(n1083), .Y(mult_x_1_n114) );
  NOR2XL U552 ( .A(n1092), .B(n1091), .Y(mult_x_1_n125) );
  NAND2XL U553 ( .A(n1092), .B(n1091), .Y(mult_x_1_n126) );
  NOR2XL U554 ( .A(n1056), .B(n1055), .Y(mult_x_1_n134) );
  NAND2XL U555 ( .A(n1056), .B(n1055), .Y(mult_x_1_n135) );
  NAND2XL U556 ( .A(n1040), .B(n1039), .Y(mult_x_1_n150) );
  NOR2XL U557 ( .A(n927), .B(mult_x_1_n312), .Y(mult_x_1_n305) );
  NAND2XL U558 ( .A(n1003), .B(n1002), .Y(mult_x_1_n80) );
  INVXL U559 ( .A(n1001), .Y(n1003) );
  OAI21XL U560 ( .A0(n927), .A1(mult_x_1_n313), .B0(n928), .Y(mult_x_1_n306)
         );
  AND2XL U561 ( .A(n1154), .B(n1153), .Y(n1258) );
  XOR2XL U562 ( .A(n1150), .B(n1153), .Y(n1257) );
  NAND2XL U563 ( .A(n1149), .B(n1148), .Y(n1150) );
  INVXL U564 ( .A(n1147), .Y(n1149) );
  XNOR2XL U565 ( .A(n1146), .B(n1145), .Y(n1256) );
  NAND2XL U566 ( .A(n120), .B(n1144), .Y(n1146) );
  NAND2XL U567 ( .A(n1159), .B(n1158), .Y(n1161) );
  NAND2XL U568 ( .A(n1136), .B(n1135), .Y(n1138) );
  AOI21XL U569 ( .A0(n1137), .A1(n1136), .B0(n1130), .Y(n1134) );
  NAND2XL U570 ( .A(n1132), .B(n1131), .Y(n1133) );
  NOR2BXL U571 ( .AN(B[0]), .B(n1000), .Y(n1259) );
  NAND2XL U572 ( .A(n1126), .B(n1125), .Y(n1127) );
  INVXL U573 ( .A(n1124), .Y(n1126) );
  OR2X2 U574 ( .A(n194), .B(n193), .Y(n36) );
  BUFX3 U575 ( .A(A[7]), .Y(n757) );
  XOR2X1 U576 ( .A(n756), .B(n364), .Y(n46) );
  AOI21X1 U577 ( .A0(n993), .A1(n5), .B0(n987), .Y(n990) );
  OAI21XL U578 ( .A0(n147), .A1(n1129), .B0(n146), .Y(n994) );
  AOI21X1 U579 ( .A0(n1132), .A1(n1130), .B0(n145), .Y(n146) );
  XNOR2X1 U580 ( .A(n437), .B(n743), .Y(n78) );
  CMPR22X1 U581 ( .A(n89), .B(n88), .CO(n82), .S(n97) );
  OAI22X1 U582 ( .A0(n784), .A1(n93), .B0(n73), .B1(n1000), .Y(n89) );
  OAI22X1 U583 ( .A0(n557), .A1(n207), .B0(n209), .B1(n1000), .Y(n212) );
  XNOR2X1 U584 ( .A(n205), .B(B[16]), .Y(n209) );
  OAI22X1 U585 ( .A0(n1118), .A1(n558), .B0(n1116), .B1(n519), .Y(n554) );
  OAI22X1 U586 ( .A0(n787), .A1(n623), .B0(n1116), .B1(n591), .Y(n620) );
  OAI22X1 U587 ( .A0(n787), .A1(n664), .B0(n1116), .B1(n623), .Y(n661) );
  OAI22X1 U588 ( .A0(n807), .A1(n169), .B0(n805), .B1(n173), .Y(n178) );
  OAI22X1 U589 ( .A0(n1029), .A1(n788), .B0(n1030), .B1(n747), .Y(n810) );
  XNOR2X1 U590 ( .A(n757), .B(B[21]), .Y(n481) );
  OAI22X1 U591 ( .A0(n716), .A1(n376), .B0(n805), .B1(n371), .Y(n390) );
  BUFX1 U592 ( .A(n106), .Y(n37) );
  OAI22X1 U593 ( .A0(n784), .A1(n283), .B0(n265), .B1(n1000), .Y(n282) );
  XOR2X1 U594 ( .A(n924), .B(n1223), .Y(PRODUCT[16]) );
  OAI22X1 U595 ( .A0(n1118), .A1(n591), .B0(n1116), .B1(n558), .Y(n588) );
  OAI22X1 U596 ( .A0(n787), .A1(n703), .B0(n1116), .B1(n664), .Y(n699) );
  OAI22X1 U597 ( .A0(n792), .A1(n70), .B0(n791), .B1(n172), .Y(n181) );
  ADDFX2 U598 ( .A(n165), .B(n164), .CI(n163), .CO(n182), .S(n190) );
  OAI22X1 U599 ( .A0(n807), .A1(n74), .B0(n805), .B1(n169), .Y(n165) );
  CMPR22X1 U600 ( .A(n555), .B(n554), .CO(n564), .S(n597) );
  OAI22X1 U601 ( .A0(n557), .A1(n556), .B0(n518), .B1(n1000), .Y(n555) );
  CMPR22X1 U602 ( .A(n230), .B(n229), .CO(n869), .S(n226) );
  CMPR22X1 U603 ( .A(n212), .B(n211), .CO(n225), .S(n253) );
  BUFX3 U604 ( .A(A[9]), .Y(n746) );
  XOR2X1 U605 ( .A(n40), .B(n863), .Y(n881) );
  NAND2XL U606 ( .A(n494), .B(n44), .Y(n41) );
  XOR2X1 U607 ( .A(n493), .B(n43), .Y(n552) );
  XOR2X1 U608 ( .A(n494), .B(n44), .Y(n43) );
  OAI22X1 U609 ( .A0(n492), .A1(n801), .B0(n799), .B1(n452), .Y(n44) );
  OAI22X1 U610 ( .A0(n801), .A1(n446), .B0(n799), .B1(n366), .Y(n417) );
  ADDFHX4 U611 ( .A(n255), .B(n254), .CI(n253), .CO(n270), .S(n333) );
  OAI22X1 U612 ( .A0(n784), .A1(n73), .B0(n72), .B1(n1000), .Y(n76) );
  XNOR2X2 U613 ( .A(n485), .B(B[14]), .Y(n251) );
  XNOR2X4 U614 ( .A(n547), .B(n546), .Y(PRODUCT[29]) );
  OAI22XL U615 ( .A0(n1029), .A1(n624), .B0(n1030), .B1(n592), .Y(n635) );
  INVX1 U616 ( .A(n645), .Y(n770) );
  AOI21XL U617 ( .A0(n346), .A1(n1004), .B0(n1009), .Y(n347) );
  AOI21XL U618 ( .A0(n1010), .A1(n1009), .B0(n1008), .Y(n1011) );
  NAND2XL U619 ( .A(n649), .B(n770), .Y(n651) );
  XNOR2XL U620 ( .A(n1096), .B(B[22]), .Y(n1072) );
  NOR2X1 U621 ( .A(n917), .B(n916), .Y(mult_x_1_n299) );
  XOR2XL U622 ( .A(A[6]), .B(A[7]), .Y(n59) );
  XNOR2XL U623 ( .A(A[6]), .B(A[5]), .Y(n60) );
  NAND2X1 U624 ( .A(n59), .B(n60), .Y(n716) );
  BUFX3 U625 ( .A(n716), .Y(n807) );
  XNOR2XL U626 ( .A(n757), .B(B[2]), .Y(n74) );
  BUFX3 U627 ( .A(n60), .Y(n805) );
  XNOR2X1 U628 ( .A(n757), .B(n257), .Y(n169) );
  XOR2XL U629 ( .A(A[8]), .B(A[9]), .Y(n61) );
  BUFX3 U630 ( .A(n666), .Y(n1029) );
  XNOR2XL U631 ( .A(n746), .B(B[0]), .Y(n63) );
  BUFX3 U632 ( .A(n62), .Y(n1030) );
  XNOR2XL U633 ( .A(n746), .B(B[1]), .Y(n162) );
  XOR2XL U634 ( .A(A[4]), .B(A[5]), .Y(n64) );
  XNOR2XL U635 ( .A(A[4]), .B(A[3]), .Y(n65) );
  BUFX3 U636 ( .A(n303), .Y(n801) );
  BUFX3 U637 ( .A(n65), .Y(n799) );
  BUFX3 U638 ( .A(B[5]), .Y(n743) );
  XNOR2X1 U639 ( .A(n365), .B(n743), .Y(n171) );
  XOR2XL U640 ( .A(A[2]), .B(A[3]), .Y(n66) );
  XNOR2X1 U641 ( .A(A[2]), .B(n485), .Y(n524) );
  NAND2X1 U642 ( .A(n66), .B(n524), .Y(n707) );
  BUFX3 U643 ( .A(n707), .Y(n792) );
  BUFX3 U644 ( .A(n524), .Y(n791) );
  BUFX3 U645 ( .A(B[6]), .Y(n702) );
  XNOR2X1 U646 ( .A(n437), .B(n702), .Y(n70) );
  OAI22XL U647 ( .A0(n792), .A1(n78), .B0(n791), .B1(n70), .Y(n84) );
  XNOR2X1 U648 ( .A(n365), .B(n257), .Y(n81) );
  OAI22XL U649 ( .A0(n303), .A1(n81), .B0(n799), .B1(n67), .Y(n83) );
  NAND2X1 U650 ( .A(A[1]), .B(n68), .Y(n557) );
  BUFX3 U651 ( .A(n557), .Y(n784) );
  XNOR2X1 U652 ( .A(n485), .B(B[7]), .Y(n73) );
  BUFX3 U653 ( .A(n68), .Y(n1000) );
  OAI22X1 U654 ( .A0(n807), .A1(n369), .B0(n805), .B1(n69), .Y(n88) );
  XNOR2X1 U655 ( .A(n485), .B(B[9]), .Y(n160) );
  OAI22X1 U656 ( .A0(n784), .A1(n72), .B0(n160), .B1(n1000), .Y(n158) );
  OAI22X1 U657 ( .A0(n1029), .A1(n368), .B0(n1030), .B1(n71), .Y(n157) );
  XNOR2XL U658 ( .A(n757), .B(B[1]), .Y(n79) );
  CMPR32X1 U659 ( .A(n77), .B(n76), .C(n75), .CO(n179), .S(n87) );
  XNOR2XL U660 ( .A(n437), .B(B[4]), .Y(n98) );
  XNOR2XL U661 ( .A(n757), .B(B[0]), .Y(n80) );
  XNOR2XL U662 ( .A(n365), .B(B[2]), .Y(n94) );
  CMPR32X1 U663 ( .A(n84), .B(n83), .C(n82), .CO(n189), .S(n85) );
  CMPR32X1 U664 ( .A(n92), .B(n91), .C(n90), .CO(n86), .S(n96) );
  XNOR2X1 U665 ( .A(n485), .B(n743), .Y(n99) );
  OAI22XL U666 ( .A0(n784), .A1(n99), .B0(n93), .B1(n1000), .Y(n102) );
  XNOR2XL U667 ( .A(n365), .B(B[1]), .Y(n109) );
  NOR2XL U668 ( .A(n995), .B(n1124), .Y(n153) );
  XNOR2XL U669 ( .A(n485), .B(B[4]), .Y(n124) );
  OAI22XL U670 ( .A0(n784), .A1(n124), .B0(n99), .B1(n1000), .Y(n112) );
  CMPR32X1 U671 ( .A(n103), .B(n102), .C(n101), .CO(n95), .S(n105) );
  NOR2X1 U672 ( .A(n144), .B(n143), .Y(n104) );
  XNOR2XL U673 ( .A(n437), .B(B[2]), .Y(n126) );
  XNOR2XL U674 ( .A(n365), .B(B[0]), .Y(n110) );
  ADDHXL U675 ( .A(n112), .B(n111), .CO(n106), .S(n132) );
  OR2X2 U676 ( .A(n142), .B(n141), .Y(n1136) );
  NAND2XL U677 ( .A(n1132), .B(n1136), .Y(n147) );
  XNOR2XL U678 ( .A(n485), .B(B[1]), .Y(n113) );
  XNOR2XL U679 ( .A(n485), .B(B[2]), .Y(n117) );
  OAI21XL U680 ( .A0(n1147), .A1(n1153), .B0(n1148), .Y(n1145) );
  OAI22X1 U681 ( .A0(n784), .A1(n117), .B0(n125), .B1(n1000), .Y(n129) );
  XNOR2XL U682 ( .A(n437), .B(B[0]), .Y(n118) );
  XNOR2XL U683 ( .A(n437), .B(B[1]), .Y(n127) );
  OAI22X1 U684 ( .A0(n792), .A1(n118), .B0(n791), .B1(n127), .Y(n128) );
  CMPR22X1 U685 ( .A(n129), .B(n128), .CO(n130), .S(n122) );
  OAI21XL U686 ( .A0(n1142), .A1(n1139), .B0(n1140), .Y(n1160) );
  CMPR32X1 U687 ( .A(n134), .B(n133), .C(n132), .CO(n141), .S(n139) );
  CMPR32X1 U688 ( .A(n137), .B(n136), .C(n135), .CO(n138), .S(n131) );
  OR2X2 U689 ( .A(n139), .B(n138), .Y(n1159) );
  NAND2XL U690 ( .A(n142), .B(n141), .Y(n1135) );
  INVXL U691 ( .A(n1135), .Y(n1130) );
  NAND2XL U692 ( .A(n144), .B(n143), .Y(n1131) );
  INVXL U693 ( .A(n1131), .Y(n145) );
  NAND2XL U694 ( .A(n151), .B(n150), .Y(n996) );
  OAI21XL U695 ( .A0(n995), .A1(n1125), .B0(n996), .Y(n152) );
  AOI21X1 U696 ( .A0(n153), .A1(n994), .B0(n152), .Y(n986) );
  XNOR2X1 U697 ( .A(n365), .B(n702), .Y(n170) );
  XNOR2X1 U698 ( .A(n365), .B(B[7]), .Y(n289) );
  OAI22XL U699 ( .A0(n303), .A1(n170), .B0(n799), .B1(n289), .Y(n941) );
  XNOR2XL U700 ( .A(n746), .B(B[2]), .Y(n161) );
  XNOR2X1 U701 ( .A(n746), .B(n257), .Y(n317) );
  OAI22XL U702 ( .A0(n1029), .A1(n161), .B0(n1030), .B1(n317), .Y(n940) );
  BUFX3 U703 ( .A(B[11]), .Y(n745) );
  BUFX3 U704 ( .A(n1075), .Y(n1051) );
  BUFX3 U705 ( .A(n155), .Y(n1076) );
  OAI22X1 U706 ( .A0(n1051), .A1(n361), .B0(n1076), .B1(n156), .Y(n318) );
  CMPR22X1 U707 ( .A(n158), .B(n157), .CO(n184), .S(n180) );
  OAI22X1 U708 ( .A0(n784), .A1(n160), .B0(n159), .B1(n1000), .Y(n167) );
  ADDFHX1 U709 ( .A(n168), .B(n167), .CI(n166), .CO(n953), .S(n183) );
  OAI22X1 U710 ( .A0(n801), .A1(n171), .B0(n799), .B1(n170), .Y(n177) );
  BUFX3 U711 ( .A(B[8]), .Y(n708) );
  XNOR2X1 U712 ( .A(n437), .B(n708), .Y(n175) );
  OAI22XL U713 ( .A0(n792), .A1(n172), .B0(n791), .B1(n175), .Y(n176) );
  XNOR2X1 U714 ( .A(n757), .B(n743), .Y(n287) );
  OAI22XL U715 ( .A0(n807), .A1(n173), .B0(n805), .B1(n287), .Y(n938) );
  XNOR2XL U716 ( .A(n1049), .B(B[0]), .Y(n174) );
  XNOR2XL U717 ( .A(n1049), .B(B[1]), .Y(n285) );
  OAI22XL U718 ( .A0(n792), .A1(n175), .B0(n791), .B1(n288), .Y(n936) );
  CMPR32X1 U719 ( .A(n187), .B(n186), .C(n185), .CO(n193), .S(n192) );
  CMPR32X1 U720 ( .A(n190), .B(n189), .C(n188), .CO(n191), .S(n151) );
  NAND2XL U721 ( .A(n36), .B(n5), .Y(n197) );
  NAND2X1 U722 ( .A(n192), .B(n191), .Y(n991) );
  NAND2XL U723 ( .A(n194), .B(n193), .Y(n988) );
  INVXL U724 ( .A(n988), .Y(n195) );
  AOI21X1 U725 ( .A0(n36), .A1(n987), .B0(n195), .Y(n196) );
  BUFX3 U726 ( .A(B[12]), .Y(n704) );
  XNOR2X1 U727 ( .A(n365), .B(n704), .Y(n219) );
  BUFX3 U728 ( .A(B[13]), .Y(n756) );
  XNOR2X1 U729 ( .A(n1049), .B(B[7]), .Y(n200) );
  XOR2XL U730 ( .A(A[12]), .B(A[13]), .Y(n198) );
  BUFX3 U731 ( .A(n1100), .Y(n1079) );
  BUFX1 U732 ( .A(A[13]), .Y(n1067) );
  XNOR2X1 U733 ( .A(A[13]), .B(n743), .Y(n234) );
  BUFX3 U734 ( .A(n199), .Y(n1101) );
  XNOR2X1 U735 ( .A(n1049), .B(n708), .Y(n803) );
  OAI22XL U736 ( .A0(n1051), .A1(n200), .B0(n1076), .B1(n803), .Y(n844) );
  XNOR2X1 U737 ( .A(n746), .B(n702), .Y(n256) );
  XNOR2X1 U738 ( .A(n746), .B(B[7]), .Y(n213) );
  XOR2XL U739 ( .A(A[14]), .B(A[15]), .Y(n202) );
  XNOR2XL U740 ( .A(A[14]), .B(A[13]), .Y(n203) );
  NAND2X1 U741 ( .A(n202), .B(n203), .Y(n787) );
  BUFX3 U742 ( .A(n787), .Y(n1118) );
  CLKINVX3 U743 ( .A(n362), .Y(n1114) );
  XNOR2XL U744 ( .A(n1114), .B(B[0]), .Y(n204) );
  BUFX3 U745 ( .A(n203), .Y(n1116) );
  XNOR2XL U746 ( .A(n1114), .B(B[1]), .Y(n208) );
  XNOR2X1 U747 ( .A(A[13]), .B(n257), .Y(n214) );
  XNOR2X1 U748 ( .A(n205), .B(B[15]), .Y(n207) );
  OAI22X1 U749 ( .A0(n784), .A1(n251), .B0(n207), .B1(n1000), .Y(n250) );
  OAI22X1 U750 ( .A0(n1118), .A1(n362), .B0(n1116), .B1(n206), .Y(n249) );
  XNOR2XL U751 ( .A(n1114), .B(B[2]), .Y(n210) );
  OAI22X1 U752 ( .A0(n1118), .A1(n208), .B0(n1116), .B1(n210), .Y(n211) );
  OAI22X1 U753 ( .A0(n557), .A1(n209), .B0(n227), .B1(n1000), .Y(n230) );
  OAI22X1 U754 ( .A0(n1118), .A1(n210), .B0(n1116), .B1(n228), .Y(n229) );
  XNOR2X1 U755 ( .A(n746), .B(n708), .Y(n232) );
  OAI22XL U756 ( .A0(n1029), .A1(n213), .B0(n1030), .B1(n232), .Y(n218) );
  XNOR2X1 U757 ( .A(n437), .B(n756), .Y(n215) );
  XNOR2X1 U758 ( .A(n437), .B(B[14]), .Y(n233) );
  OAI22XL U759 ( .A0(n792), .A1(n215), .B0(n791), .B1(n233), .Y(n217) );
  XNOR2XL U760 ( .A(A[13]), .B(B[4]), .Y(n235) );
  XNOR2X1 U761 ( .A(n437), .B(n704), .Y(n259) );
  OAI22XL U762 ( .A0(n792), .A1(n259), .B0(n791), .B1(n215), .Y(n292) );
  XNOR2XL U763 ( .A(n1049), .B(B[4]), .Y(n258) );
  CMPR32X1 U764 ( .A(n218), .B(n217), .C(n216), .CO(n224), .S(n327) );
  XNOR2X1 U765 ( .A(n365), .B(n745), .Y(n248) );
  OAI22XL U766 ( .A0(n801), .A1(n248), .B0(n799), .B1(n219), .Y(n238) );
  OAI22XL U767 ( .A0(n1051), .A1(n221), .B0(n1076), .B1(n220), .Y(n237) );
  OAI22X1 U768 ( .A0(n784), .A1(n227), .B0(n783), .B1(n1000), .Y(n836) );
  XNOR2XL U769 ( .A(n1114), .B(B[4]), .Y(n786) );
  OAI22X1 U770 ( .A0(n1118), .A1(n228), .B0(n1116), .B1(n786), .Y(n835) );
  CMPR32X1 U771 ( .A(n238), .B(n237), .C(n236), .CO(n247), .S(n326) );
  CMPR32X1 U772 ( .A(n241), .B(n240), .C(n239), .CO(n868), .S(n246) );
  CMPR32X1 U773 ( .A(n244), .B(n243), .C(n242), .CO(n876), .S(n245) );
  CMPR32X1 U774 ( .A(n247), .B(n246), .C(n245), .CO(n891), .S(n912) );
  OAI22XL U775 ( .A0(n801), .A1(n263), .B0(n799), .B1(n248), .Y(n295) );
  CMPR22X1 U776 ( .A(n250), .B(n249), .CO(n254), .S(n294) );
  XNOR2X1 U777 ( .A(n485), .B(B[13]), .Y(n265) );
  OAI22X1 U778 ( .A0(n784), .A1(n265), .B0(n251), .B1(n1000), .Y(n297) );
  XNOR2XL U779 ( .A(n1067), .B(B[1]), .Y(n275) );
  XNOR2X1 U780 ( .A(n746), .B(n743), .Y(n299) );
  CMPR32X1 U781 ( .A(n262), .B(n261), .C(n260), .CO(n255), .S(n272) );
  OAI22XL U782 ( .A0(n801), .A1(n301), .B0(n799), .B1(n263), .Y(n280) );
  OAI22XL U783 ( .A0(n807), .A1(n274), .B0(n805), .B1(n264), .Y(n279) );
  XNOR2X1 U784 ( .A(n485), .B(n704), .Y(n283) );
  OAI22X1 U785 ( .A0(n1079), .A1(n267), .B0(n1101), .B1(n266), .Y(n281) );
  CMPR32X1 U786 ( .A(n273), .B(n272), .C(n271), .CO(n332), .S(n337) );
  XNOR2XL U787 ( .A(n1067), .B(B[0]), .Y(n276) );
  XNOR2XL U788 ( .A(n1049), .B(B[2]), .Y(n284) );
  CMPR22X1 U789 ( .A(n282), .B(n281), .CO(n278), .S(n935) );
  XNOR2X1 U790 ( .A(n437), .B(B[10]), .Y(n300) );
  OAI22XL U791 ( .A0(n792), .A1(n288), .B0(n791), .B1(n300), .Y(n943) );
  OAI22XL U792 ( .A0(n801), .A1(n289), .B0(n799), .B1(n302), .Y(n942) );
  CMPR32X1 U793 ( .A(n292), .B(n291), .C(n290), .CO(n328), .S(n331) );
  CMPR32X1 U794 ( .A(n295), .B(n294), .C(n293), .CO(n334), .S(n330) );
  XNOR2XL U795 ( .A(n746), .B(B[4]), .Y(n316) );
  OAI22XL U796 ( .A0(n1029), .A1(n316), .B0(n1030), .B1(n299), .Y(n315) );
  OAI22XL U797 ( .A0(n303), .A1(n302), .B0(n799), .B1(n301), .Y(n313) );
  CMPR32X1 U798 ( .A(n309), .B(n308), .C(n307), .CO(n329), .S(n966) );
  CMPR32X1 U799 ( .A(n312), .B(n311), .C(n310), .CO(n325), .S(n947) );
  ADDFHX1 U800 ( .A(n315), .B(n314), .CI(n313), .CO(n308), .S(n946) );
  CMPR22X1 U801 ( .A(n319), .B(n318), .CO(n949), .S(n939) );
  ADDFHX1 U802 ( .A(n322), .B(n321), .CI(n320), .CO(n934), .S(n948) );
  NAND2XL U803 ( .A(n926), .B(n925), .Y(mult_x_1_n313) );
  CMPR32X1 U804 ( .A(n328), .B(n327), .C(n326), .CO(n268), .S(n915) );
  CMPR32X1 U805 ( .A(n331), .B(n330), .C(n329), .CO(n914), .S(n335) );
  CMPR32X1 U806 ( .A(n337), .B(n336), .C(n335), .CO(n338), .S(n926) );
  NAND2X1 U807 ( .A(n644), .B(n341), .Y(n343) );
  INVXL U808 ( .A(n1005), .Y(n400) );
  NAND2XL U809 ( .A(n404), .B(n1004), .Y(n348) );
  NOR2XL U810 ( .A(n400), .B(n348), .Y(n350) );
  NAND2XL U811 ( .A(n430), .B(n350), .Y(n352) );
  OAI21XL U812 ( .A0(n1197), .A1(n1200), .B0(n1198), .Y(n504) );
  OAI21XL U813 ( .A0(n1193), .A1(n1196), .B0(n1194), .Y(n344) );
  OAI21XL U814 ( .A0(n1189), .A1(n1192), .B0(n1190), .Y(n1015) );
  INVXL U815 ( .A(n1015), .Y(n401) );
  OAI21XL U816 ( .A0(n401), .A1(n348), .B0(n347), .Y(n349) );
  AOI21XL U817 ( .A0(n470), .A1(n350), .B0(n349), .Y(n351) );
  OAI21XL U818 ( .A0(n1172), .A1(n352), .B0(n351), .Y(n354) );
  NOR2XL U819 ( .A(n400), .B(n1187), .Y(n356) );
  NAND2XL U820 ( .A(n430), .B(n356), .Y(n358) );
  OAI21XL U821 ( .A0(n401), .A1(n1187), .B0(n1188), .Y(n355) );
  AOI21XL U822 ( .A0(n470), .A1(n356), .B0(n355), .Y(n357) );
  OAI21XL U823 ( .A0(n1172), .A1(n358), .B0(n357), .Y(n360) );
  XNOR2X1 U824 ( .A(n360), .B(n359), .Y(PRODUCT[34]) );
  XNOR2X1 U825 ( .A(n1096), .B(B[16]), .Y(n410) );
  XNOR2X1 U826 ( .A(n365), .B(B[25]), .Y(n446) );
  BUFX3 U827 ( .A(B[26]), .Y(n1113) );
  OAI22XL U828 ( .A0(n1029), .A1(n407), .B0(n1030), .B1(n375), .Y(n380) );
  XNOR2X1 U829 ( .A(n757), .B(B[25]), .Y(n376) );
  INVXL U830 ( .A(n390), .Y(n379) );
  OAI22XL U831 ( .A0(n807), .A1(n409), .B0(n805), .B1(n376), .Y(n415) );
  OAI22XL U832 ( .A0(n1051), .A1(n408), .B0(n1076), .B1(n378), .Y(n413) );
  CMPR32X1 U833 ( .A(n381), .B(n380), .C(n379), .CO(n397), .S(n423) );
  CMPR32X1 U834 ( .A(n384), .B(n383), .C(n382), .CO(n427), .S(n422) );
  OAI22X1 U835 ( .A0(n1029), .A1(n387), .B0(n1030), .B1(n1027), .Y(n1045) );
  CMPR32X1 U836 ( .A(n391), .B(n390), .C(n389), .CO(n1037), .S(n396) );
  CMPR32X1 U837 ( .A(n394), .B(n393), .C(n392), .CO(n1036), .S(n395) );
  CMPR32X1 U838 ( .A(n397), .B(n396), .C(n395), .CO(n1023), .S(n426) );
  NOR2XL U839 ( .A(n399), .B(n398), .Y(mult_x_1_n162) );
  NAND2XL U840 ( .A(n399), .B(n398), .Y(mult_x_1_n163) );
  NAND2XL U841 ( .A(n430), .B(n1005), .Y(n403) );
  AOI21XL U842 ( .A0(n470), .A1(n1005), .B0(n1015), .Y(n402) );
  OAI21XL U843 ( .A0(n1172), .A1(n403), .B0(n402), .Y(n406) );
  XNOR2X2 U844 ( .A(n406), .B(n405), .Y(PRODUCT[33]) );
  INVXL U845 ( .A(n417), .Y(n443) );
  OAI22XL U846 ( .A0(n1118), .A1(n436), .B0(n1116), .B1(n410), .Y(n442) );
  OAI22XL U847 ( .A0(n1100), .A1(n447), .B0(n1101), .B1(n411), .Y(n441) );
  CMPR32X1 U848 ( .A(n415), .B(n414), .C(n413), .CO(n424), .S(n464) );
  CMPR32X1 U849 ( .A(n418), .B(n417), .C(n416), .CO(n382), .S(n463) );
  CMPR32X1 U850 ( .A(n427), .B(n426), .C(n425), .CO(n399), .S(n428) );
  NOR2XL U851 ( .A(n429), .B(n428), .Y(mult_x_1_n173) );
  NAND2XL U852 ( .A(n429), .B(n428), .Y(mult_x_1_n174) );
  NAND2XL U853 ( .A(n430), .B(n471), .Y(n432) );
  XNOR2X2 U854 ( .A(n435), .B(n434), .Y(PRODUCT[32]) );
  OAI22XL U855 ( .A0(n1118), .A1(n454), .B0(n1116), .B1(n436), .Y(n458) );
  XNOR2X1 U856 ( .A(n437), .B(B[25]), .Y(n490) );
  INVXL U857 ( .A(n438), .Y(n439) );
  CMPR32X1 U858 ( .A(n442), .B(n441), .C(n440), .CO(n419), .S(n478) );
  CMPR32X1 U859 ( .A(n445), .B(n444), .C(n443), .CO(n420), .S(n477) );
  XNOR2X1 U860 ( .A(n365), .B(B[24]), .Y(n452) );
  OAI22XL U861 ( .A0(n801), .A1(n452), .B0(n799), .B1(n446), .Y(n461) );
  OAI22XL U862 ( .A0(n1079), .A1(n480), .B0(n1101), .B1(n447), .Y(n460) );
  OAI22XL U863 ( .A0(n807), .A1(n453), .B0(n805), .B1(n448), .Y(n459) );
  OAI22XL U864 ( .A0(n1029), .A1(n455), .B0(n1030), .B1(n449), .Y(n489) );
  XNOR2X1 U865 ( .A(n1049), .B(B[18]), .Y(n451) );
  OAI22XL U866 ( .A0(n1075), .A1(n451), .B0(n1076), .B1(n450), .Y(n488) );
  XNOR2X1 U867 ( .A(n1049), .B(B[17]), .Y(n491) );
  OAI22X1 U868 ( .A0(n1051), .A1(n491), .B0(n1076), .B1(n451), .Y(n494) );
  XNOR2X1 U869 ( .A(n365), .B(B[23]), .Y(n492) );
  INVXL U870 ( .A(n457), .Y(n493) );
  CMPR32X1 U871 ( .A(n461), .B(n460), .C(n459), .CO(n500), .S(n515) );
  CMPR32X1 U872 ( .A(n467), .B(n466), .C(n465), .CO(n429), .S(n468) );
  NOR2XL U873 ( .A(n469), .B(n468), .Y(mult_x_1_n184) );
  NAND2XL U874 ( .A(n469), .B(n468), .Y(mult_x_1_n185) );
  XNOR2X2 U875 ( .A(n473), .B(n472), .Y(PRODUCT[31]) );
  CMPR32X1 U876 ( .A(n479), .B(n478), .C(n477), .CO(n476), .S(n514) );
  XNOR2X1 U877 ( .A(n1067), .B(n753), .Y(n482) );
  XNOR2X1 U878 ( .A(n757), .B(B[20]), .Y(n531) );
  OAI22X1 U879 ( .A0(n807), .A1(n531), .B0(n805), .B1(n481), .Y(n521) );
  OAI22XL U880 ( .A0(n1079), .A1(n525), .B0(n1101), .B1(n482), .Y(n520) );
  INVXL U881 ( .A(n518), .Y(n486) );
  CMPR32X1 U882 ( .A(n489), .B(n488), .C(n487), .CO(n499), .S(n539) );
  XNOR2X1 U883 ( .A(n437), .B(B[24]), .Y(n523) );
  XNOR2X1 U884 ( .A(n365), .B(B[22]), .Y(n529) );
  OAI22XL U885 ( .A0(n801), .A1(n529), .B0(n799), .B1(n492), .Y(n535) );
  NAND2XL U886 ( .A(n502), .B(n501), .Y(mult_x_1_n192) );
  INVXL U887 ( .A(n503), .Y(n544) );
  NAND2XL U888 ( .A(n503), .B(n545), .Y(n508) );
  INVXL U889 ( .A(n504), .Y(n505) );
  INVXL U890 ( .A(n505), .Y(n543) );
  AOI21XL U891 ( .A0(n543), .A1(n545), .B0(n506), .Y(n507) );
  NAND2X1 U892 ( .A(n509), .B(n1194), .Y(n510) );
  XNOR2X2 U893 ( .A(n511), .B(n510), .Y(PRODUCT[30]) );
  CMPR32X1 U894 ( .A(n517), .B(n516), .C(n515), .CO(n498), .S(n550) );
  XNOR2X1 U895 ( .A(n205), .B(B[25]), .Y(n556) );
  XNOR2X1 U896 ( .A(n1114), .B(n745), .Y(n558) );
  OAI22XL U897 ( .A0(n1029), .A1(n559), .B0(n1030), .B1(n522), .Y(n570) );
  OAI22X1 U898 ( .A0(n792), .A1(n560), .B0(n524), .B1(n523), .Y(n569) );
  XNOR2X1 U899 ( .A(n365), .B(B[21]), .Y(n565) );
  XNOR2X1 U900 ( .A(n1049), .B(n753), .Y(n566) );
  OAI22XL U901 ( .A0(n1051), .A1(n566), .B0(n1076), .B1(n530), .Y(n572) );
  CMPR32X1 U902 ( .A(n537), .B(n536), .C(n535), .CO(n553), .S(n585) );
  NOR2XL U903 ( .A(n542), .B(n541), .Y(mult_x_1_n202) );
  NAND2XL U904 ( .A(n542), .B(n541), .Y(mult_x_1_n203) );
  NAND2X1 U905 ( .A(n545), .B(n1196), .Y(n546) );
  CMPR32X1 U906 ( .A(n550), .B(n549), .C(n548), .CO(n541), .S(n578) );
  CMPR32X1 U907 ( .A(n553), .B(n552), .C(n551), .CO(n538), .S(n584) );
  XNOR2X1 U908 ( .A(n205), .B(B[24]), .Y(n590) );
  OAI22X1 U909 ( .A0(n557), .A1(n590), .B0(n556), .B1(n1000), .Y(n589) );
  XNOR2X1 U910 ( .A(n437), .B(B[22]), .Y(n593) );
  XNOR2X1 U911 ( .A(n365), .B(B[20]), .Y(n598) );
  OAI22XL U912 ( .A0(n1051), .A1(n599), .B0(n1076), .B1(n566), .Y(n605) );
  CMPR32X1 U913 ( .A(n573), .B(n572), .C(n571), .CO(n587), .S(n617) );
  NOR2XL U914 ( .A(n578), .B(n577), .Y(mult_x_1_n209) );
  NAND2XL U915 ( .A(n578), .B(n577), .Y(mult_x_1_n210) );
  INVXL U916 ( .A(n1197), .Y(n579) );
  CMPR32X1 U917 ( .A(n584), .B(n583), .C(n582), .CO(n577), .S(n611) );
  CMPR32X1 U918 ( .A(n587), .B(n586), .C(n585), .CO(n574), .S(n616) );
  CMPR22X1 U919 ( .A(n589), .B(n588), .CO(n596), .S(n629) );
  OAI22X1 U920 ( .A0(n784), .A1(n622), .B0(n590), .B1(n1000), .Y(n621) );
  XNOR2X1 U921 ( .A(n746), .B(n753), .Y(n624) );
  XNOR2X1 U922 ( .A(n437), .B(B[21]), .Y(n625) );
  CMPR32X1 U923 ( .A(n597), .B(n596), .C(n595), .CO(n609), .S(n640) );
  XNOR2X1 U924 ( .A(n365), .B(B[19]), .Y(n630) );
  XNOR2X1 U925 ( .A(n1049), .B(n756), .Y(n631) );
  OAI22XL U926 ( .A0(n716), .A1(n632), .B0(n805), .B1(n600), .Y(n636) );
  CMPR32X1 U927 ( .A(n606), .B(n605), .C(n604), .CO(n619), .S(n658) );
  NOR2XL U928 ( .A(n611), .B(n610), .Y(mult_x_1_n220) );
  NAND2XL U929 ( .A(n611), .B(n610), .Y(mult_x_1_n221) );
  INVXL U930 ( .A(n1199), .Y(n612) );
  NAND2XL U931 ( .A(n612), .B(n1200), .Y(n613) );
  CMPR32X1 U932 ( .A(n619), .B(n618), .C(n617), .CO(n607), .S(n657) );
  CMPR22X1 U933 ( .A(n621), .B(n620), .CO(n628), .S(n671) );
  XNOR2X1 U934 ( .A(n205), .B(B[22]), .Y(n663) );
  OAI22X1 U935 ( .A0(n784), .A1(n663), .B0(n622), .B1(n1000), .Y(n662) );
  OAI22XL U936 ( .A0(n1029), .A1(n665), .B0(n1030), .B1(n624), .Y(n677) );
  XNOR2X1 U937 ( .A(n437), .B(B[20]), .Y(n667) );
  OAI22X1 U938 ( .A0(n707), .A1(n667), .B0(n791), .B1(n625), .Y(n676) );
  XNOR2X1 U939 ( .A(A[13]), .B(B[10]), .Y(n668) );
  ADDFHX1 U940 ( .A(n635), .B(n634), .CI(n633), .CO(n627), .S(n697) );
  CMPR32X1 U941 ( .A(n641), .B(n640), .C(n639), .CO(n615), .S(n655) );
  NOR2XL U942 ( .A(n643), .B(n642), .Y(mult_x_1_n223) );
  NAND2XL U943 ( .A(n643), .B(n642), .Y(mult_x_1_n224) );
  INVXL U944 ( .A(n644), .Y(n686) );
  NOR2XL U945 ( .A(n686), .B(n1203), .Y(n649) );
  INVXL U946 ( .A(n647), .Y(n687) );
  OAI21XL U947 ( .A0(n687), .A1(n1203), .B0(n1204), .Y(n648) );
  AOI21XL U948 ( .A0(n6), .A1(n649), .B0(n648), .Y(n650) );
  OAI21XL U949 ( .A0(n26), .A1(n651), .B0(n650), .Y(n654) );
  CMPR32X1 U950 ( .A(n657), .B(n656), .C(n655), .CO(n642), .S(n685) );
  CMPR32X1 U951 ( .A(n660), .B(n659), .C(n658), .CO(n639), .S(n695) );
  CMPR22X1 U952 ( .A(n662), .B(n661), .CO(n670), .S(n712) );
  XNOR2X1 U953 ( .A(n205), .B(B[21]), .Y(n701) );
  XNOR2X1 U954 ( .A(n746), .B(n756), .Y(n705) );
  OAI22XL U955 ( .A0(n666), .A1(n705), .B0(n1030), .B1(n665), .Y(n719) );
  XNOR2X1 U956 ( .A(n437), .B(B[19]), .Y(n706) );
  OAI22X1 U957 ( .A0(n707), .A1(n706), .B0(n791), .B1(n667), .Y(n718) );
  XNOR2X1 U958 ( .A(A[13]), .B(B[9]), .Y(n709) );
  ADDFHX1 U959 ( .A(n677), .B(n676), .CI(n675), .CO(n669), .S(n738) );
  CMPR32X1 U960 ( .A(n683), .B(n682), .C(n681), .CO(n656), .S(n693) );
  NOR2XL U961 ( .A(n685), .B(n684), .Y(mult_x_1_n232) );
  NAND2XL U962 ( .A(n685), .B(n684), .Y(mult_x_1_n233) );
  AOI21XL U963 ( .A0(n6), .A1(n644), .B0(n647), .Y(n688) );
  OAI21XL U964 ( .A0(n26), .A1(n689), .B0(n688), .Y(n692) );
  XNOR2X2 U965 ( .A(n692), .B(n691), .Y(PRODUCT[25]) );
  CMPR32X1 U966 ( .A(n698), .B(n697), .C(n696), .CO(n681), .S(n736) );
  CMPR22X1 U967 ( .A(n700), .B(n699), .CO(n711), .S(n752) );
  XNOR2X1 U968 ( .A(n205), .B(B[20]), .Y(n742) );
  OAI22X1 U969 ( .A0(n784), .A1(n742), .B0(n701), .B1(n1000), .Y(n741) );
  OAI22X1 U970 ( .A0(n1118), .A1(n744), .B0(n1116), .B1(n703), .Y(n740) );
  XNOR2X1 U971 ( .A(n746), .B(n704), .Y(n747) );
  OAI22XL U972 ( .A0(n1029), .A1(n747), .B0(n1030), .B1(n705), .Y(n761) );
  XNOR2X1 U973 ( .A(n437), .B(B[18]), .Y(n748) );
  OAI22X1 U974 ( .A0(n707), .A1(n748), .B0(n791), .B1(n706), .Y(n760) );
  XNOR2X1 U975 ( .A(A[13]), .B(n708), .Y(n749) );
  NOR2XL U976 ( .A(n727), .B(n726), .Y(mult_x_1_n241) );
  OAI21XL U977 ( .A0(n26), .A1(n730), .B0(n729), .Y(n733) );
  NAND2X1 U978 ( .A(n731), .B(n1206), .Y(n732) );
  CMPR32X1 U979 ( .A(n736), .B(n735), .C(n734), .CO(n726), .S(n769) );
  CMPR32X1 U980 ( .A(n739), .B(n738), .C(n737), .CO(n723), .S(n776) );
  CMPR22X1 U981 ( .A(n741), .B(n740), .CO(n751), .S(n797) );
  XNOR2X1 U982 ( .A(n205), .B(B[19]), .Y(n782) );
  OAI22X1 U983 ( .A0(n784), .A1(n782), .B0(n742), .B1(n1000), .Y(n781) );
  OAI22X1 U984 ( .A0(n1118), .A1(n785), .B0(n1116), .B1(n744), .Y(n780) );
  XNOR2X1 U985 ( .A(n746), .B(n745), .Y(n788) );
  XNOR2X1 U986 ( .A(n437), .B(B[17]), .Y(n790) );
  OAI22X1 U987 ( .A0(n792), .A1(n790), .B0(n791), .B1(n748), .Y(n809) );
  XNOR2X1 U988 ( .A(A[13]), .B(B[7]), .Y(n793) );
  XNOR2X1 U989 ( .A(n365), .B(n753), .Y(n798) );
  OAI22XL U990 ( .A0(n801), .A1(n798), .B0(n799), .B1(n754), .Y(n813) );
  XNOR2X1 U991 ( .A(n1049), .B(B[9]), .Y(n802) );
  OAI22XL U992 ( .A0(n1051), .A1(n802), .B0(n1076), .B1(n755), .Y(n812) );
  CMPR32X1 U993 ( .A(n761), .B(n760), .C(n759), .CO(n750), .S(n831) );
  NOR2XL U994 ( .A(n769), .B(n768), .Y(mult_x_1_n252) );
  NAND2XL U995 ( .A(n769), .B(n768), .Y(mult_x_1_n253) );
  CMPR32X1 U996 ( .A(n776), .B(n775), .C(n774), .CO(n768), .S(n818) );
  CMPR32X1 U997 ( .A(n779), .B(n778), .C(n777), .CO(n765), .S(n829) );
  CMPR22X1 U998 ( .A(n781), .B(n780), .CO(n796), .S(n842) );
  OAI22X1 U999 ( .A0(n784), .A1(n783), .B0(n782), .B1(n1000), .Y(n834) );
  OAI22X1 U1000 ( .A0(n787), .A1(n786), .B0(n1116), .B1(n785), .Y(n833) );
  OAI22XL U1001 ( .A0(n801), .A1(n800), .B0(n799), .B1(n798), .Y(n851) );
  OAI22XL U1002 ( .A0(n1051), .A1(n803), .B0(n1076), .B1(n802), .Y(n850) );
  CMPR32X1 U1003 ( .A(n813), .B(n812), .C(n811), .CO(n832), .S(n865) );
  NOR2XL U1004 ( .A(n818), .B(n817), .Y(mult_x_1_n259) );
  NAND2XL U1005 ( .A(n818), .B(n817), .Y(mult_x_1_n260) );
  NAND2XL U1006 ( .A(n857), .B(n821), .Y(n823) );
  INVXL U1007 ( .A(n1212), .Y(n820) );
  AOI21XL U1008 ( .A0(n819), .A1(n821), .B0(n820), .Y(n822) );
  INVXL U1009 ( .A(n1209), .Y(n824) );
  CMPR32X1 U1010 ( .A(n829), .B(n828), .C(n827), .CO(n817), .S(n856) );
  CMPR32X1 U1011 ( .A(n832), .B(n831), .C(n830), .CO(n814), .S(n864) );
  CMPR22X1 U1012 ( .A(n834), .B(n833), .CO(n841), .S(n873) );
  CMPR22X1 U1013 ( .A(n836), .B(n835), .CO(n872), .S(n870) );
  CMPR32X1 U1014 ( .A(n845), .B(n844), .C(n843), .CO(n890), .S(n874) );
  CMPR32X1 U1015 ( .A(n851), .B(n850), .C(n849), .CO(n867), .S(n888) );
  CMPR32X1 U1016 ( .A(n854), .B(n853), .C(n852), .CO(n828), .S(n862) );
  NOR2XL U1017 ( .A(n856), .B(n855), .Y(mult_x_1_n270) );
  NAND2XL U1018 ( .A(n856), .B(n855), .Y(mult_x_1_n271) );
  NAND2X1 U1019 ( .A(n821), .B(n1212), .Y(n860) );
  CMPR32X1 U1020 ( .A(n870), .B(n869), .C(n868), .CO(n896), .S(n892) );
  CMPR32X1 U1021 ( .A(n873), .B(n872), .C(n871), .CO(n879), .S(n895) );
  CMPR32X1 U1022 ( .A(n876), .B(n875), .C(n874), .CO(n894), .S(n904) );
  CMPR32X1 U1023 ( .A(n879), .B(n878), .C(n877), .CO(n863), .S(n885) );
  NOR2XL U1024 ( .A(n881), .B(n880), .Y(mult_x_1_n277) );
  NAND2XL U1025 ( .A(n881), .B(n880), .Y(mult_x_1_n278) );
  OAI21X1 U1026 ( .A0(n26), .A1(n1215), .B0(n1216), .Y(n884) );
  NAND2X1 U1027 ( .A(n882), .B(n1214), .Y(n883) );
  XNOR2X2 U1028 ( .A(n884), .B(n883), .Y(PRODUCT[20]) );
  CMPR32X1 U1029 ( .A(n887), .B(n886), .C(n885), .CO(n880), .S(n898) );
  CMPR32X1 U1030 ( .A(n896), .B(n895), .C(n894), .CO(n886), .S(n899) );
  NOR2XL U1031 ( .A(n898), .B(n897), .Y(mult_x_1_n288) );
  NAND2XL U1032 ( .A(n898), .B(n897), .Y(mult_x_1_n289) );
  CMPR32X1 U1033 ( .A(n901), .B(n900), .C(n899), .CO(n897), .S(n906) );
  NOR2XL U1034 ( .A(n906), .B(n905), .Y(mult_x_1_n291) );
  NAND2XL U1035 ( .A(n906), .B(n905), .Y(mult_x_1_n292) );
  AOI21X2 U1036 ( .A0(n932), .A1(n1222), .B0(n1229), .Y(n920) );
  OAI21XL U1037 ( .A0(n920), .A1(n1220), .B0(n1221), .Y(n909) );
  INVXL U1038 ( .A(n1218), .Y(n907) );
  CMPR32X1 U1039 ( .A(n915), .B(n914), .C(n913), .CO(n921), .S(n339) );
  NOR2XL U1040 ( .A(mult_x_1_n302), .B(mult_x_1_n299), .Y(mult_x_1_n297) );
  NAND2XL U1041 ( .A(n917), .B(n916), .Y(mult_x_1_n300) );
  INVXL U1042 ( .A(n1220), .Y(n918) );
  NAND2X1 U1043 ( .A(n918), .B(n1221), .Y(n919) );
  NAND2XL U1044 ( .A(n922), .B(n921), .Y(mult_x_1_n303) );
  INVXL U1045 ( .A(n1225), .Y(n923) );
  INVXL U1046 ( .A(n927), .Y(n929) );
  NAND2XL U1047 ( .A(n929), .B(n928), .Y(mult_x_1_n78) );
  NAND2XL U1048 ( .A(n930), .B(n1225), .Y(n931) );
  XNOR2X1 U1049 ( .A(n932), .B(n931), .Y(PRODUCT[15]) );
  XNOR2X1 U1050 ( .A(n1231), .B(n1227), .Y(PRODUCT[14]) );
  CMPR32X1 U1051 ( .A(n935), .B(n934), .C(n933), .CO(n323), .S(n969) );
  CMPR32X1 U1052 ( .A(n938), .B(n937), .C(n936), .CO(n956), .S(n951) );
  CMPR32X1 U1053 ( .A(n941), .B(n940), .C(n939), .CO(n955), .S(n962) );
  CMPR32X1 U1054 ( .A(n944), .B(n943), .C(n942), .CO(n933), .S(n954) );
  CMPR32X1 U1055 ( .A(n947), .B(n946), .C(n945), .CO(n965), .S(n967) );
  CMPR32X1 U1056 ( .A(n950), .B(n949), .C(n948), .CO(n945), .S(n959) );
  CMPR32X1 U1057 ( .A(n953), .B(n952), .C(n951), .CO(n958), .S(n960) );
  CMPR32X1 U1058 ( .A(n959), .B(n958), .C(n957), .CO(n972), .S(n971) );
  NAND2XL U1059 ( .A(n980), .B(n983), .Y(n978) );
  NOR2XL U1060 ( .A(n978), .B(n1001), .Y(mult_x_1_n316) );
  INVXL U1061 ( .A(n981), .Y(n984) );
  NAND2XL U1062 ( .A(n973), .B(n972), .Y(n979) );
  INVXL U1063 ( .A(n979), .Y(n974) );
  OAI21XL U1064 ( .A0(n977), .A1(n1001), .B0(n1002), .Y(mult_x_1_n317) );
  XNOR2X1 U1065 ( .A(n1232), .B(n1228), .Y(PRODUCT[13]) );
  INVX1 U1066 ( .A(mult_x_1_n335), .Y(n985) );
  OAI21XL U1067 ( .A0(n985), .A1(n978), .B0(n977), .Y(mult_x_1_n320) );
  NAND2XL U1068 ( .A(n980), .B(n979), .Y(mult_x_1_n81) );
  NAND2XL U1069 ( .A(n983), .B(n981), .Y(n982) );
  XOR2X1 U1070 ( .A(n985), .B(n982), .Y(n1247) );
  OAI21XL U1071 ( .A0(n985), .A1(n963), .B0(n981), .Y(mult_x_1_n327) );
  NAND2XL U1072 ( .A(n36), .B(n988), .Y(n989) );
  XOR2X1 U1073 ( .A(n990), .B(n989), .Y(n1248) );
  NAND2XL U1074 ( .A(n5), .B(n991), .Y(n992) );
  INVXL U1075 ( .A(n994), .Y(n1128) );
  OAI21XL U1076 ( .A0(n1128), .A1(n1124), .B0(n1125), .Y(n999) );
  INVXL U1077 ( .A(n995), .Y(n997) );
  OAI21XL U1078 ( .A0(n1012), .A1(n1188), .B0(n1011), .Y(n1013) );
  AOI21XL U1079 ( .A0(n1015), .A1(n1014), .B0(n1013), .Y(n1016) );
  AOI21XL U1080 ( .A0(n1169), .A1(n1156), .B0(n1059), .Y(n1019) );
  OAI21XL U1081 ( .A0(n1172), .A1(n1020), .B0(n1019), .Y(n1022) );
  CMPR32X1 U1082 ( .A(n1035), .B(n1034), .C(n1033), .CO(n1052), .S(n1025) );
  CMPR32X1 U1083 ( .A(n1038), .B(n1037), .C(n1036), .CO(n1041), .S(n1024) );
  CMPR32X1 U1084 ( .A(n1046), .B(n1045), .C(n1044), .CO(n1087), .S(n1043) );
  OAI22X1 U1085 ( .A0(n1051), .A1(n1050), .B0(n1076), .B1(n1073), .Y(n1082) );
  CMPR32X1 U1086 ( .A(n1054), .B(n1053), .C(n1052), .CO(n1085), .S(n1042) );
  AOI21XL U1087 ( .A0(n1169), .A1(n1061), .B0(n1060), .Y(n1062) );
  OAI21XL U1088 ( .A0(n1172), .A1(n1063), .B0(n1062), .Y(n1066) );
  CMPR32X1 U1089 ( .A(n1071), .B(n1070), .C(n1069), .CO(n1089), .S(n1086) );
  OAI22X1 U1090 ( .A0(n1079), .A1(n1078), .B0(n1101), .B1(n1098), .Y(n1112) );
  CMPR32X1 U1091 ( .A(n1082), .B(n1081), .C(n1080), .CO(n1093), .S(n1088) );
  CMPR32X1 U1092 ( .A(n1087), .B(n1086), .C(n1085), .CO(n1092), .S(n1055) );
  CMPR32X1 U1093 ( .A(n1090), .B(n1089), .C(n1088), .CO(n1084), .S(n1091) );
  CMPR32X1 U1094 ( .A(n1095), .B(n1094), .C(n1093), .CO(n1103), .S(n1083) );
  OAI21XL U1095 ( .A0(n1105), .A1(n1177), .B0(n1178), .Y(n1165) );
  AOI21XL U1096 ( .A0(n1169), .A1(n1162), .B0(n1165), .Y(n1106) );
  OAI21XL U1097 ( .A0(n1172), .A1(n1107), .B0(n1106), .Y(n1109) );
  CMPR32X1 U1098 ( .A(n1112), .B(n1111), .C(n1110), .CO(n1121), .S(n1102) );
  XNOR2XL U1099 ( .A(n1114), .B(n1113), .Y(n1115) );
  XNOR2XL U1100 ( .A(n1161), .B(n1160), .Y(n1254) );
  AOI21XL U1101 ( .A0(n1169), .A1(n1168), .B0(n1167), .Y(n1170) );
  OAI21XL U1102 ( .A0(n1172), .A1(n1171), .B0(n1170), .Y(n1173) );
  XNOR2XL U1103 ( .A(n1173), .B(n1174), .Y(PRODUCT[40]) );
endmodule


module FFT2048_DW02_mult_2_stage_J1_12 ( A, B, TC, CLK, PRODUCT );
  input [25:0] A;
  input [16:0] B;
  output [42:0] PRODUCT;
  input TC, CLK;
  wire   n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         mult_x_1_n749, mult_x_1_n738, mult_x_1_n737, mult_x_1_n726,
         mult_x_1_n725, mult_x_1_n713, mult_x_1_n712, mult_x_1_n711,
         mult_x_1_n702, mult_x_1_n700, mult_x_1_n699, mult_x_1_n686,
         mult_x_1_n684, mult_x_1_n683, mult_x_1_n670, mult_x_1_n669,
         mult_x_1_n668, mult_x_1_n667, mult_x_1_n653, mult_x_1_n652,
         mult_x_1_n651, mult_x_1_n637, mult_x_1_n636, mult_x_1_n635,
         mult_x_1_n621, mult_x_1_n620, mult_x_1_n619, mult_x_1_n605,
         mult_x_1_n604, mult_x_1_n603, mult_x_1_n589, mult_x_1_n588,
         mult_x_1_n587, mult_x_1_n573, mult_x_1_n572, mult_x_1_n571,
         mult_x_1_n557, mult_x_1_n556, mult_x_1_n555, mult_x_1_n540,
         mult_x_1_n539, mult_x_1_n528, mult_x_1_n525, mult_x_1_n524,
         mult_x_1_n523, mult_x_1_n513, mult_x_1_n510, mult_x_1_n509,
         mult_x_1_n496, mult_x_1_n495, mult_x_1_n486, mult_x_1_n484,
         mult_x_1_n483, mult_x_1_n474, mult_x_1_n472, mult_x_1_n460,
         mult_x_1_n459, mult_x_1_n450, mult_x_1_n449, mult_x_1_n442,
         mult_x_1_n338, mult_x_1_n331, mult_x_1_n329, mult_x_1_n328,
         mult_x_1_n326, mult_x_1_n325, mult_x_1_n320, mult_x_1_n319,
         mult_x_1_n152, mult_x_1_n151, mult_x_1_n137, mult_x_1_n136,
         mult_x_1_n130, mult_x_1_n129, mult_x_1_n121, mult_x_1_n120,
         mult_x_1_n89, mult_x_1_n59, n5, n6, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299;

  DFFHQXL mult_x_1_clk_r_REG24_S1 ( .D(mult_x_1_n151), .CK(CLK), .Q(n1229) );
  DFFHQX1 mult_x_1_clk_r_REG66_S1 ( .D(mult_x_1_n737), .CK(CLK), .Q(n1297) );
  DFFHQX1 mult_x_1_clk_r_REG64_S1 ( .D(mult_x_1_n726), .CK(CLK), .Q(n1296) );
  DFFHQX1 mult_x_1_clk_r_REG63_S1 ( .D(mult_x_1_n725), .CK(CLK), .Q(n1295) );
  DFFHQX1 mult_x_1_clk_r_REG57_S1 ( .D(mult_x_1_n700), .CK(CLK), .Q(n1290) );
  DFFHQX4 mult_x_1_clk_r_REG53_S1 ( .D(mult_x_1_n686), .CK(CLK), .Q(n1288) );
  DFFHQX1 mult_x_1_clk_r_REG59_S1 ( .D(mult_x_1_n684), .CK(CLK), .Q(n1287) );
  DFFHQX2 mult_x_1_clk_r_REG58_S1 ( .D(mult_x_1_n683), .CK(CLK), .Q(n1286) );
  DFFHQX4 mult_x_1_clk_r_REG44_S1 ( .D(mult_x_1_n635), .CK(CLK), .Q(n1276) );
  DFFHQX2 mult_x_1_clk_r_REG41_S1 ( .D(mult_x_1_n619), .CK(CLK), .Q(n1273) );
  DFFHQX1 mult_x_1_clk_r_REG39_S1 ( .D(mult_x_1_n604), .CK(CLK), .Q(n1271) );
  DFFHQX2 mult_x_1_clk_r_REG38_S1 ( .D(mult_x_1_n603), .CK(CLK), .Q(n1270) );
  DFFHQX1 mult_x_1_clk_r_REG36_S1 ( .D(mult_x_1_n588), .CK(CLK), .Q(n1268) );
  DFFHQX4 mult_x_1_clk_r_REG32_S1 ( .D(mult_x_1_n571), .CK(CLK), .Q(n1264) );
  DFFHQX1 mult_x_1_clk_r_REG6_S1 ( .D(mult_x_1_n525), .CK(CLK), .Q(n1257) );
  DFFHQXL mult_x_1_clk_r_REG28_S1 ( .D(mult_x_1_n129), .CK(CLK), .Q(n1225) );
  DFFHQXL mult_x_1_clk_r_REG27_S1 ( .D(mult_x_1_n130), .CK(CLK), .Q(n1226) );
  DFFHQXL mult_x_1_clk_r_REG48_S1 ( .D(mult_x_1_n652), .CK(CLK), .Q(n1280) );
  DFFHQXL mult_x_1_clk_r_REG1_S1 ( .D(mult_x_1_n556), .CK(CLK), .Q(n1262) );
  DFFHQXL mult_x_1_clk_r_REG45_S1 ( .D(mult_x_1_n636), .CK(CLK), .Q(n1277) );
  DFFHQXL mult_x_1_clk_r_REG9_S1 ( .D(mult_x_1_n510), .CK(CLK), .Q(n1253) );
  DFFHQXL mult_x_1_clk_r_REG25_S1 ( .D(mult_x_1_n137), .CK(CLK), .Q(n1228) );
  DFFHQXL mult_x_1_clk_r_REG8_S1 ( .D(mult_x_1_n509), .CK(CLK), .Q(n1252) );
  DFFHQXL mult_x_1_clk_r_REG22_S1 ( .D(mult_x_1_n442), .CK(CLK), .Q(n1240) );
  DFFHQXL mult_x_1_clk_r_REG5_S1 ( .D(mult_x_1_n524), .CK(CLK), .Q(n1256) );
  DFFHQXL mult_x_1_clk_r_REG17_S1 ( .D(mult_x_1_n459), .CK(CLK), .Q(n1243) );
  DFFHQXL mult_x_1_clk_r_REG18_S1 ( .D(mult_x_1_n460), .CK(CLK), .Q(n1244) );
  DFFHQXL mult_x_1_clk_r_REG11_S1 ( .D(mult_x_1_n495), .CK(CLK), .Q(n1250) );
  DFFHQXL mult_x_1_clk_r_REG3_S1 ( .D(mult_x_1_n540), .CK(CLK), .Q(n1260) );
  DFFHQXL mult_x_1_clk_r_REG23_S1 ( .D(mult_x_1_n152), .CK(CLK), .Q(n1230) );
  DFFHQXL mult_x_1_clk_r_REG21_S1 ( .D(mult_x_1_n450), .CK(CLK), .Q(n1242) );
  DFFHQXL clk_r_REG80_S1 ( .D(n1312), .CK(CLK), .Q(PRODUCT[6]) );
  DFFHQXL mult_x_1_clk_r_REG26_S1 ( .D(mult_x_1_n136), .CK(CLK), .Q(n1227) );
  DFFHQX4 mult_x_1_clk_r_REG65_S1 ( .D(mult_x_1_n702), .CK(CLK), .Q(n1291) );
  DFFHQXL clk_r_REG77_S1 ( .D(n1310), .CK(CLK), .Q(PRODUCT[8]) );
  DFFHQXL clk_r_REG79_S1 ( .D(n1311), .CK(CLK), .Q(PRODUCT[7]) );
  DFFHQXL clk_r_REG81_S1 ( .D(n1313), .CK(CLK), .Q(PRODUCT[5]) );
  DFFHQXL clk_r_REG82_S1 ( .D(n1314), .CK(CLK), .Q(PRODUCT[4]) );
  DFFHQXL clk_r_REG83_S1 ( .D(n1315), .CK(CLK), .Q(PRODUCT[3]) );
  DFFHQXL clk_r_REG84_S1 ( .D(n1316), .CK(CLK), .Q(PRODUCT[2]) );
  DFFHQXL clk_r_REG85_S1 ( .D(n1317), .CK(CLK), .Q(PRODUCT[1]) );
  DFFHQXL clk_r_REG86_S1 ( .D(n1318), .CK(CLK), .Q(PRODUCT[0]) );
  DFFHQXL mult_x_1_clk_r_REG70_S1 ( .D(mult_x_1_n319), .CK(CLK), .Q(n1231) );
  DFFHQX1 mult_x_1_clk_r_REG68_S1 ( .D(mult_x_1_n749), .CK(CLK), .Q(n1299) );
  DFFHQX2 mult_x_1_clk_r_REG60_S1 ( .D(mult_x_1_n713), .CK(CLK), .Q(n1294) );
  DFFHQX2 mult_x_1_clk_r_REG56_S1 ( .D(mult_x_1_n699), .CK(CLK), .Q(n1289) );
  DFFHQX2 mult_x_1_clk_r_REG55_S1 ( .D(mult_x_1_n670), .CK(CLK), .Q(n1285) );
  DFFHQX2 mult_x_1_clk_r_REG54_S1 ( .D(mult_x_1_n669), .CK(CLK), .Q(n1284) );
  DFFHQX1 mult_x_1_clk_r_REG37_S1 ( .D(mult_x_1_n573), .CK(CLK), .Q(n1266) );
  DFFHQXL mult_x_1_clk_r_REG33_S1 ( .D(mult_x_1_n572), .CK(CLK), .Q(n1265) );
  DFFHQX1 mult_x_1_clk_r_REG34_S1 ( .D(mult_x_1_n557), .CK(CLK), .Q(n1263) );
  DFFHQX1 mult_x_1_clk_r_REG2_S1 ( .D(mult_x_1_n539), .CK(CLK), .Q(n1259) );
  DFFHQX1 mult_x_1_clk_r_REG7_S1 ( .D(mult_x_1_n528), .CK(CLK), .Q(n1258) );
  DFFHQX1 mult_x_1_clk_r_REG4_S1 ( .D(mult_x_1_n523), .CK(CLK), .Q(n1255) );
  DFFHQXL mult_x_1_clk_r_REG10_S1 ( .D(mult_x_1_n513), .CK(CLK), .Q(n1254) );
  DFFHQX1 mult_x_1_clk_r_REG12_S1 ( .D(mult_x_1_n496), .CK(CLK), .Q(n1251) );
  DFFHQXL mult_x_1_clk_r_REG16_S1 ( .D(mult_x_1_n472), .CK(CLK), .Q(n1245) );
  DFFHQXL mult_x_1_clk_r_REG20_S1 ( .D(mult_x_1_n449), .CK(CLK), .Q(n1241) );
  DFFHQXL mult_x_1_clk_r_REG78_S1 ( .D(mult_x_1_n338), .CK(CLK), .Q(n1239) );
  DFFHQXL mult_x_1_clk_r_REG76_S1 ( .D(mult_x_1_n331), .CK(CLK), .Q(n1238) );
  DFFHQXL mult_x_1_clk_r_REG75_S1 ( .D(mult_x_1_n89), .CK(CLK), .Q(n1237) );
  DFFHQXL mult_x_1_clk_r_REG73_S1 ( .D(mult_x_1_n329), .CK(CLK), .Q(n1236) );
  DFFHQXL mult_x_1_clk_r_REG71_S1 ( .D(mult_x_1_n326), .CK(CLK), .Q(n1234) );
  DFFHQXL mult_x_1_clk_r_REG72_S1 ( .D(mult_x_1_n325), .CK(CLK), .Q(n1233) );
  DFFHQXL mult_x_1_clk_r_REG69_S1 ( .D(mult_x_1_n320), .CK(CLK), .Q(n1232) );
  DFFHQXL mult_x_1_clk_r_REG29_S1 ( .D(mult_x_1_n121), .CK(CLK), .Q(n1224) );
  DFFHQXL mult_x_1_clk_r_REG31_S1 ( .D(mult_x_1_n59), .CK(CLK), .Q(n1222) );
  DFFHQXL mult_x_1_clk_r_REG15_S1 ( .D(mult_x_1_n486), .CK(CLK), .Q(n1249) );
  DFFHQXL mult_x_1_clk_r_REG19_S1 ( .D(mult_x_1_n474), .CK(CLK), .Q(n1246) );
  DFFHQXL mult_x_1_clk_r_REG30_S1 ( .D(mult_x_1_n120), .CK(CLK), .Q(n1223) );
  DFFHQXL mult_x_1_clk_r_REG61_S1 ( .D(mult_x_1_n711), .CK(CLK), .Q(n1292) );
  DFFHQX1 mult_x_1_clk_r_REG50_S1 ( .D(mult_x_1_n667), .CK(CLK), .Q(n1282) );
  DFFHQXL mult_x_1_clk_r_REG62_S1 ( .D(mult_x_1_n712), .CK(CLK), .Q(n1293) );
  DFFHQXL mult_x_1_clk_r_REG42_S1 ( .D(mult_x_1_n620), .CK(CLK), .Q(n1274) );
  DFFHQX1 mult_x_1_clk_r_REG74_S1 ( .D(mult_x_1_n328), .CK(CLK), .Q(n1235) );
  DFFHQXL mult_x_1_clk_r_REG13_S1 ( .D(mult_x_1_n483), .CK(CLK), .Q(n1247) );
  DFFHQX1 mult_x_1_clk_r_REG40_S1 ( .D(mult_x_1_n589), .CK(CLK), .Q(n1269) );
  DFFHQX1 mult_x_1_clk_r_REG43_S1 ( .D(mult_x_1_n605), .CK(CLK), .Q(n1272) );
  DFFHQX1 mult_x_1_clk_r_REG14_S1 ( .D(mult_x_1_n484), .CK(CLK), .Q(n1248) );
  DFFHQX1 mult_x_1_clk_r_REG35_S1 ( .D(mult_x_1_n587), .CK(CLK), .Q(n1267) );
  DFFHQX1 mult_x_1_clk_r_REG67_S1 ( .D(mult_x_1_n738), .CK(CLK), .Q(n1298) );
  DFFHQX1 mult_x_1_clk_r_REG47_S1 ( .D(mult_x_1_n651), .CK(CLK), .Q(n1279) );
  DFFHQX2 mult_x_1_clk_r_REG49_S1 ( .D(mult_x_1_n637), .CK(CLK), .Q(n1278) );
  DFFHQX2 mult_x_1_clk_r_REG52_S1 ( .D(mult_x_1_n653), .CK(CLK), .Q(n1281) );
  DFFHQX2 mult_x_1_clk_r_REG46_S1 ( .D(mult_x_1_n621), .CK(CLK), .Q(n1275) );
  DFFHQX1 mult_x_1_clk_r_REG0_S1 ( .D(mult_x_1_n555), .CK(CLK), .Q(n1261) );
  DFFHQX1 mult_x_1_clk_r_REG51_S1 ( .D(mult_x_1_n668), .CK(CLK), .Q(n1283) );
  CMPR32X1 U1 ( .A(n988), .B(n987), .C(n986), .CO(mult_x_1_n725), .S(
        mult_x_1_n726) );
  CMPR32X1 U2 ( .A(n1157), .B(n1156), .C(n1155), .CO(mult_x_1_n749), .S(n1083)
         );
  ADDFHX2 U3 ( .A(n513), .B(n512), .CI(n511), .CO(n506), .S(n532) );
  ADDFX2 U4 ( .A(n526), .B(n525), .CI(n524), .CO(n511), .S(n550) );
  BUFX3 U5 ( .A(n713), .Y(n1070) );
  BUFX3 U6 ( .A(n541), .Y(n5) );
  BUFX4 U7 ( .A(n935), .Y(n8) );
  BUFX3 U8 ( .A(n488), .Y(n9) );
  CLKINVX3 U9 ( .A(n979), .Y(n995) );
  NAND2X1 U10 ( .A(n97), .B(n406), .Y(n521) );
  XNOR2X2 U11 ( .A(B[14]), .B(B[13]), .Y(n541) );
  NAND2X1 U12 ( .A(n194), .B(n743), .Y(n949) );
  XNOR2X1 U13 ( .A(B[6]), .B(B[5]), .Y(n743) );
  OAI21XL U14 ( .A0(n1171), .A1(n22), .B0(n163), .Y(n165) );
  XNOR2X1 U15 ( .A(n302), .B(n301), .Y(PRODUCT[24]) );
  XNOR2X1 U16 ( .A(n268), .B(n267), .Y(PRODUCT[28]) );
  OAI21XL U17 ( .A0(n1171), .A1(n223), .B0(n222), .Y(n228) );
  OAI21X1 U18 ( .A0(n1171), .A1(n240), .B0(n239), .Y(n244) );
  NAND2X1 U19 ( .A(n126), .B(n322), .Y(n55) );
  OAI21X1 U20 ( .A0(n1119), .A1(n1122), .B0(n1123), .Y(n115) );
  NOR2X1 U21 ( .A(n120), .B(n119), .Y(n334) );
  NOR2X1 U22 ( .A(n294), .B(n298), .Y(n135) );
  NOR2X2 U23 ( .A(n129), .B(n130), .Y(n310) );
  ADDFHX1 U24 ( .A(n1284), .B(n1282), .CI(n1280), .CO(n123), .S(n122) );
  ADDFHX1 U25 ( .A(n1263), .B(n1261), .CI(n1260), .CO(n140), .S(n139) );
  ADDFHX1 U26 ( .A(n1266), .B(n1264), .CI(n1262), .CO(n138), .S(n137) );
  ADDFHX1 U27 ( .A(n1281), .B(n1279), .CI(n1277), .CO(n127), .S(n124) );
  ADDFHX2 U28 ( .A(n1272), .B(n1270), .CI(n1268), .CO(n133), .S(n132) );
  CMPR32X1 U29 ( .A(n1249), .B(n1248), .C(n1250), .CO(n153), .S(n151) );
  ADDFHX1 U30 ( .A(n1269), .B(n1267), .CI(n1265), .CO(n136), .S(n134) );
  NOR2X1 U31 ( .A(n143), .B(n142), .Y(n264) );
  OAI21X1 U32 ( .A0(n222), .A1(n162), .B0(n161), .Y(n1168) );
  XOR2XL U33 ( .A(n1121), .B(n1112), .Y(PRODUCT[14]) );
  XNOR2XL U34 ( .A(n993), .B(n945), .Y(n419) );
  XNOR2XL U35 ( .A(n993), .B(n1003), .Y(n418) );
  XNOR2XL U36 ( .A(n993), .B(n1066), .Y(n195) );
  XNOR2XL U37 ( .A(B[16]), .B(n950), .Y(n588) );
  XNOR2XL U38 ( .A(n1064), .B(n1000), .Y(n682) );
  XOR2XL U39 ( .A(n739), .B(n40), .Y(n39) );
  BUFX1 U40 ( .A(A[7]), .Y(n953) );
  XOR2XL U41 ( .A(B[11]), .B(B[10]), .Y(n30) );
  CLKINVX3 U42 ( .A(n472), .Y(n1001) );
  XNOR2XL U43 ( .A(n1067), .B(n874), .Y(n518) );
  XOR2XL U44 ( .A(n415), .B(n650), .Y(n484) );
  XNOR2XL U45 ( .A(n1064), .B(n928), .Y(n515) );
  XNOR2XL U46 ( .A(n993), .B(n739), .Y(n604) );
  XNOR2X2 U47 ( .A(B[10]), .B(B[9]), .Y(n640) );
  XOR2XL U48 ( .A(n415), .B(n709), .Y(n520) );
  XNOR2XL U49 ( .A(B[16]), .B(n974), .Y(n593) );
  XNOR2XL U50 ( .A(n993), .B(n850), .Y(n742) );
  BUFX3 U51 ( .A(n406), .Y(n6) );
  ADDFX2 U52 ( .A(n960), .B(n959), .CI(n958), .CO(mult_x_1_n713), .S(n961) );
  ADDFX2 U53 ( .A(n554), .B(n553), .CI(n552), .CO(mult_x_1_n495), .S(
        mult_x_1_n496) );
  INVX1 U54 ( .A(B[13]), .Y(n931) );
  NAND2XL U55 ( .A(n443), .B(n445), .Y(n37) );
  NAND2XL U56 ( .A(n638), .B(n639), .Y(n25) );
  OAI21XL U57 ( .A0(n638), .A1(n639), .B0(n637), .Y(n26) );
  INVX1 U58 ( .A(n444), .Y(n443) );
  OAI21XL U59 ( .A0(n756), .A1(n755), .B0(n754), .Y(n41) );
  INVX1 U60 ( .A(n38), .Y(n445) );
  INVXL U61 ( .A(n32), .Y(n31) );
  NOR2X1 U62 ( .A(n436), .B(n435), .Y(n38) );
  INVX1 U63 ( .A(n436), .Y(n36) );
  INVX1 U64 ( .A(n435), .Y(n35) );
  NOR2BXL U65 ( .AN(n747), .B(n34), .Y(n32) );
  OAI21XL U66 ( .A0(n6), .A1(n51), .B0(n50), .Y(n175) );
  NOR2X1 U67 ( .A(n14), .B(n13), .Y(n34) );
  OAI21XL U68 ( .A0(n889), .A1(n997), .B0(n28), .Y(n895) );
  OR2XL U69 ( .A(n821), .B(n640), .Y(n63) );
  NOR2BX1 U70 ( .AN(n1020), .B(n9), .Y(n880) );
  NAND2BXL U71 ( .AN(n64), .B(n29), .Y(n28) );
  NOR2X1 U72 ( .A(n9), .B(n540), .Y(n596) );
  NOR2X1 U73 ( .A(n9), .B(n593), .Y(n608) );
  NOR2X1 U74 ( .A(n9), .B(n81), .Y(n167) );
  OAI22X1 U75 ( .A0(n997), .A1(n101), .B0(n978), .B1(n73), .Y(n90) );
  NOR2X1 U76 ( .A(n9), .B(n453), .Y(n477) );
  NOR2BX1 U77 ( .AN(n1020), .B(n5), .Y(n913) );
  XOR2XL U78 ( .A(n415), .B(n680), .Y(n514) );
  XOR2XL U79 ( .A(n415), .B(n739), .Y(n559) );
  XNOR2X1 U80 ( .A(n228), .B(n227), .Y(PRODUCT[33]) );
  XNOR2X1 U81 ( .A(n1133), .B(n1132), .Y(PRODUCT[37]) );
  NOR2BX1 U82 ( .AN(n1020), .B(n6), .Y(n422) );
  XNOR2X1 U83 ( .A(B[1]), .B(A[24]), .Y(n589) );
  NAND2XL U84 ( .A(n21), .B(n19), .Y(n18) );
  XNOR2X1 U85 ( .A(n931), .B(n16), .Y(n714) );
  INVX2 U86 ( .A(n877), .Y(n482) );
  NAND2XL U87 ( .A(n21), .B(B[0]), .Y(n20) );
  XOR2X1 U88 ( .A(n415), .B(A[24]), .Y(n200) );
  XNOR2X1 U89 ( .A(B[1]), .B(n1063), .Y(n651) );
  XOR2XL U90 ( .A(n680), .B(B[1]), .Y(n21) );
  INVX1 U91 ( .A(n640), .Y(n29) );
  BUFX3 U92 ( .A(A[22]), .Y(n650) );
  NOR2BX1 U93 ( .AN(n1020), .B(n1033), .Y(n397) );
  CLKINVX3 U94 ( .A(B[9]), .Y(n415) );
  XOR2X1 U95 ( .A(n319), .B(n318), .Y(PRODUCT[21]) );
  INVX1 U96 ( .A(n1168), .Y(n163) );
  INVX2 U97 ( .A(n472), .Y(n954) );
  INVXL U98 ( .A(n950), .Y(n17) );
  INVX1 U99 ( .A(n1024), .Y(n19) );
  INVXL U100 ( .A(B[3]), .Y(n40) );
  INVX1 U101 ( .A(n1165), .Y(n22) );
  XOR2X1 U102 ( .A(n1151), .B(n1150), .Y(PRODUCT[13]) );
  NOR2X1 U103 ( .A(n223), .B(n162), .Y(n1165) );
  INVX1 U104 ( .A(n256), .Y(n287) );
  NAND2X1 U105 ( .A(n252), .B(n251), .Y(n253) );
  NAND2X1 U106 ( .A(n312), .B(n311), .Y(n313) );
  INVX1 U107 ( .A(n278), .Y(n290) );
  INVX1 U108 ( .A(n299), .Y(n24) );
  INVX1 U109 ( .A(n241), .Y(n11) );
  AOI21X1 U110 ( .A0(n1149), .A1(n1147), .B0(n110), .Y(n111) );
  NOR2X2 U111 ( .A(n134), .B(n133), .Y(n298) );
  ADDFHX1 U112 ( .A(n1258), .B(n1259), .CI(n1256), .CO(n142), .S(n141) );
  ADDFHX1 U113 ( .A(n1257), .B(n1255), .CI(n1253), .CO(n150), .S(n143) );
  NAND2XL U114 ( .A(n26), .B(n25), .Y(mult_x_1_n539) );
  OAI2BB1XL U115 ( .A0N(n755), .A1N(n756), .B0(n41), .Y(mult_x_1_n603) );
  XNOR2X1 U116 ( .A(n1118), .B(n1117), .Y(n1311) );
  NOR2X1 U117 ( .A(n36), .B(n35), .Y(n444) );
  ADDFHX1 U118 ( .A(n985), .B(n984), .CI(n983), .CO(n962), .S(n986) );
  OR2X2 U119 ( .A(n438), .B(n437), .Y(n1100) );
  XNOR2X1 U120 ( .A(n501), .B(n500), .Y(n46) );
  XOR2X1 U121 ( .A(n15), .B(n34), .Y(n758) );
  NOR2X1 U122 ( .A(n403), .B(n402), .Y(n1114) );
  ADDFHX1 U123 ( .A(n566), .B(n565), .CI(n564), .CO(n553), .S(n577) );
  OAI2BB1XL U124 ( .A0N(n942), .A1N(n8), .B0(n88), .Y(n1072) );
  NAND2X1 U125 ( .A(n401), .B(n400), .Y(n1176) );
  NOR2X1 U126 ( .A(n401), .B(n400), .Y(n1175) );
  INVX1 U127 ( .A(n98), .Y(n51) );
  NAND2BXL U128 ( .AN(n996), .B(n27), .Y(n60) );
  NOR2X1 U129 ( .A(n9), .B(n859), .Y(n1190) );
  NOR2X1 U130 ( .A(n9), .B(n801), .Y(n828) );
  NOR2X1 U131 ( .A(n9), .B(n772), .Y(n797) );
  NOR2X1 U132 ( .A(n9), .B(n831), .Y(n866) );
  NOR2X1 U133 ( .A(n9), .B(n489), .Y(n525) );
  OR2X2 U134 ( .A(n200), .B(n521), .Y(n50) );
  XNOR2X1 U135 ( .A(n1066), .B(n415), .Y(n98) );
  XNOR2XL U136 ( .A(B[13]), .B(n1063), .Y(n95) );
  INVX1 U137 ( .A(n997), .Y(n27) );
  OAI22XL U138 ( .A0(n1024), .A1(n770), .B0(n740), .B1(n769), .Y(n768) );
  XOR2X1 U139 ( .A(n415), .B(n953), .Y(n881) );
  XOR2X1 U140 ( .A(n415), .B(A[18]), .Y(n598) );
  XOR2X1 U141 ( .A(n415), .B(n799), .Y(n599) );
  XNOR2X1 U142 ( .A(n931), .B(n17), .Y(n745) );
  BUFX3 U143 ( .A(n640), .Y(n978) );
  BUFX3 U144 ( .A(B[11]), .Y(n72) );
  INVX1 U145 ( .A(n974), .Y(n16) );
  BUFX3 U146 ( .A(n956), .Y(n1033) );
  AOI21X1 U147 ( .A0(n342), .A1(n322), .B0(n321), .Y(n332) );
  INVX1 U148 ( .A(n288), .Y(n258) );
  BUFX2 U149 ( .A(A[4]), .Y(n992) );
  INVX1 U150 ( .A(n343), .Y(n1121) );
  INVX1 U151 ( .A(n160), .Y(n161) );
  NAND2BX1 U152 ( .AN(n233), .B(n11), .Y(n48) );
  AOI21X1 U153 ( .A0(n346), .A1(n344), .B0(n113), .Y(n1119) );
  INVXL U154 ( .A(n339), .Y(n10) );
  BUFX3 U155 ( .A(A[0]), .Y(n1020) );
  NOR2X1 U156 ( .A(n315), .B(n310), .Y(n293) );
  NOR2X1 U157 ( .A(n250), .B(n245), .Y(n229) );
  NOR2X1 U158 ( .A(n154), .B(n153), .Y(n230) );
  NAND2X1 U159 ( .A(n134), .B(n133), .Y(n299) );
  NAND2X1 U160 ( .A(n120), .B(n119), .Y(n335) );
  NAND2X1 U161 ( .A(n118), .B(n117), .Y(n340) );
  INVXL U162 ( .A(n1295), .Y(n52) );
  ADDFHX2 U163 ( .A(n1275), .B(n1273), .CI(n1271), .CO(n131), .S(n130) );
  NOR2X1 U164 ( .A(n1243), .B(n1242), .Y(n224) );
  XNOR2X1 U165 ( .A(n446), .B(n37), .Y(n1310) );
  INVXL U166 ( .A(n469), .Y(n57) );
  OAI2BB1X1 U167 ( .A0N(n501), .A1N(n500), .B0(n43), .Y(n469) );
  AOI21XL U168 ( .A0(n1100), .A1(n444), .B0(n439), .Y(n440) );
  NAND2XL U169 ( .A(n68), .B(n1043), .Y(n67) );
  OAI2BB1X1 U170 ( .A0N(n746), .A1N(n33), .B0(n31), .Y(n729) );
  XNOR2X1 U171 ( .A(n499), .B(n46), .Y(n502) );
  OR2XL U172 ( .A(n1079), .B(n1078), .Y(n1081) );
  OAI2BB1X1 U173 ( .A0N(n45), .A1N(n44), .B0(n499), .Y(n43) );
  INVX1 U174 ( .A(n756), .Y(n42) );
  ADDFHX2 U175 ( .A(n507), .B(n506), .CI(n505), .CO(n503), .S(mult_x_1_n472)
         );
  INVXL U176 ( .A(n500), .Y(n45) );
  ADDFHX1 U177 ( .A(n849), .B(n848), .CI(n847), .CO(mult_x_1_n653), .S(n845)
         );
  INVXL U178 ( .A(n501), .Y(n44) );
  NAND2BXL U179 ( .AN(n747), .B(n34), .Y(n33) );
  XNOR2X1 U180 ( .A(n747), .B(n746), .Y(n15) );
  OAI2BB1XL U181 ( .A0N(n743), .A1N(n1031), .B0(n196), .Y(n459) );
  OAI21XL U182 ( .A0(n997), .A1(n61), .B0(n59), .Y(n980) );
  OAI2BB1XL U183 ( .A0N(n6), .A1N(n521), .B0(n98), .Y(n174) );
  NAND2XL U184 ( .A(n516), .B(n70), .Y(n69) );
  OAI2BB1XL U185 ( .A0N(n1037), .A1N(n1039), .B0(n516), .Y(n570) );
  NOR2X1 U186 ( .A(n744), .B(n713), .Y(n14) );
  NOR2X1 U187 ( .A(n712), .B(n5), .Y(n13) );
  OAI22XL U188 ( .A0(n1031), .A1(n890), .B0(n1029), .B1(n863), .Y(n894) );
  OAI22XL U189 ( .A0(n1039), .A1(n731), .B0(n1037), .B1(n39), .Y(n734) );
  OAI21XL U190 ( .A0(n740), .A1(n1024), .B0(n20), .Y(n738) );
  OR2X2 U191 ( .A(n390), .B(n389), .Y(n388) );
  OAI22XL U192 ( .A0(n1039), .A1(n39), .B0(n1037), .B1(n672), .Y(n704) );
  OAI21XL U193 ( .A0(n681), .A1(n769), .B0(n18), .Y(n708) );
  OAI22X1 U194 ( .A0(n1027), .A1(n484), .B0(n6), .B1(n452), .Y(n479) );
  XNOR2X1 U195 ( .A(n165), .B(n164), .Y(PRODUCT[36]) );
  XOR2X1 U196 ( .A(n415), .B(n1063), .Y(n452) );
  BUFX3 U197 ( .A(B[16]), .Y(n1064) );
  XOR2X2 U198 ( .A(n249), .B(n248), .Y(PRODUCT[30]) );
  AND2XL U199 ( .A(n1221), .B(n1220), .Y(n1317) );
  OR2XL U200 ( .A(n1219), .B(n1218), .Y(n1221) );
  INVX2 U201 ( .A(B[11]), .Y(n979) );
  OR2XL U202 ( .A(n375), .B(n374), .Y(n1215) );
  INVX2 U203 ( .A(B[7]), .Y(n351) );
  BUFX2 U204 ( .A(A[19]), .Y(n739) );
  BUFX2 U205 ( .A(A[21]), .Y(n680) );
  INVXL U206 ( .A(n1000), .Y(n65) );
  INVXL U207 ( .A(n1037), .Y(n70) );
  INVXL U208 ( .A(n945), .Y(n62) );
  NAND2X1 U209 ( .A(n354), .B(n355), .Y(n952) );
  XOR2X1 U210 ( .A(B[2]), .B(B[3]), .Y(n354) );
  BUFX2 U211 ( .A(A[1]), .Y(n945) );
  XNOR2X1 U212 ( .A(B[2]), .B(B[1]), .Y(n355) );
  NAND2X1 U213 ( .A(n48), .B(n234), .Y(n47) );
  NAND2X1 U214 ( .A(n156), .B(n229), .Y(n223) );
  AND2X2 U215 ( .A(n247), .B(n246), .Y(n248) );
  BUFX2 U216 ( .A(A[2]), .Y(n1003) );
  OR2X2 U217 ( .A(n245), .B(n251), .Y(n49) );
  NAND2XL U218 ( .A(n226), .B(n225), .Y(n227) );
  AND2XL U219 ( .A(n1167), .B(n1172), .Y(n1161) );
  NAND2X1 U220 ( .A(n132), .B(n131), .Y(n306) );
  NAND2X2 U221 ( .A(n128), .B(n127), .Y(n316) );
  NAND2X2 U222 ( .A(n129), .B(n130), .Y(n311) );
  NOR2X1 U223 ( .A(n137), .B(n136), .Y(n278) );
  NOR2X1 U224 ( .A(n141), .B(n140), .Y(n255) );
  NOR2X1 U225 ( .A(n152), .B(n151), .Y(n245) );
  NAND2XL U226 ( .A(n219), .B(n218), .Y(n220) );
  ADDFHX2 U227 ( .A(n1291), .B(n1294), .CI(n1290), .CO(n117), .S(n114) );
  ADDFHX2 U228 ( .A(n1285), .B(n1286), .CI(n1283), .CO(n121), .S(n120) );
  ADDFHX2 U229 ( .A(n1288), .B(n1289), .CI(n1287), .CO(n119), .S(n118) );
  NAND2X1 U230 ( .A(n293), .B(n135), .Y(n256) );
  AOI21X1 U231 ( .A0(n1238), .A1(n109), .B0(n108), .Y(n1146) );
  XNOR2X1 U232 ( .A(n995), .B(n1003), .Y(n946) );
  NOR2X1 U233 ( .A(n233), .B(n230), .Y(n156) );
  OAI21XL U234 ( .A0(n222), .A1(n224), .B0(n225), .Y(n215) );
  XNOR2X1 U235 ( .A(n190), .B(n189), .Y(PRODUCT[35]) );
  XNOR2X1 U236 ( .A(n1067), .B(n953), .Y(n744) );
  XNOR2X1 U237 ( .A(n975), .B(n739), .Y(n770) );
  OAI22X1 U238 ( .A0(n8), .A1(n486), .B0(n942), .B1(n451), .Y(n480) );
  CLKINVX3 U239 ( .A(B[15]), .Y(n877) );
  BUFX2 U240 ( .A(n942), .Y(n12) );
  NAND2X4 U241 ( .A(n77), .B(n942), .Y(n935) );
  OAI22X1 U242 ( .A0(n8), .A1(n745), .B0(n12), .B1(n714), .Y(n746) );
  NOR2X1 U243 ( .A(n155), .B(n1244), .Y(n233) );
  XNOR3X2 U244 ( .A(n755), .B(n754), .C(n42), .Y(mult_x_1_n604) );
  OAI2BB1X2 U245 ( .A0N(n303), .A1N(n135), .B0(n23), .Y(n288) );
  AOI2BB1X2 U246 ( .A0N(n298), .A1N(n306), .B0(n24), .Y(n23) );
  OAI21X2 U247 ( .A0(n310), .A1(n316), .B0(n311), .Y(n303) );
  XOR3X2 U248 ( .A(n637), .B(n639), .C(n638), .Y(mult_x_1_n540) );
  NAND2X4 U249 ( .A(n640), .B(n30), .Y(n997) );
  XOR2X1 U250 ( .A(n979), .B(n947), .Y(n889) );
  AOI21X4 U251 ( .A0(n156), .A1(n238), .B0(n47), .Y(n222) );
  NAND2X2 U252 ( .A(n246), .B(n49), .Y(n238) );
  NAND2BX1 U253 ( .AN(n1293), .B(n52), .Y(n346) );
  AOI21X4 U254 ( .A0(n148), .A1(n257), .B0(n53), .Y(n1171) );
  OAI21X2 U255 ( .A0(n258), .A1(n147), .B0(n146), .Y(n53) );
  NAND2XL U256 ( .A(n254), .B(n145), .Y(n147) );
  OAI21X4 U257 ( .A0(n320), .A1(n55), .B0(n54), .Y(n257) );
  AOI21X2 U258 ( .A0(n321), .A1(n126), .B0(n125), .Y(n54) );
  AOI21X4 U259 ( .A0(n116), .A1(n343), .B0(n115), .Y(n320) );
  NOR2X1 U260 ( .A(n334), .B(n339), .Y(n322) );
  NOR2X1 U261 ( .A(n118), .B(n117), .Y(n339) );
  XNOR3X2 U262 ( .A(n58), .B(n468), .C(n469), .Y(mult_x_1_n450) );
  XOR2X2 U263 ( .A(n1171), .B(n253), .Y(PRODUCT[29]) );
  NAND2X2 U264 ( .A(n75), .B(n541), .Y(n713) );
  XOR2X1 U265 ( .A(B[14]), .B(B[15]), .Y(n75) );
  OAI21X2 U266 ( .A0(n1146), .A1(n112), .B0(n111), .Y(n343) );
  XNOR2X2 U267 ( .A(B[4]), .B(B[3]), .Y(n956) );
  INVX1 U268 ( .A(B[5]), .Y(n472) );
  INVXL U269 ( .A(n1227), .Y(n1128) );
  BUFX3 U270 ( .A(A[10]), .Y(n974) );
  AOI21XL U271 ( .A0(n185), .A1(n188), .B0(n157), .Y(n158) );
  BUFX3 U272 ( .A(A[25]), .Y(n1066) );
  BUFX3 U273 ( .A(A[23]), .Y(n1063) );
  OAI21XL U274 ( .A0(n282), .A1(n289), .B0(n283), .Y(n259) );
  NAND2XL U275 ( .A(n141), .B(n140), .Y(n274) );
  XNOR2XL U276 ( .A(n72), .B(A[24]), .Y(n101) );
  XNOR2XL U277 ( .A(n482), .B(n739), .Y(n172) );
  XNOR2XL U278 ( .A(n72), .B(n1063), .Y(n173) );
  BUFX2 U279 ( .A(A[20]), .Y(n709) );
  BUFX3 U280 ( .A(A[14]), .Y(n874) );
  BUFX3 U281 ( .A(A[15]), .Y(n850) );
  XNOR2XL U282 ( .A(n975), .B(A[16]), .Y(n851) );
  XNOR2XL U283 ( .A(n975), .B(n850), .Y(n875) );
  XNOR2XL U284 ( .A(n975), .B(A[13]), .Y(n929) );
  BUFX3 U285 ( .A(A[6]), .Y(n1000) );
  BUFX3 U286 ( .A(A[5]), .Y(n947) );
  BUFX3 U287 ( .A(A[9]), .Y(n950) );
  BUFX3 U288 ( .A(A[8]), .Y(n998) );
  CLKINVX3 U289 ( .A(n415), .Y(n1004) );
  XNOR2XL U290 ( .A(n1001), .B(n947), .Y(n1034) );
  XNOR2XL U291 ( .A(B[3]), .B(n953), .Y(n1038) );
  XNOR2XL U292 ( .A(n1004), .B(n945), .Y(n1026) );
  XNOR2XL U293 ( .A(n482), .B(n680), .Y(n80) );
  XNOR2XL U294 ( .A(n975), .B(n1003), .Y(n377) );
  XNOR2XL U295 ( .A(n975), .B(n992), .Y(n382) );
  XNOR2XL U296 ( .A(n975), .B(A[3]), .Y(n383) );
  XNOR2XL U297 ( .A(n1001), .B(n945), .Y(n368) );
  XNOR2XL U298 ( .A(B[3]), .B(n992), .Y(n358) );
  NAND2XL U299 ( .A(n1149), .B(n1148), .Y(n1150) );
  NAND2XL U300 ( .A(n346), .B(n345), .Y(n347) );
  NAND2XL U301 ( .A(n188), .B(n1230), .Y(n189) );
  OAI21XL U302 ( .A0(n1171), .A1(n187), .B0(n186), .Y(n190) );
  NAND2XL U303 ( .A(n1128), .B(n1228), .Y(n164) );
  BUFX3 U304 ( .A(A[17]), .Y(n799) );
  INVXL U305 ( .A(n1074), .Y(n83) );
  OAI22XL U306 ( .A0(n1070), .A1(n79), .B0(n5), .B1(n82), .Y(n85) );
  NOR2XL U307 ( .A(n9), .B(n76), .Y(n84) );
  XNOR2XL U308 ( .A(n1001), .B(n974), .Y(n925) );
  BUFX3 U309 ( .A(n1035), .Y(n957) );
  NAND2X1 U310 ( .A(n353), .B(n956), .Y(n1035) );
  XOR2XL U311 ( .A(B[4]), .B(B[5]), .Y(n353) );
  BUFX3 U312 ( .A(n952), .Y(n1039) );
  BUFX3 U313 ( .A(n743), .Y(n1029) );
  NAND2BXL U314 ( .AN(n1020), .B(n995), .Y(n977) );
  NOR2BXL U315 ( .AN(n1020), .B(n942), .Y(n982) );
  XNOR2XL U316 ( .A(n975), .B(n945), .Y(n372) );
  NOR2XL U317 ( .A(n9), .B(n86), .Y(n1073) );
  INVXL U318 ( .A(n87), .Y(n88) );
  OR2X2 U319 ( .A(n1045), .B(n1044), .Y(n68) );
  NAND2XL U320 ( .A(n1149), .B(n1186), .Y(n112) );
  XNOR2XL U321 ( .A(n995), .B(n1066), .Y(n73) );
  XNOR2XL U322 ( .A(n1185), .B(n1184), .Y(PRODUCT[11]) );
  NAND2XL U323 ( .A(n1183), .B(n1234), .Y(n1184) );
  XOR2XL U324 ( .A(n1182), .B(n1181), .Y(PRODUCT[10]) );
  NAND2XL U325 ( .A(n124), .B(n123), .Y(n324) );
  INVXL U326 ( .A(n323), .Y(n325) );
  NOR2XL U327 ( .A(n1227), .B(n1225), .Y(n1167) );
  INVXL U328 ( .A(n73), .Y(n74) );
  XNOR2XL U329 ( .A(B[3]), .B(n947), .Y(n408) );
  XNOR2XL U330 ( .A(n1001), .B(A[3]), .Y(n410) );
  XNOR2XL U331 ( .A(n1004), .B(n1020), .Y(n407) );
  XNOR2XL U332 ( .A(n1001), .B(n992), .Y(n409) );
  XNOR2XL U333 ( .A(B[3]), .B(n1000), .Y(n413) );
  XNOR2XL U334 ( .A(n482), .B(A[18]), .Y(n201) );
  XNOR2X1 U335 ( .A(B[1]), .B(n1066), .Y(n587) );
  XNOR2XL U336 ( .A(n995), .B(n874), .Y(n622) );
  XNOR2XL U337 ( .A(B[3]), .B(n650), .Y(n623) );
  XNOR2XL U338 ( .A(n954), .B(n709), .Y(n624) );
  XNOR2XL U339 ( .A(n995), .B(A[13]), .Y(n641) );
  XNOR2XL U340 ( .A(B[3]), .B(n680), .Y(n642) );
  XNOR2XL U341 ( .A(n954), .B(n739), .Y(n643) );
  XNOR2XL U342 ( .A(n995), .B(n950), .Y(n760) );
  XNOR2XL U343 ( .A(B[3]), .B(n799), .Y(n761) );
  XNOR2XL U344 ( .A(n1001), .B(n850), .Y(n762) );
  XNOR2XL U345 ( .A(n1067), .B(n945), .Y(n882) );
  XNOR2XL U346 ( .A(n1067), .B(n1020), .Y(n883) );
  BUFX3 U347 ( .A(A[11]), .Y(n943) );
  XNOR2XL U348 ( .A(n1004), .B(n1000), .Y(n914) );
  XNOR2XL U349 ( .A(B[3]), .B(n943), .Y(n918) );
  NAND2BXL U350 ( .AN(n1020), .B(n1004), .Y(n414) );
  XNOR2XL U351 ( .A(B[3]), .B(n945), .Y(n385) );
  OAI22XL U352 ( .A0(n1024), .A1(n417), .B0(n416), .B1(n1021), .Y(n421) );
  NAND2BXL U353 ( .AN(n1020), .B(n993), .Y(n350) );
  XNOR2XL U354 ( .A(n1188), .B(n1187), .Y(PRODUCT[12]) );
  NAND2XL U355 ( .A(n1186), .B(n1232), .Y(n1187) );
  NAND2XL U356 ( .A(n284), .B(n283), .Y(n285) );
  OAI21XL U357 ( .A0(n319), .A1(n281), .B0(n280), .Y(n286) );
  NAND2XL U358 ( .A(n275), .B(n274), .Y(n276) );
  OAI21XL U359 ( .A0(n319), .A1(n273), .B0(n272), .Y(n277) );
  INVXL U360 ( .A(n1159), .Y(n1160) );
  AOI21XL U361 ( .A0(n1166), .A1(n1172), .B0(n1158), .Y(n1159) );
  INVXL U362 ( .A(n1224), .Y(n1158) );
  NAND2XL U363 ( .A(n1165), .B(n1167), .Y(n1170) );
  INVXL U364 ( .A(n1223), .Y(n1172) );
  NOR2X1 U365 ( .A(n256), .B(n147), .Y(n148) );
  INVXL U366 ( .A(n1228), .Y(n1127) );
  NAND2XL U367 ( .A(n1165), .B(n1128), .Y(n1130) );
  INVXL U368 ( .A(n1225), .Y(n1131) );
  XNOR2XL U369 ( .A(B[3]), .B(n874), .Y(n852) );
  OAI22XL U370 ( .A0(n997), .A1(n173), .B0(n978), .B1(n101), .Y(n177) );
  XNOR2XL U371 ( .A(n482), .B(n799), .Y(n454) );
  XNOR2XL U372 ( .A(n72), .B(A[18]), .Y(n523) );
  XNOR2X1 U373 ( .A(n954), .B(n1066), .Y(n473) );
  OAI22X1 U374 ( .A0(n957), .A1(n517), .B0(n1033), .B1(n473), .Y(n494) );
  OAI22XL U375 ( .A0(n1070), .A1(n80), .B0(n5), .B1(n79), .Y(n93) );
  OAI22XL U376 ( .A0(n8), .A1(n95), .B0(n942), .B1(n78), .Y(n94) );
  XNOR2XL U377 ( .A(n72), .B(n680), .Y(n455) );
  XNOR2XL U378 ( .A(n72), .B(n650), .Y(n450) );
  NOR2XL U379 ( .A(n9), .B(n193), .Y(n461) );
  XNOR2XL U380 ( .A(n482), .B(A[16]), .Y(n483) );
  XNOR2XL U381 ( .A(n482), .B(n850), .Y(n491) );
  XNOR2XL U382 ( .A(n72), .B(n709), .Y(n485) );
  XNOR2XL U383 ( .A(n72), .B(n739), .Y(n492) );
  OAI22XL U384 ( .A0(n1031), .A1(n539), .B0(n743), .B1(n519), .Y(n543) );
  BUFX3 U385 ( .A(A[12]), .Y(n928) );
  XNOR2XL U386 ( .A(B[3]), .B(A[24]), .Y(n555) );
  XNOR2XL U387 ( .A(B[3]), .B(n1063), .Y(n583) );
  XNOR2XL U388 ( .A(n72), .B(n850), .Y(n582) );
  XNOR2XL U389 ( .A(n954), .B(n650), .Y(n591) );
  XNOR2XL U390 ( .A(n954), .B(n1063), .Y(n558) );
  OAI21XL U391 ( .A0(n555), .A1(n1039), .B0(n69), .Y(n571) );
  OAI22XL U392 ( .A0(n1070), .A1(n605), .B0(n5), .B1(n563), .Y(n602) );
  OAI22XL U393 ( .A0(n1031), .A1(n604), .B0(n743), .B1(n562), .Y(n603) );
  XNOR2XL U394 ( .A(n72), .B(A[16]), .Y(n561) );
  XNOR2XL U395 ( .A(n72), .B(n799), .Y(n560) );
  XNOR2XL U396 ( .A(n1004), .B(A[16]), .Y(n647) );
  XNOR2XL U397 ( .A(n1004), .B(n850), .Y(n677) );
  XNOR2XL U398 ( .A(n1067), .B(n974), .Y(n654) );
  XNOR2XL U399 ( .A(n1004), .B(n874), .Y(n706) );
  XNOR2XL U400 ( .A(n1004), .B(A[13]), .Y(n736) );
  XNOR2XL U401 ( .A(n1004), .B(n928), .Y(n766) );
  XNOR2XL U402 ( .A(n1004), .B(n943), .Y(n796) );
  XNOR2XL U403 ( .A(n1067), .B(n1000), .Y(n774) );
  XNOR2XL U404 ( .A(n1004), .B(n974), .Y(n823) );
  XNOR2XL U405 ( .A(n1001), .B(n874), .Y(n824) );
  XNOR2XL U406 ( .A(n1001), .B(A[13]), .Y(n825) );
  XNOR2XL U407 ( .A(n995), .B(n953), .Y(n821) );
  XNOR2XL U408 ( .A(n995), .B(n998), .Y(n791) );
  XNOR2XL U409 ( .A(B[3]), .B(A[16]), .Y(n792) );
  XNOR2XL U410 ( .A(n1067), .B(n992), .Y(n804) );
  XNOR2XL U411 ( .A(n1004), .B(n950), .Y(n864) );
  XNOR2XL U412 ( .A(n1004), .B(n998), .Y(n865) );
  OAI22XL U413 ( .A0(n1024), .A1(n851), .B0(n830), .B1(n1021), .Y(n867) );
  NAND2BXL U414 ( .AN(n1020), .B(B[16]), .Y(n831) );
  XNOR2XL U415 ( .A(n1001), .B(n943), .Y(n906) );
  NAND2BXL U416 ( .AN(n1020), .B(n1067), .Y(n876) );
  XNOR2XL U417 ( .A(B[3]), .B(A[13]), .Y(n888) );
  XNOR2XL U418 ( .A(B[3]), .B(n928), .Y(n917) );
  OAI22XL U419 ( .A0(n1024), .A1(n929), .B0(n909), .B1(n1021), .Y(n912) );
  OAI22XL U420 ( .A0(n957), .A1(n926), .B0(n1033), .B1(n925), .Y(n939) );
  OAI22XL U421 ( .A0(n949), .A1(n932), .B0(n1029), .B1(n927), .Y(n938) );
  OAI22XL U422 ( .A0(n1039), .A1(n1038), .B0(n1037), .B1(n1036), .Y(n1089) );
  OAI22XL U423 ( .A0(n1035), .A1(n1034), .B0(n1033), .B1(n1032), .Y(n1090) );
  OAI22XL U424 ( .A0(n1031), .A1(n1030), .B0(n1029), .B1(n1028), .Y(n1091) );
  NOR2BXL U425 ( .AN(n1020), .B(n640), .Y(n1053) );
  OAI22XL U426 ( .A0(n1024), .A1(n1023), .B0(n1022), .B1(n1021), .Y(n1052) );
  OAI22XL U427 ( .A0(n1027), .A1(n1026), .B0(n6), .B1(n1025), .Y(n1051) );
  INVXL U428 ( .A(B[1]), .Y(n349) );
  BUFX3 U429 ( .A(n771), .Y(n1024) );
  NOR2BXL U430 ( .AN(n1020), .B(n1037), .Y(n374) );
  OAI22XL U431 ( .A0(n1024), .A1(n372), .B0(n377), .B1(n1021), .Y(n375) );
  OAI22XL U432 ( .A0(n1039), .A1(n384), .B0(n1037), .B1(n367), .Y(n394) );
  OAI22XL U433 ( .A0(n957), .A1(n369), .B0(n1033), .B1(n368), .Y(n393) );
  XNOR2XL U434 ( .A(n1001), .B(n1020), .Y(n369) );
  OAI22XL U435 ( .A0(n1039), .A1(n367), .B0(n1037), .B1(n358), .Y(n366) );
  ADDFX2 U436 ( .A(n431), .B(n430), .CI(n429), .CO(n437), .S(n436) );
  INVXL U437 ( .A(n1071), .Y(n1076) );
  OAI22XL U438 ( .A0(n1070), .A1(n1069), .B0(n5), .B1(n1068), .Y(n1071) );
  XNOR2XL U439 ( .A(n1067), .B(n1066), .Y(n1068) );
  NOR2XL U440 ( .A(n9), .B(n1065), .Y(n1077) );
  OAI22XL U441 ( .A0(n1070), .A1(n82), .B0(n5), .B1(n1069), .Y(n1062) );
  NAND2XL U442 ( .A(n438), .B(n437), .Y(n1101) );
  ADDFX2 U443 ( .A(n870), .B(n869), .CI(n868), .CO(n846), .S(n871) );
  OAI22XL U444 ( .A0(n957), .A1(n1002), .B0(n1033), .B1(n955), .Y(n1008) );
  OAI22XL U445 ( .A0(n952), .A1(n999), .B0(n1037), .B1(n951), .Y(n1009) );
  OAI22XL U446 ( .A0(n1035), .A1(n1032), .B0(n1033), .B1(n1002), .Y(n1048) );
  OAI22XL U447 ( .A0(n1039), .A1(n1036), .B0(n1037), .B1(n999), .Y(n1040) );
  OAI22XL U448 ( .A0(n1031), .A1(n1028), .B0(n1029), .B1(n994), .Y(n1042) );
  OAI21XL U449 ( .A0(n640), .A1(n61), .B0(n60), .Y(n1041) );
  OAI22XL U450 ( .A0(n1027), .A1(n1005), .B0(n6), .B1(n973), .Y(n1019) );
  OAI22XL U451 ( .A0(n1024), .A1(n1020), .B0(n372), .B1(n1021), .Y(n1219) );
  NAND2XL U452 ( .A(n373), .B(n1024), .Y(n1218) );
  NAND2BXL U453 ( .AN(n1020), .B(n975), .Y(n373) );
  NAND2XL U454 ( .A(n1219), .B(n1218), .Y(n1220) );
  NAND2XL U455 ( .A(n375), .B(n374), .Y(n1214) );
  INVXL U456 ( .A(n1220), .Y(n1216) );
  INVXL U457 ( .A(n1113), .Y(n1178) );
  NAND2XL U458 ( .A(n1083), .B(n1082), .Y(mult_x_1_n320) );
  INVXL U459 ( .A(n1238), .Y(n1182) );
  NOR2X1 U460 ( .A(n132), .B(n131), .Y(n294) );
  NOR2XL U461 ( .A(n255), .B(n264), .Y(n145) );
  XNOR2XL U462 ( .A(n975), .B(n998), .Y(n416) );
  XNOR2XL U463 ( .A(B[1]), .B(n953), .Y(n417) );
  INVXL U464 ( .A(n1231), .Y(n1186) );
  NAND2X1 U465 ( .A(n114), .B(n1292), .Y(n1123) );
  INVXL U466 ( .A(n340), .Y(n333) );
  INVXL U467 ( .A(n334), .Y(n336) );
  INVXL U468 ( .A(n294), .Y(n307) );
  INVXL U469 ( .A(n298), .Y(n300) );
  AOI21XL U470 ( .A0(n288), .A1(n290), .B0(n279), .Y(n280) );
  INVXL U471 ( .A(n282), .Y(n284) );
  AOI21XL U472 ( .A0(n288), .A1(n261), .B0(n260), .Y(n262) );
  INVXL U473 ( .A(n264), .Y(n266) );
  INVXL U474 ( .A(n233), .Y(n235) );
  INVXL U475 ( .A(n224), .Y(n226) );
  NAND2XL U476 ( .A(n1241), .B(n1240), .Y(n218) );
  INVXL U477 ( .A(n218), .Y(n185) );
  INVXL U478 ( .A(n1230), .Y(n157) );
  NAND2XL U479 ( .A(n219), .B(n188), .Y(n159) );
  NAND2XL U480 ( .A(n1243), .B(n1242), .Y(n225) );
  INVXL U481 ( .A(n1229), .Y(n188) );
  XNOR2XL U482 ( .A(n1064), .B(A[18]), .Y(n96) );
  XNOR2XL U483 ( .A(B[13]), .B(A[24]), .Y(n78) );
  XNOR2XL U484 ( .A(n1064), .B(A[16]), .Y(n193) );
  XNOR2XL U485 ( .A(B[1]), .B(n650), .Y(n681) );
  XNOR2XL U486 ( .A(n995), .B(n928), .Y(n671) );
  XNOR2XL U487 ( .A(B[3]), .B(n709), .Y(n672) );
  XNOR2XL U488 ( .A(n954), .B(A[18]), .Y(n673) );
  XNOR2XL U489 ( .A(n995), .B(n943), .Y(n701) );
  XNOR2XL U490 ( .A(n954), .B(n799), .Y(n702) );
  XNOR2XL U491 ( .A(B[1]), .B(n709), .Y(n740) );
  XNOR2XL U492 ( .A(n995), .B(n974), .Y(n730) );
  XNOR2XL U493 ( .A(B[3]), .B(A[18]), .Y(n731) );
  XNOR2XL U494 ( .A(n1001), .B(A[16]), .Y(n732) );
  XNOR2XL U495 ( .A(n975), .B(A[18]), .Y(n800) );
  XNOR2XL U496 ( .A(B[1]), .B(n799), .Y(n830) );
  XNOR2XL U497 ( .A(n975), .B(n874), .Y(n909) );
  XNOR2XL U498 ( .A(n1001), .B(n950), .Y(n926) );
  XNOR2XL U499 ( .A(n975), .B(n943), .Y(n976) );
  XNOR2XL U500 ( .A(n975), .B(n974), .Y(n1022) );
  XNOR2XL U501 ( .A(n975), .B(n950), .Y(n1023) );
  XNOR2XL U502 ( .A(B[3]), .B(A[3]), .Y(n367) );
  NAND2BXL U503 ( .AN(n1020), .B(n1001), .Y(n360) );
  NOR2BXL U504 ( .AN(n1020), .B(n1029), .Y(n363) );
  OAI22XL U505 ( .A0(n1035), .A1(n357), .B0(n1033), .B1(n410), .Y(n423) );
  OAI22X1 U506 ( .A0(n949), .A1(n356), .B0(n1029), .B1(n419), .Y(n424) );
  OAI22XL U507 ( .A0(n1039), .A1(n358), .B0(n1037), .B1(n408), .Y(n425) );
  XOR2X1 U508 ( .A(n338), .B(n337), .Y(PRODUCT[18]) );
  NAND2XL U509 ( .A(n336), .B(n335), .Y(n337) );
  AOI21X1 U510 ( .A0(n342), .A1(n10), .B0(n333), .Y(n338) );
  XOR2X1 U511 ( .A(n332), .B(n331), .Y(PRODUCT[19]) );
  XNOR2X1 U512 ( .A(n327), .B(n326), .Y(PRODUCT[20]) );
  NAND2XL U513 ( .A(n325), .B(n324), .Y(n326) );
  OAI21XL U514 ( .A0(n332), .A1(n328), .B0(n329), .Y(n327) );
  NAND2XL U515 ( .A(n317), .B(n316), .Y(n318) );
  XNOR2X1 U516 ( .A(n237), .B(n236), .Y(PRODUCT[32]) );
  NAND2XL U517 ( .A(n235), .B(n234), .Y(n236) );
  OAI21X1 U518 ( .A0(n1171), .A1(n232), .B0(n231), .Y(n237) );
  XNOR2X1 U519 ( .A(B[13]), .B(n1066), .Y(n87) );
  XNOR2XL U520 ( .A(n482), .B(n1063), .Y(n82) );
  NOR2XL U521 ( .A(n9), .B(n71), .Y(n91) );
  OAI2BB1XL U522 ( .A0N(n978), .A1N(n997), .B0(n74), .Y(n89) );
  XNOR2XL U523 ( .A(n1064), .B(n709), .Y(n71) );
  OAI22XL U524 ( .A0(n952), .A1(n408), .B0(n1037), .B1(n413), .Y(n428) );
  OAI22XL U525 ( .A0(n957), .A1(n410), .B0(n1033), .B1(n409), .Y(n427) );
  OAI22XL U526 ( .A0(n957), .A1(n409), .B0(n956), .B1(n1034), .Y(n1054) );
  OAI22XL U527 ( .A0(n1031), .A1(n418), .B0(n1029), .B1(n1030), .Y(n1056) );
  OAI22XL U528 ( .A0(n1027), .A1(n407), .B0(n6), .B1(n1026), .Y(n1055) );
  OAI22XL U529 ( .A0(n1039), .A1(n413), .B0(n1037), .B1(n1038), .Y(n1094) );
  OAI22XL U530 ( .A0(n997), .A1(n450), .B0(n978), .B1(n173), .Y(n204) );
  OAI22XL U531 ( .A0(n1070), .A1(n201), .B0(n5), .B1(n172), .Y(n205) );
  OAI22XL U532 ( .A0(n8), .A1(n451), .B0(n942), .B1(n202), .Y(n456) );
  OAI22XL U533 ( .A0(n521), .A1(n452), .B0(n6), .B1(n200), .Y(n458) );
  OAI22XL U534 ( .A0(n997), .A1(n560), .B0(n978), .B1(n523), .Y(n546) );
  OAI22XL U535 ( .A0(n521), .A1(n559), .B0(n6), .B1(n520), .Y(n548) );
  OAI22XL U536 ( .A0(n8), .A1(n522), .B0(n942), .B1(n487), .Y(n526) );
  XOR2XL U537 ( .A(n1066), .B(B[3]), .Y(n516) );
  OAI22XL U538 ( .A0(n1027), .A1(n647), .B0(n6), .B1(n599), .Y(n630) );
  OAI22XL U539 ( .A0(n957), .A1(n624), .B0(n956), .B1(n592), .Y(n625) );
  OAI22XL U540 ( .A0(n997), .A1(n622), .B0(n978), .B1(n582), .Y(n627) );
  OAI22XL U541 ( .A0(n1039), .A1(n623), .B0(n1037), .B1(n583), .Y(n626) );
  OAI22XL U542 ( .A0(n957), .A1(n643), .B0(n956), .B1(n624), .Y(n644) );
  OAI22XL U543 ( .A0(n1039), .A1(n642), .B0(n1037), .B1(n623), .Y(n645) );
  OAI22XL U544 ( .A0(n997), .A1(n641), .B0(n978), .B1(n622), .Y(n646) );
  ADDFX2 U545 ( .A(n676), .B(n675), .CI(n674), .CO(n694), .S(n722) );
  OAI22XL U546 ( .A0(n957), .A1(n673), .B0(n956), .B1(n643), .Y(n674) );
  OAI22XL U547 ( .A0(n1039), .A1(n672), .B0(n1037), .B1(n642), .Y(n675) );
  OAI22XL U548 ( .A0(n997), .A1(n671), .B0(n640), .B1(n641), .Y(n676) );
  ADDFX2 U549 ( .A(n705), .B(n704), .CI(n703), .CO(n723), .S(n752) );
  OAI22XL U550 ( .A0(n957), .A1(n702), .B0(n956), .B1(n673), .Y(n703) );
  OAI22XL U551 ( .A0(n997), .A1(n701), .B0(n978), .B1(n671), .Y(n705) );
  ADDFX2 U552 ( .A(n735), .B(n734), .CI(n733), .CO(n753), .S(n783) );
  OAI22XL U553 ( .A0(n957), .A1(n732), .B0(n956), .B1(n702), .Y(n733) );
  OAI22XL U554 ( .A0(n997), .A1(n730), .B0(n978), .B1(n701), .Y(n735) );
  ADDFX2 U555 ( .A(n765), .B(n764), .CI(n763), .CO(n784), .S(n813) );
  OAI22XL U556 ( .A0(n957), .A1(n762), .B0(n956), .B1(n732), .Y(n763) );
  OAI22XL U557 ( .A0(n1039), .A1(n761), .B0(n1037), .B1(n731), .Y(n764) );
  OAI22XL U558 ( .A0(n997), .A1(n760), .B0(n640), .B1(n730), .Y(n765) );
  OAI22XL U559 ( .A0(n957), .A1(n824), .B0(n956), .B1(n762), .Y(n793) );
  OAI22XL U560 ( .A0(n1039), .A1(n792), .B0(n1037), .B1(n761), .Y(n794) );
  OAI22XL U561 ( .A0(n997), .A1(n791), .B0(n640), .B1(n760), .Y(n795) );
  OAI22XL U562 ( .A0(n957), .A1(n856), .B0(n956), .B1(n825), .Y(n853) );
  OAI22XL U563 ( .A0(n1039), .A1(n852), .B0(n1037), .B1(n822), .Y(n854) );
  XOR2XL U564 ( .A(n995), .B(n65), .Y(n64) );
  XNOR2XL U565 ( .A(n1001), .B(n928), .Y(n856) );
  OAI22XL U566 ( .A0(n1024), .A1(n875), .B0(n851), .B1(n1021), .Y(n879) );
  OAI22XL U567 ( .A0(n1070), .A1(n882), .B0(n5), .B1(n858), .Y(n878) );
  OAI22XL U568 ( .A0(n935), .A1(n910), .B0(n942), .B1(n884), .Y(n922) );
  OAI22XL U569 ( .A0(n1027), .A1(n914), .B0(n6), .B1(n881), .Y(n924) );
  OAI22XL U570 ( .A0(n1070), .A1(n883), .B0(n5), .B1(n882), .Y(n923) );
  OAI22XL U571 ( .A0(n1039), .A1(n918), .B0(n1037), .B1(n917), .Y(n919) );
  OAI22XL U572 ( .A0(n1024), .A1(n944), .B0(n929), .B1(n1021), .Y(n941) );
  NAND2BXL U573 ( .AN(n1020), .B(B[13]), .Y(n930) );
  OAI22XL U574 ( .A0(n997), .A1(n946), .B0(n640), .B1(n936), .Y(n967) );
  OAI22XL U575 ( .A0(n1031), .A1(n948), .B0(n1029), .B1(n932), .Y(n969) );
  XNOR2XL U576 ( .A(n993), .B(n1000), .Y(n948) );
  XNOR2XL U577 ( .A(n1001), .B(n998), .Y(n955) );
  XNOR2XL U578 ( .A(n954), .B(n953), .Y(n1002) );
  XNOR2XL U579 ( .A(n1001), .B(n1000), .Y(n1032) );
  XNOR2XL U580 ( .A(n1004), .B(n1003), .Y(n1025) );
  XOR2XL U581 ( .A(n995), .B(n62), .Y(n61) );
  XNOR2XL U582 ( .A(n993), .B(n947), .Y(n994) );
  XNOR2XL U583 ( .A(n993), .B(n992), .Y(n1028) );
  XNOR2XL U584 ( .A(B[3]), .B(n950), .Y(n999) );
  XNOR2XL U585 ( .A(B[3]), .B(n998), .Y(n1036) );
  XNOR2XL U586 ( .A(n1004), .B(n992), .Y(n973) );
  OAI22XL U587 ( .A0(n1070), .A1(n99), .B0(n5), .B1(n80), .Y(n168) );
  OAI22XL U588 ( .A0(n8), .A1(n100), .B0(n942), .B1(n95), .Y(n171) );
  OAI22XL U589 ( .A0(n1039), .A1(n40), .B0(n1037), .B1(n379), .Y(n380) );
  NAND2BXL U590 ( .AN(n1020), .B(B[3]), .Y(n379) );
  XNOR2XL U591 ( .A(B[3]), .B(n1020), .Y(n378) );
  OAI22XL U592 ( .A0(n1024), .A1(n383), .B0(n382), .B1(n1021), .Y(n396) );
  OAI22XL U593 ( .A0(n952), .A1(n385), .B0(n1037), .B1(n384), .Y(n395) );
  XNOR2XL U594 ( .A(n1164), .B(n1222), .Y(PRODUCT[39]) );
  XNOR2XL U595 ( .A(n1174), .B(n1173), .Y(PRODUCT[38]) );
  NAND2XL U596 ( .A(n1172), .B(n1224), .Y(n1173) );
  NAND2XL U597 ( .A(n1131), .B(n1226), .Y(n1132) );
  OAI22XL U598 ( .A0(n1039), .A1(n888), .B0(n1037), .B1(n852), .Y(n892) );
  OAI22XL U599 ( .A0(n1027), .A1(n881), .B0(n6), .B1(n865), .Y(n893) );
  NOR2XL U600 ( .A(n9), .B(n192), .Y(n207) );
  OAI22XL U601 ( .A0(n8), .A1(n202), .B0(n942), .B1(n191), .Y(n208) );
  XNOR2XL U602 ( .A(n1064), .B(n799), .Y(n192) );
  ADDFX2 U603 ( .A(n480), .B(n479), .CI(n478), .CO(n463), .S(n508) );
  OAI22XL U604 ( .A0(n997), .A1(n485), .B0(n978), .B1(n455), .Y(n475) );
  OAI22XL U605 ( .A0(n1070), .A1(n483), .B0(n5), .B1(n454), .Y(n476) );
  OAI22XL U606 ( .A0(n1070), .A1(n563), .B0(n5), .B1(n542), .Y(n595) );
  OAI22XL U607 ( .A0(n1031), .A1(n562), .B0(n1029), .B1(n539), .Y(n597) );
  OAI22XL U608 ( .A0(n1027), .A1(n599), .B0(n6), .B1(n598), .Y(n612) );
  XNOR2XL U609 ( .A(n603), .B(n602), .Y(n610) );
  OAI22XL U610 ( .A0(n957), .A1(n592), .B0(n1033), .B1(n591), .Y(n609) );
  OAI22XL U611 ( .A0(n8), .A1(n606), .B0(n942), .B1(n594), .Y(n607) );
  OAI22XL U612 ( .A0(n997), .A1(n523), .B0(n978), .B1(n492), .Y(n527) );
  OAI22X1 U613 ( .A0(n1070), .A1(n518), .B0(n5), .B1(n491), .Y(n528) );
  OAI22XL U614 ( .A0(n1031), .A1(n519), .B0(n1029), .B1(n490), .Y(n529) );
  ADDFX2 U615 ( .A(n495), .B(n494), .CI(n493), .CO(n510), .S(n534) );
  OAI2BB1XL U616 ( .A0N(n956), .A1N(n957), .B0(n474), .Y(n493) );
  ADDFX2 U617 ( .A(n464), .B(n463), .CI(n462), .CO(n470), .S(n499) );
  OAI22XL U618 ( .A0(n997), .A1(n455), .B0(n978), .B1(n450), .Y(n464) );
  ADDFX2 U619 ( .A(n467), .B(n466), .CI(n465), .CO(n447), .S(n468) );
  INVX1 U620 ( .A(n470), .Y(n58) );
  OAI22XL U621 ( .A0(n521), .A1(n514), .B0(n6), .B1(n484), .Y(n496) );
  OAI22XL U622 ( .A0(n1070), .A1(n491), .B0(n5), .B1(n483), .Y(n497) );
  OAI22XL U623 ( .A0(n1027), .A1(n520), .B0(n6), .B1(n514), .Y(n538) );
  OAI2BB1XL U624 ( .A0N(n1021), .A1N(n771), .B0(n556), .Y(n584) );
  OAI22XL U625 ( .A0(n997), .A1(n582), .B0(n978), .B1(n561), .Y(n586) );
  OAI22XL U626 ( .A0(n957), .A1(n591), .B0(n1033), .B1(n558), .Y(n568) );
  OAI22XL U627 ( .A0(n1027), .A1(n598), .B0(n6), .B1(n559), .Y(n575) );
  OAI22XL U628 ( .A0(n997), .A1(n561), .B0(n978), .B1(n560), .Y(n574) );
  OAI22XL U629 ( .A0(n1031), .A1(n653), .B0(n743), .B1(n604), .Y(n658) );
  OAI22XL U630 ( .A0(n1027), .A1(n677), .B0(n6), .B1(n647), .Y(n661) );
  OAI22XL U631 ( .A0(n1027), .A1(n706), .B0(n6), .B1(n677), .Y(n691) );
  OAI22XL U632 ( .A0(n1031), .A1(n683), .B0(n743), .B1(n653), .Y(n688) );
  CMPR32X1 U633 ( .A(n723), .B(n722), .C(n721), .CO(n697), .S(n724) );
  OAI22XL U634 ( .A0(n1027), .A1(n736), .B0(n6), .B1(n706), .Y(n720) );
  OAI22XL U635 ( .A0(n1031), .A1(n711), .B0(n743), .B1(n683), .Y(n717) );
  ADDFX2 U636 ( .A(n753), .B(n752), .CI(n751), .CO(n726), .S(n754) );
  OAI22XL U637 ( .A0(n1027), .A1(n766), .B0(n6), .B1(n736), .Y(n750) );
  OAI22XL U638 ( .A0(n1031), .A1(n742), .B0(n1029), .B1(n711), .Y(n747) );
  ADDFX2 U639 ( .A(n784), .B(n783), .CI(n782), .CO(n756), .S(n785) );
  OAI22XL U640 ( .A0(n1027), .A1(n796), .B0(n6), .B1(n766), .Y(n781) );
  OAI22XL U641 ( .A0(n1031), .A1(n773), .B0(n743), .B1(n742), .Y(n778) );
  ADDFX2 U642 ( .A(n814), .B(n813), .CI(n812), .CO(n787), .S(n815) );
  OAI22XL U643 ( .A0(n1027), .A1(n823), .B0(n6), .B1(n796), .Y(n811) );
  OAI22XL U644 ( .A0(n1031), .A1(n802), .B0(n1029), .B1(n773), .Y(n808) );
  OAI22XL U645 ( .A0(n1031), .A1(n862), .B0(n1029), .B1(n827), .Y(n840) );
  OAI22XL U646 ( .A0(n957), .A1(n825), .B0(n1033), .B1(n824), .Y(n833) );
  OAI22XL U647 ( .A0(n935), .A1(n860), .B0(n942), .B1(n826), .Y(n832) );
  OAI22XL U648 ( .A0(n1027), .A1(n864), .B0(n6), .B1(n823), .Y(n834) );
  OAI22XL U649 ( .A0(n949), .A1(n827), .B0(n1029), .B1(n802), .Y(n837) );
  OAI22XL U650 ( .A0(n935), .A1(n826), .B0(n942), .B1(n805), .Y(n835) );
  OAI22XL U651 ( .A0(n1039), .A1(n822), .B0(n1037), .B1(n792), .Y(n1195) );
  OAI22XL U652 ( .A0(n997), .A1(n821), .B0(n640), .B1(n791), .Y(n1197) );
  OAI22XL U653 ( .A0(n1031), .A1(n863), .B0(n1029), .B1(n862), .Y(n1194) );
  OAI22XL U654 ( .A0(n1027), .A1(n865), .B0(n6), .B1(n864), .Y(n1193) );
  OAI22XL U655 ( .A0(n957), .A1(n925), .B0(n956), .B1(n906), .Y(n1136) );
  OAI22XL U656 ( .A0(n1031), .A1(n927), .B0(n1029), .B1(n890), .Y(n903) );
  OAI22XL U657 ( .A0(n1039), .A1(n917), .B0(n1037), .B1(n888), .Y(n905) );
  NOR2XL U658 ( .A(n381), .B(n380), .Y(n1209) );
  NAND2XL U659 ( .A(n381), .B(n380), .Y(n1210) );
  AOI21XL U660 ( .A0(n1215), .A1(n1216), .B0(n376), .Y(n1212) );
  INVXL U661 ( .A(n1214), .Y(n376) );
  NAND2XL U662 ( .A(n390), .B(n389), .Y(n1206) );
  AOI21XL U663 ( .A0(n1207), .A1(n388), .B0(n391), .Y(n1204) );
  INVXL U664 ( .A(n1206), .Y(n391) );
  NOR2XL U665 ( .A(n399), .B(n398), .Y(n1201) );
  NAND2XL U666 ( .A(n399), .B(n398), .Y(n1202) );
  XOR2XL U667 ( .A(n1179), .B(n1178), .Y(n1312) );
  NAND2XL U668 ( .A(n1177), .B(n1176), .Y(n1179) );
  INVXL U669 ( .A(n1175), .Y(n1177) );
  NOR2XL U670 ( .A(n1085), .B(n1084), .Y(mult_x_1_n120) );
  ADDFX2 U671 ( .A(n510), .B(n509), .CI(n508), .CO(n504), .S(mult_x_1_n474) );
  NAND2XL U672 ( .A(n1081), .B(n1080), .Y(mult_x_1_n59) );
  NAND2XL U673 ( .A(n1079), .B(n1078), .Y(n1080) );
  NOR2XL U674 ( .A(n1099), .B(n1098), .Y(mult_x_1_n325) );
  NAND2XL U675 ( .A(n1099), .B(n1098), .Y(mult_x_1_n326) );
  NOR2XL U676 ( .A(n1109), .B(n1108), .Y(mult_x_1_n328) );
  NAND2XL U677 ( .A(n1109), .B(n1108), .Y(mult_x_1_n329) );
  NAND2XL U678 ( .A(n1100), .B(n1101), .Y(mult_x_1_n89) );
  INVXL U679 ( .A(n1101), .Y(n439) );
  OAI21XL U680 ( .A0(n58), .A1(n57), .B0(n56), .Y(mult_x_1_n449) );
  OAI21XL U681 ( .A0(n469), .A1(n470), .B0(n468), .Y(n56) );
  NAND2X1 U682 ( .A(n67), .B(n66), .Y(n1015) );
  NAND2XL U683 ( .A(n1045), .B(n1044), .Y(n66) );
  NOR2XL U684 ( .A(n1083), .B(n1082), .Y(mult_x_1_n319) );
  NOR2BXL U685 ( .AN(n1020), .B(n1021), .Y(n1318) );
  NAND2XL U686 ( .A(n1215), .B(n1214), .Y(n1217) );
  XOR2XL U687 ( .A(n1213), .B(n1212), .Y(n1315) );
  NAND2XL U688 ( .A(n1211), .B(n1210), .Y(n1213) );
  INVXL U689 ( .A(n1209), .Y(n1211) );
  XNOR2XL U690 ( .A(n1208), .B(n1207), .Y(n1314) );
  NAND2XL U691 ( .A(n388), .B(n1206), .Y(n1208) );
  XOR2XL U692 ( .A(n1205), .B(n1204), .Y(n1313) );
  NAND2XL U693 ( .A(n1203), .B(n1202), .Y(n1205) );
  INVXL U694 ( .A(n1201), .Y(n1203) );
  NAND2XL U695 ( .A(n1116), .B(n1115), .Y(n1117) );
  INVXL U696 ( .A(n1114), .Y(n1116) );
  CMPR22X1 U697 ( .A(n679), .B(n678), .CO(n659), .S(n690) );
  CMPR22X1 U698 ( .A(n738), .B(n737), .CO(n718), .S(n749) );
  CMPR22X1 U699 ( .A(n829), .B(n828), .CO(n809), .S(n839) );
  CMPR22X1 U700 ( .A(n1007), .B(n1006), .CO(n1018), .S(n1046) );
  OAI22X1 U701 ( .A0(n771), .A1(n589), .B0(n587), .B1(n1021), .Y(n601) );
  OAI22X1 U702 ( .A0(n1031), .A1(n481), .B0(n1029), .B1(n195), .Y(n460) );
  CMPR22X1 U703 ( .A(n601), .B(n600), .CO(n611), .S(n629) );
  CMPR22X1 U704 ( .A(n371), .B(n370), .CO(n365), .S(n392) );
  CMPR22X1 U705 ( .A(n908), .B(n907), .CO(n1139), .S(n1135) );
  XNOR2X1 U706 ( .A(n292), .B(n291), .Y(PRODUCT[25]) );
  NAND2X1 U707 ( .A(n290), .B(n289), .Y(n291) );
  XNOR2X1 U708 ( .A(n314), .B(n313), .Y(PRODUCT[22]) );
  AOI21XL U709 ( .A0(n1168), .A1(n1161), .B0(n1160), .Y(n1162) );
  AOI21XL U710 ( .A0(n1168), .A1(n1167), .B0(n1166), .Y(n1169) );
  AOI21XL U711 ( .A0(n1168), .A1(n1128), .B0(n1127), .Y(n1129) );
  OAI21XL U712 ( .A0(n997), .A1(n64), .B0(n63), .Y(n855) );
  OAI22X1 U713 ( .A0(n8), .A1(n934), .B0(n12), .B1(n933), .Y(n968) );
  OAI22X1 U714 ( .A0(n1027), .A1(n973), .B0(n6), .B1(n915), .Y(n972) );
  XOR2X1 U715 ( .A(B[13]), .B(B[12]), .Y(n77) );
  OR2X2 U716 ( .A(n946), .B(n640), .Y(n59) );
  XOR3X2 U717 ( .A(n1043), .B(n1044), .C(n1045), .Y(n1155) );
  XNOR2X4 U718 ( .A(B[11]), .B(B[12]), .Y(n942) );
  CLKINVX3 U719 ( .A(n349), .Y(n975) );
  OAI21X1 U720 ( .A0(n334), .A1(n340), .B0(n335), .Y(n321) );
  NOR2X2 U721 ( .A(n139), .B(n138), .Y(n282) );
  XNOR2XL U722 ( .A(B[3]), .B(n1003), .Y(n384) );
  XNOR2XL U723 ( .A(n482), .B(n650), .Y(n79) );
  XNOR2X1 U724 ( .A(B[13]), .B(A[16]), .Y(n522) );
  XNOR2XL U725 ( .A(B[16]), .B(A[3]), .Y(n772) );
  XNOR2XL U726 ( .A(n482), .B(n709), .Y(n99) );
  XNOR2XL U727 ( .A(B[16]), .B(n943), .Y(n540) );
  XNOR2XL U728 ( .A(B[3]), .B(n850), .Y(n822) );
  BUFX3 U729 ( .A(n949), .Y(n1031) );
  BUFX4 U730 ( .A(n521), .Y(n1027) );
  XNOR2XL U731 ( .A(n1217), .B(n1216), .Y(n1316) );
  XNOR2X1 U732 ( .A(B[16]), .B(B[15]), .Y(n488) );
  XNOR2XL U733 ( .A(n1064), .B(n680), .Y(n76) );
  OAI22X1 U734 ( .A0(n8), .A1(n78), .B0(n942), .B1(n87), .Y(n1074) );
  XNOR2X1 U735 ( .A(n1064), .B(n739), .Y(n81) );
  INVXL U736 ( .A(n90), .Y(n166) );
  XNOR2XL U737 ( .A(n482), .B(A[24]), .Y(n1069) );
  CMPR32X1 U738 ( .A(n85), .B(n84), .C(n83), .CO(n1061), .S(n103) );
  XNOR2XL U739 ( .A(n1064), .B(n650), .Y(n86) );
  NAND2XL U740 ( .A(n1085), .B(n1084), .Y(mult_x_1_n121) );
  CMPR32X1 U741 ( .A(n91), .B(n89), .C(n90), .CO(n104), .S(n182) );
  CMPR32X1 U742 ( .A(n94), .B(n93), .C(n92), .CO(n102), .S(n181) );
  XNOR2XL U743 ( .A(B[13]), .B(n650), .Y(n100) );
  NOR2X1 U744 ( .A(n9), .B(n96), .Y(n176) );
  XOR2X1 U745 ( .A(B[8]), .B(B[9]), .Y(n97) );
  XNOR2X1 U746 ( .A(B[8]), .B(B[7]), .Y(n406) );
  OAI22XL U747 ( .A0(n1070), .A1(n172), .B0(n5), .B1(n99), .Y(n179) );
  XNOR2XL U748 ( .A(B[13]), .B(n680), .Y(n191) );
  OAI22XL U749 ( .A0(n8), .A1(n191), .B0(n942), .B1(n100), .Y(n178) );
  CMPR32X1 U750 ( .A(n104), .B(n103), .C(n102), .CO(n1085), .S(n105) );
  NOR2XL U751 ( .A(n106), .B(n105), .Y(mult_x_1_n129) );
  NAND2XL U752 ( .A(n106), .B(n105), .Y(mult_x_1_n130) );
  NOR2X1 U753 ( .A(n128), .B(n127), .Y(n315) );
  ADDFHX2 U754 ( .A(n1278), .B(n1276), .CI(n1274), .CO(n129), .S(n128) );
  NOR2XL U755 ( .A(n278), .B(n282), .Y(n254) );
  NOR2X2 U756 ( .A(n122), .B(n121), .Y(n328) );
  NOR2X2 U757 ( .A(n124), .B(n123), .Y(n323) );
  NOR2X2 U758 ( .A(n328), .B(n323), .Y(n126) );
  NOR2XL U759 ( .A(n1296), .B(n1297), .Y(n107) );
  INVXL U760 ( .A(n107), .Y(n1111) );
  NAND2XL U761 ( .A(n346), .B(n1111), .Y(n1120) );
  NOR2X2 U762 ( .A(n114), .B(n1292), .Y(n1122) );
  NOR2X1 U763 ( .A(n1120), .B(n1122), .Y(n116) );
  NOR2XL U764 ( .A(n1233), .B(n1235), .Y(n109) );
  OAI21XL U765 ( .A0(n1233), .A1(n1236), .B0(n1234), .Y(n108) );
  OR2X2 U766 ( .A(n1298), .B(n1299), .Y(n1149) );
  INVXL U767 ( .A(n1232), .Y(n1147) );
  NAND2XL U768 ( .A(n1298), .B(n1299), .Y(n1148) );
  INVXL U769 ( .A(n1148), .Y(n110) );
  NAND2XL U770 ( .A(n1296), .B(n1297), .Y(n1110) );
  INVXL U771 ( .A(n1110), .Y(n344) );
  NAND2XL U772 ( .A(n1293), .B(n1295), .Y(n345) );
  INVXL U773 ( .A(n345), .Y(n113) );
  NAND2X1 U774 ( .A(n122), .B(n121), .Y(n329) );
  OAI21X1 U775 ( .A0(n323), .A1(n329), .B0(n324), .Y(n125) );
  NAND2X1 U776 ( .A(n137), .B(n136), .Y(n289) );
  NAND2X1 U777 ( .A(n139), .B(n138), .Y(n283) );
  NAND2XL U778 ( .A(n143), .B(n142), .Y(n265) );
  OAI21XL U779 ( .A0(n264), .A1(n274), .B0(n265), .Y(n144) );
  AOI21XL U780 ( .A0(n145), .A1(n259), .B0(n144), .Y(n146) );
  NOR2X1 U781 ( .A(n150), .B(n149), .Y(n250) );
  CMPR32X1 U782 ( .A(n1254), .B(n1251), .C(n1252), .CO(n152), .S(n149) );
  CMPR32X1 U783 ( .A(n1246), .B(n1247), .C(n1245), .CO(n155), .S(n154) );
  OR2X2 U784 ( .A(n1241), .B(n1240), .Y(n219) );
  OR2X2 U785 ( .A(n159), .B(n224), .Y(n162) );
  NAND2X1 U786 ( .A(n150), .B(n149), .Y(n251) );
  NAND2XL U787 ( .A(n152), .B(n151), .Y(n246) );
  NAND2XL U788 ( .A(n154), .B(n153), .Y(n241) );
  NAND2XL U789 ( .A(n155), .B(n1244), .Y(n234) );
  OAI21XL U790 ( .A0(n159), .A1(n225), .B0(n158), .Y(n160) );
  CMPR32X1 U791 ( .A(n168), .B(n167), .C(n166), .CO(n92), .S(n211) );
  CMPR32X1 U792 ( .A(n171), .B(n170), .C(n169), .CO(n180), .S(n210) );
  INVXL U793 ( .A(n175), .Y(n203) );
  CMPR32X1 U794 ( .A(n176), .B(n175), .C(n174), .CO(n170), .S(n198) );
  CMPR32X1 U795 ( .A(n179), .B(n178), .C(n177), .CO(n169), .S(n197) );
  CMPR32X1 U796 ( .A(n182), .B(n181), .C(n180), .CO(n106), .S(n183) );
  NOR2XL U797 ( .A(n184), .B(n183), .Y(mult_x_1_n136) );
  NAND2XL U798 ( .A(n184), .B(n183), .Y(mult_x_1_n137) );
  NOR2XL U799 ( .A(n223), .B(n224), .Y(n214) );
  NAND2XL U800 ( .A(n214), .B(n219), .Y(n187) );
  AOI21XL U801 ( .A0(n215), .A1(n219), .B0(n185), .Y(n186) );
  XNOR2X1 U802 ( .A(B[13]), .B(n709), .Y(n202) );
  XOR2X1 U803 ( .A(B[6]), .B(B[7]), .Y(n194) );
  XNOR2XL U804 ( .A(B[7]), .B(A[24]), .Y(n481) );
  INVX8 U805 ( .A(n351), .Y(n993) );
  INVXL U806 ( .A(n195), .Y(n196) );
  CMPR32X1 U807 ( .A(n199), .B(n198), .C(n197), .CO(n209), .S(n448) );
  OAI22XL U808 ( .A0(n1070), .A1(n454), .B0(n5), .B1(n201), .Y(n457) );
  XNOR2X1 U809 ( .A(B[13]), .B(n739), .Y(n451) );
  CMPR32X1 U810 ( .A(n205), .B(n204), .C(n203), .CO(n199), .S(n466) );
  CMPR32X1 U811 ( .A(n208), .B(n207), .C(n206), .CO(n449), .S(n465) );
  CMPR32X1 U812 ( .A(n211), .B(n210), .C(n209), .CO(n184), .S(n212) );
  NOR2XL U813 ( .A(n213), .B(n212), .Y(mult_x_1_n151) );
  NAND2XL U814 ( .A(n213), .B(n212), .Y(mult_x_1_n152) );
  INVXL U815 ( .A(n214), .Y(n217) );
  INVXL U816 ( .A(n215), .Y(n216) );
  OAI21X1 U817 ( .A0(n1171), .A1(n217), .B0(n216), .Y(n221) );
  XNOR2X1 U818 ( .A(n221), .B(n220), .Y(PRODUCT[34]) );
  INVXL U819 ( .A(n230), .Y(n242) );
  NAND2XL U820 ( .A(n229), .B(n242), .Y(n232) );
  AOI21XL U821 ( .A0(n238), .A1(n242), .B0(n11), .Y(n231) );
  INVXL U822 ( .A(n229), .Y(n240) );
  INVXL U823 ( .A(n238), .Y(n239) );
  NAND2X1 U824 ( .A(n242), .B(n241), .Y(n243) );
  XNOR2X2 U825 ( .A(n244), .B(n243), .Y(PRODUCT[31]) );
  OAI21X2 U826 ( .A0(n1171), .A1(n250), .B0(n251), .Y(n249) );
  INVXL U827 ( .A(n245), .Y(n247) );
  INVXL U828 ( .A(n250), .Y(n252) );
  INVXL U829 ( .A(n254), .Y(n269) );
  INVXL U830 ( .A(n255), .Y(n275) );
  NOR2XL U831 ( .A(n269), .B(n255), .Y(n261) );
  NAND2XL U832 ( .A(n261), .B(n287), .Y(n263) );
  INVX4 U833 ( .A(n257), .Y(n319) );
  INVXL U834 ( .A(n259), .Y(n270) );
  OAI21XL U835 ( .A0(n270), .A1(n255), .B0(n274), .Y(n260) );
  OAI21XL U836 ( .A0(n263), .A1(n319), .B0(n262), .Y(n268) );
  NAND2X1 U837 ( .A(n266), .B(n265), .Y(n267) );
  INVXL U838 ( .A(n269), .Y(n271) );
  NAND2XL U839 ( .A(n287), .B(n271), .Y(n273) );
  AOI21XL U840 ( .A0(n288), .A1(n271), .B0(n259), .Y(n272) );
  XNOR2X1 U841 ( .A(n277), .B(n276), .Y(PRODUCT[27]) );
  NAND2XL U842 ( .A(n287), .B(n290), .Y(n281) );
  INVXL U843 ( .A(n289), .Y(n279) );
  XNOR2X1 U844 ( .A(n286), .B(n285), .Y(PRODUCT[26]) );
  OAI21X1 U845 ( .A0(n319), .A1(n256), .B0(n258), .Y(n292) );
  NAND2XL U846 ( .A(n293), .B(n307), .Y(n297) );
  INVXL U847 ( .A(n306), .Y(n295) );
  AOI21XL U848 ( .A0(n303), .A1(n307), .B0(n295), .Y(n296) );
  OAI21XL U849 ( .A0(n319), .A1(n297), .B0(n296), .Y(n302) );
  NAND2X1 U850 ( .A(n300), .B(n299), .Y(n301) );
  INVXL U851 ( .A(n293), .Y(n305) );
  INVXL U852 ( .A(n303), .Y(n304) );
  OAI21XL U853 ( .A0(n319), .A1(n305), .B0(n304), .Y(n309) );
  NAND2X1 U854 ( .A(n307), .B(n306), .Y(n308) );
  XNOR2X1 U855 ( .A(n309), .B(n308), .Y(PRODUCT[23]) );
  OAI21XL U856 ( .A0(n319), .A1(n315), .B0(n316), .Y(n314) );
  INVXL U857 ( .A(n310), .Y(n312) );
  INVXL U858 ( .A(n315), .Y(n317) );
  INVX1 U859 ( .A(n320), .Y(n342) );
  INVXL U860 ( .A(n328), .Y(n330) );
  NAND2XL U861 ( .A(n330), .B(n329), .Y(n331) );
  NAND2XL U862 ( .A(n10), .B(n340), .Y(n341) );
  XNOR2X1 U863 ( .A(n342), .B(n341), .Y(PRODUCT[17]) );
  OAI21XL U864 ( .A0(n1121), .A1(n107), .B0(n1110), .Y(n348) );
  XNOR2X1 U865 ( .A(n348), .B(n347), .Y(PRODUCT[15]) );
  INVX1 U866 ( .A(B[0]), .Y(n769) );
  NAND2X1 U867 ( .A(B[1]), .B(n769), .Y(n771) );
  XNOR2XL U868 ( .A(n975), .B(n1000), .Y(n352) );
  BUFX3 U869 ( .A(n769), .Y(n1021) );
  OAI22X1 U870 ( .A0(n1024), .A1(n352), .B0(n417), .B1(n1021), .Y(n412) );
  OAI22X1 U871 ( .A0(n1031), .A1(n351), .B0(n1029), .B1(n350), .Y(n411) );
  XNOR2XL U872 ( .A(n975), .B(n947), .Y(n359) );
  OAI22XL U873 ( .A0(n1024), .A1(n359), .B0(n352), .B1(n1021), .Y(n362) );
  XNOR2XL U874 ( .A(n1001), .B(n1003), .Y(n357) );
  OAI22XL U875 ( .A0(n957), .A1(n368), .B0(n1033), .B1(n357), .Y(n361) );
  BUFX3 U876 ( .A(n355), .Y(n1037) );
  XNOR2XL U877 ( .A(n993), .B(n1020), .Y(n356) );
  OAI22X1 U878 ( .A0(n1024), .A1(n382), .B0(n359), .B1(n1021), .Y(n371) );
  OAI22X1 U879 ( .A0(n957), .A1(n472), .B0(n1033), .B1(n360), .Y(n370) );
  CMPR32X1 U880 ( .A(n363), .B(n362), .C(n361), .CO(n433), .S(n364) );
  CMPR32X1 U881 ( .A(n366), .B(n365), .C(n364), .CO(n402), .S(n401) );
  NOR2XL U882 ( .A(n1114), .B(n1175), .Y(n405) );
  OAI22X1 U883 ( .A0(n1024), .A1(n377), .B0(n383), .B1(n1021), .Y(n387) );
  OAI22X1 U884 ( .A0(n952), .A1(n378), .B0(n1037), .B1(n385), .Y(n386) );
  OAI21XL U885 ( .A0(n1212), .A1(n1209), .B0(n1210), .Y(n1207) );
  CMPR22X1 U886 ( .A(n387), .B(n386), .CO(n389), .S(n381) );
  CMPR32X1 U887 ( .A(n394), .B(n393), .C(n392), .CO(n400), .S(n399) );
  CMPR32X1 U888 ( .A(n397), .B(n396), .C(n395), .CO(n398), .S(n390) );
  OAI21XL U889 ( .A0(n1204), .A1(n1201), .B0(n1202), .Y(n1113) );
  NAND2XL U890 ( .A(n403), .B(n402), .Y(n1115) );
  OAI21XL U891 ( .A0(n1114), .A1(n1176), .B0(n1115), .Y(n404) );
  AOI21XL U892 ( .A0(n405), .A1(n1113), .B0(n404), .Y(n442) );
  XNOR2X1 U893 ( .A(n993), .B(A[3]), .Y(n1030) );
  CMPR22X1 U894 ( .A(n412), .B(n411), .CO(n426), .S(n434) );
  OAI22X1 U895 ( .A0(n1024), .A1(n416), .B0(n1023), .B1(n1021), .Y(n1050) );
  OAI22X1 U896 ( .A0(n1027), .A1(n415), .B0(n6), .B1(n414), .Y(n1049) );
  OAI22XL U897 ( .A0(n1031), .A1(n419), .B0(n1029), .B1(n418), .Y(n420) );
  CMPR32X1 U898 ( .A(n422), .B(n421), .C(n420), .CO(n1092), .S(n431) );
  CMPR32X1 U899 ( .A(n425), .B(n424), .C(n423), .CO(n430), .S(n432) );
  CMPR32X1 U900 ( .A(n428), .B(n427), .C(n426), .CO(n1106), .S(n429) );
  CMPR32X1 U901 ( .A(n434), .B(n433), .C(n432), .CO(n435), .S(n403) );
  NAND2XL U902 ( .A(n1100), .B(n445), .Y(n441) );
  OAI21XL U903 ( .A0(n442), .A1(n441), .B0(n440), .Y(mult_x_1_n331) );
  INVXL U904 ( .A(n442), .Y(n446) );
  AOI21XL U905 ( .A0(n446), .A1(n445), .B0(n444), .Y(mult_x_1_n338) );
  CMPR32X1 U906 ( .A(n449), .B(n448), .C(n447), .CO(n213), .S(mult_x_1_n442)
         );
  XNOR2X1 U907 ( .A(B[13]), .B(A[18]), .Y(n486) );
  INVXL U908 ( .A(n460), .Y(n478) );
  XNOR2X1 U909 ( .A(n1064), .B(n850), .Y(n453) );
  CMPR32X1 U910 ( .A(n458), .B(n457), .C(n456), .CO(n467), .S(n501) );
  CMPR32X1 U911 ( .A(n461), .B(n460), .C(n459), .CO(n206), .S(n500) );
  XNOR2XL U912 ( .A(n1064), .B(n874), .Y(n471) );
  NOR2XL U913 ( .A(n9), .B(n471), .Y(n495) );
  XNOR2XL U914 ( .A(n954), .B(A[24]), .Y(n517) );
  INVXL U915 ( .A(n473), .Y(n474) );
  CMPR32X1 U916 ( .A(n477), .B(n476), .C(n475), .CO(n462), .S(n509) );
  XNOR2X1 U917 ( .A(n993), .B(n1063), .Y(n490) );
  OAI22XL U918 ( .A0(n1031), .A1(n490), .B0(n1029), .B1(n481), .Y(n498) );
  OAI22X1 U919 ( .A0(n997), .A1(n492), .B0(n978), .B1(n485), .Y(n513) );
  XNOR2X1 U920 ( .A(B[13]), .B(n799), .Y(n487) );
  OAI22X2 U921 ( .A0(n8), .A1(n487), .B0(n942), .B1(n486), .Y(n512) );
  XNOR2X1 U922 ( .A(n1064), .B(A[13]), .Y(n489) );
  INVXL U923 ( .A(n494), .Y(n524) );
  XNOR2X1 U924 ( .A(B[7]), .B(n650), .Y(n519) );
  CLKINVX3 U925 ( .A(n877), .Y(n1067) );
  CMPR32X1 U926 ( .A(n498), .B(n497), .C(n496), .CO(n507), .S(n533) );
  CMPR32X1 U927 ( .A(n504), .B(n503), .C(n502), .CO(mult_x_1_n459), .S(
        mult_x_1_n460) );
  NOR2X1 U928 ( .A(n9), .B(n515), .Y(n572) );
  OAI22XL U929 ( .A0(n957), .A1(n558), .B0(n1033), .B1(n517), .Y(n545) );
  XNOR2XL U930 ( .A(n1067), .B(A[13]), .Y(n542) );
  OAI22X1 U931 ( .A0(n1070), .A1(n542), .B0(n5), .B1(n518), .Y(n544) );
  XNOR2X1 U932 ( .A(n993), .B(n680), .Y(n539) );
  XNOR2XL U933 ( .A(B[13]), .B(n850), .Y(n557) );
  OAI22XL U934 ( .A0(n8), .A1(n557), .B0(n942), .B1(n522), .Y(n547) );
  ADDFHX1 U935 ( .A(n529), .B(n528), .CI(n527), .CO(n535), .S(n549) );
  CMPR32X1 U936 ( .A(n532), .B(n531), .C(n530), .CO(mult_x_1_n483), .S(
        mult_x_1_n484) );
  ADDFHX1 U937 ( .A(n535), .B(n534), .CI(n533), .CO(n505), .S(mult_x_1_n486)
         );
  CMPR32X1 U938 ( .A(n538), .B(n537), .C(n536), .CO(n531), .S(n554) );
  XNOR2X1 U939 ( .A(B[7]), .B(n709), .Y(n562) );
  XNOR2XL U940 ( .A(n1067), .B(n928), .Y(n563) );
  CMPR32X1 U941 ( .A(n545), .B(n544), .C(n543), .CO(n536), .S(n565) );
  CMPR32X1 U942 ( .A(n548), .B(n547), .C(n546), .CO(n551), .S(n564) );
  CMPR32X1 U943 ( .A(n551), .B(n550), .C(n549), .CO(n530), .S(n552) );
  OAI22XL U944 ( .A0(n1039), .A1(n583), .B0(n1037), .B1(n555), .Y(n585) );
  INVXL U945 ( .A(n587), .Y(n556) );
  XNOR2XL U946 ( .A(B[13]), .B(n874), .Y(n594) );
  OAI22XL U947 ( .A0(n8), .A1(n594), .B0(n942), .B1(n557), .Y(n569) );
  INVXL U948 ( .A(n571), .Y(n567) );
  XNOR2XL U949 ( .A(n1067), .B(n943), .Y(n605) );
  OR2X2 U950 ( .A(n603), .B(n602), .Y(n573) );
  CMPR32X1 U951 ( .A(n569), .B(n568), .C(n567), .CO(n581), .S(n620) );
  CMPR32X1 U952 ( .A(n572), .B(n571), .C(n570), .CO(n537), .S(n580) );
  CMPR32X1 U953 ( .A(n575), .B(n574), .C(n573), .CO(n579), .S(n619) );
  CMPR32X1 U954 ( .A(n578), .B(n577), .C(n576), .CO(mult_x_1_n509), .S(
        mult_x_1_n510) );
  CMPR32X1 U955 ( .A(n581), .B(n580), .C(n579), .CO(mult_x_1_n513), .S(n576)
         );
  XNOR2XL U956 ( .A(n954), .B(n680), .Y(n592) );
  CMPR32X1 U957 ( .A(n586), .B(n585), .C(n584), .CO(n621), .S(n632) );
  NOR2X1 U958 ( .A(n9), .B(n588), .Y(n600) );
  OAI22XL U959 ( .A0(n771), .A1(n651), .B0(n589), .B1(n1021), .Y(n649) );
  XNOR2X1 U960 ( .A(B[16]), .B(n998), .Y(n590) );
  NOR2X1 U961 ( .A(n9), .B(n590), .Y(n648) );
  XNOR2XL U962 ( .A(B[13]), .B(A[13]), .Y(n606) );
  CMPR32X1 U963 ( .A(n597), .B(n596), .C(n595), .CO(n566), .S(n617) );
  XNOR2X1 U964 ( .A(n993), .B(A[18]), .Y(n653) );
  OAI22X1 U965 ( .A0(n1070), .A1(n654), .B0(n5), .B1(n605), .Y(n657) );
  XNOR2XL U966 ( .A(B[13]), .B(n928), .Y(n655) );
  OAI22XL U967 ( .A0(n935), .A1(n655), .B0(n942), .B1(n606), .Y(n656) );
  CMPR32X1 U968 ( .A(n609), .B(n608), .C(n607), .CO(n618), .S(n635) );
  CMPR32X1 U969 ( .A(n612), .B(n611), .C(n610), .CO(n616), .S(n634) );
  CMPR32X1 U970 ( .A(n615), .B(n614), .C(n613), .CO(mult_x_1_n523), .S(
        mult_x_1_n524) );
  CMPR32X1 U971 ( .A(n618), .B(n617), .C(n616), .CO(mult_x_1_n525), .S(n614)
         );
  CMPR32X1 U972 ( .A(n621), .B(n620), .C(n619), .CO(n578), .S(mult_x_1_n528)
         );
  CMPR32X1 U973 ( .A(n627), .B(n626), .C(n625), .CO(n633), .S(n663) );
  CMPR32X1 U974 ( .A(n630), .B(n629), .C(n628), .CO(n631), .S(n662) );
  CMPR32X1 U975 ( .A(n633), .B(n632), .C(n631), .CO(n615), .S(n638) );
  CMPR32X1 U976 ( .A(n636), .B(n635), .C(n634), .CO(n613), .S(n637) );
  CMPR32X1 U977 ( .A(n646), .B(n645), .C(n644), .CO(n664), .S(n693) );
  ADDHXL U978 ( .A(n649), .B(n648), .CO(n628), .S(n660) );
  OAI22X1 U979 ( .A0(n771), .A1(n681), .B0(n651), .B1(n1021), .Y(n679) );
  XNOR2X1 U980 ( .A(B[16]), .B(n953), .Y(n652) );
  NOR2X1 U981 ( .A(n9), .B(n652), .Y(n678) );
  XNOR2X1 U982 ( .A(B[7]), .B(n799), .Y(n683) );
  XNOR2X1 U983 ( .A(n1067), .B(n950), .Y(n684) );
  OAI22X1 U984 ( .A0(n713), .A1(n684), .B0(n5), .B1(n654), .Y(n687) );
  XNOR2XL U985 ( .A(B[13]), .B(n943), .Y(n685) );
  OAI22XL U986 ( .A0(n935), .A1(n685), .B0(n942), .B1(n655), .Y(n686) );
  CMPR32X1 U987 ( .A(n658), .B(n657), .C(n656), .CO(n636), .S(n669) );
  CMPR32X1 U988 ( .A(n661), .B(n659), .C(n660), .CO(n668), .S(n692) );
  CMPR32X1 U989 ( .A(n664), .B(n663), .C(n662), .CO(n639), .S(n665) );
  CMPR32X1 U990 ( .A(n667), .B(n666), .C(n665), .CO(mult_x_1_n555), .S(
        mult_x_1_n556) );
  CMPR32X1 U991 ( .A(n670), .B(n669), .C(n668), .CO(mult_x_1_n557), .S(n666)
         );
  NOR2X1 U992 ( .A(n9), .B(n682), .Y(n707) );
  XNOR2X1 U993 ( .A(n993), .B(A[16]), .Y(n711) );
  XNOR2X1 U994 ( .A(n1067), .B(n998), .Y(n712) );
  OAI22X1 U995 ( .A0(n713), .A1(n712), .B0(n5), .B1(n684), .Y(n716) );
  OAI22XL U996 ( .A0(n935), .A1(n714), .B0(n942), .B1(n685), .Y(n715) );
  CMPR32X1 U997 ( .A(n688), .B(n687), .C(n686), .CO(n670), .S(n699) );
  CMPR32X1 U998 ( .A(n691), .B(n690), .C(n689), .CO(n698), .S(n721) );
  CMPR32X1 U999 ( .A(n694), .B(n693), .C(n692), .CO(n667), .S(n695) );
  CMPR32X1 U1000 ( .A(n697), .B(n696), .C(n695), .CO(mult_x_1_n571), .S(
        mult_x_1_n572) );
  CMPR32X1 U1001 ( .A(n700), .B(n699), .C(n698), .CO(mult_x_1_n573), .S(n696)
         );
  ADDHXL U1002 ( .A(n708), .B(n707), .CO(n689), .S(n719) );
  XNOR2X1 U1003 ( .A(B[16]), .B(n947), .Y(n710) );
  NOR2X1 U1004 ( .A(n9), .B(n710), .Y(n737) );
  CMPR32X1 U1005 ( .A(n717), .B(n716), .C(n715), .CO(n700), .S(n728) );
  CMPR32X1 U1006 ( .A(n720), .B(n718), .C(n719), .CO(n727), .S(n751) );
  CMPR32X1 U1007 ( .A(n726), .B(n725), .C(n724), .CO(mult_x_1_n587), .S(
        mult_x_1_n588) );
  CMPR32X1 U1008 ( .A(n729), .B(n728), .C(n727), .CO(mult_x_1_n589), .S(n725)
         );
  XNOR2X1 U1009 ( .A(B[16]), .B(n992), .Y(n741) );
  NOR2X1 U1010 ( .A(n9), .B(n741), .Y(n767) );
  XNOR2X1 U1011 ( .A(n993), .B(n874), .Y(n773) );
  OAI22X1 U1012 ( .A0(n1070), .A1(n774), .B0(n5), .B1(n744), .Y(n777) );
  XNOR2XL U1013 ( .A(B[13]), .B(n998), .Y(n775) );
  OAI22XL U1014 ( .A0(n8), .A1(n775), .B0(n12), .B1(n745), .Y(n776) );
  CMPR32X1 U1015 ( .A(n750), .B(n749), .C(n748), .CO(n757), .S(n782) );
  CMPR32X1 U1016 ( .A(n759), .B(n758), .C(n757), .CO(mult_x_1_n605), .S(n755)
         );
  ADDHXL U1017 ( .A(n768), .B(n767), .CO(n748), .S(n780) );
  OAI22X1 U1018 ( .A0(n771), .A1(n800), .B0(n770), .B1(n769), .Y(n798) );
  XNOR2X1 U1019 ( .A(n993), .B(A[13]), .Y(n802) );
  XNOR2X1 U1020 ( .A(n1067), .B(n947), .Y(n803) );
  OAI22X1 U1021 ( .A0(n1070), .A1(n803), .B0(n5), .B1(n774), .Y(n807) );
  XNOR2X1 U1022 ( .A(B[13]), .B(n953), .Y(n805) );
  OAI22XL U1023 ( .A0(n935), .A1(n805), .B0(n942), .B1(n775), .Y(n806) );
  CMPR32X1 U1024 ( .A(n778), .B(n777), .C(n776), .CO(n759), .S(n789) );
  CMPR32X1 U1025 ( .A(n781), .B(n779), .C(n780), .CO(n788), .S(n812) );
  CMPR32X1 U1026 ( .A(n787), .B(n786), .C(n785), .CO(mult_x_1_n619), .S(
        mult_x_1_n620) );
  CMPR32X1 U1027 ( .A(n790), .B(n789), .C(n788), .CO(mult_x_1_n621), .S(n786)
         );
  XNOR2XL U1028 ( .A(n1067), .B(A[3]), .Y(n857) );
  OAI22XL U1029 ( .A0(n1070), .A1(n857), .B0(n5), .B1(n804), .Y(n1196) );
  CMPR32X1 U1030 ( .A(n795), .B(n794), .C(n793), .CO(n814), .S(n842) );
  CMPR22X1 U1031 ( .A(n798), .B(n797), .CO(n779), .S(n810) );
  OAI22X1 U1032 ( .A0(n1024), .A1(n830), .B0(n800), .B1(n1021), .Y(n829) );
  XNOR2XL U1033 ( .A(B[16]), .B(n1003), .Y(n801) );
  XNOR2X1 U1034 ( .A(n993), .B(n928), .Y(n827) );
  OAI22XL U1035 ( .A0(n1070), .A1(n804), .B0(n5), .B1(n803), .Y(n836) );
  XNOR2X1 U1036 ( .A(B[13]), .B(n1000), .Y(n826) );
  CMPR32X1 U1037 ( .A(n808), .B(n807), .C(n806), .CO(n790), .S(n819) );
  CMPR32X1 U1038 ( .A(n811), .B(n810), .C(n809), .CO(n818), .S(n841) );
  CMPR32X1 U1039 ( .A(n817), .B(n816), .C(n815), .CO(mult_x_1_n635), .S(
        mult_x_1_n636) );
  CMPR32X1 U1040 ( .A(n820), .B(n819), .C(n818), .CO(mult_x_1_n637), .S(n816)
         );
  XNOR2XL U1041 ( .A(B[13]), .B(n947), .Y(n860) );
  XNOR2X1 U1042 ( .A(n993), .B(n943), .Y(n862) );
  CMPR32X1 U1043 ( .A(n834), .B(n833), .C(n832), .CO(n849), .S(n869) );
  CMPR32X1 U1044 ( .A(n837), .B(n836), .C(n835), .CO(n820), .S(n848) );
  CMPR32X1 U1045 ( .A(n840), .B(n839), .C(n838), .CO(n847), .S(n868) );
  CMPR32X1 U1046 ( .A(n843), .B(n842), .C(n841), .CO(n817), .S(n844) );
  CMPR32X1 U1047 ( .A(n846), .B(n845), .C(n844), .CO(mult_x_1_n651), .S(
        mult_x_1_n652) );
  XNOR2XL U1048 ( .A(n1067), .B(n1003), .Y(n858) );
  XNOR2X1 U1049 ( .A(B[13]), .B(A[3]), .Y(n884) );
  XNOR2XL U1050 ( .A(B[13]), .B(n992), .Y(n861) );
  OAI22XL U1051 ( .A0(n8), .A1(n884), .B0(n12), .B1(n861), .Y(n891) );
  CMPR32X1 U1052 ( .A(n855), .B(n854), .C(n853), .CO(n870), .S(n885) );
  OAI22X1 U1053 ( .A0(n1035), .A1(n906), .B0(n1033), .B1(n856), .Y(n896) );
  XNOR2X1 U1054 ( .A(n993), .B(n950), .Y(n890) );
  XNOR2X1 U1055 ( .A(n993), .B(n974), .Y(n863) );
  OAI22XL U1056 ( .A0(n1070), .A1(n858), .B0(n5), .B1(n857), .Y(n1191) );
  XNOR2X1 U1057 ( .A(B[16]), .B(n945), .Y(n859) );
  OAI22XL U1058 ( .A0(n935), .A1(n861), .B0(n942), .B1(n860), .Y(n1189) );
  ADDHXL U1059 ( .A(n867), .B(n866), .CO(n838), .S(n1192) );
  CMPR32X1 U1060 ( .A(n873), .B(n872), .C(n871), .CO(mult_x_1_n667), .S(
        mult_x_1_n668) );
  OAI22X1 U1061 ( .A0(n1024), .A1(n909), .B0(n875), .B1(n1021), .Y(n908) );
  OAI22X1 U1062 ( .A0(n1070), .A1(n877), .B0(n5), .B1(n876), .Y(n907) );
  CMPR32X1 U1063 ( .A(n880), .B(n879), .C(n878), .CO(n887), .S(n1138) );
  XNOR2XL U1064 ( .A(B[13]), .B(n1003), .Y(n910) );
  CMPR32X1 U1065 ( .A(n887), .B(n886), .C(n885), .CO(n873), .S(n898) );
  XNOR2XL U1066 ( .A(n995), .B(n992), .Y(n916) );
  OAI22XL U1067 ( .A0(n997), .A1(n916), .B0(n640), .B1(n889), .Y(n904) );
  XNOR2X1 U1068 ( .A(n993), .B(n998), .Y(n927) );
  CMPR32X1 U1069 ( .A(n893), .B(n892), .C(n891), .CO(n886), .S(n1153) );
  CMPR32X1 U1070 ( .A(n896), .B(n895), .C(n894), .CO(n902), .S(n1152) );
  CMPR32X1 U1071 ( .A(n899), .B(n898), .C(n897), .CO(mult_x_1_n683), .S(
        mult_x_1_n684) );
  CMPR32X1 U1072 ( .A(n902), .B(n901), .C(n900), .CO(n872), .S(mult_x_1_n686)
         );
  CMPR32X1 U1073 ( .A(n905), .B(n904), .C(n903), .CO(n1154), .S(n960) );
  XNOR2X1 U1074 ( .A(B[13]), .B(n945), .Y(n933) );
  OAI22XL U1075 ( .A0(n935), .A1(n933), .B0(n942), .B1(n910), .Y(n911) );
  CMPR32X1 U1076 ( .A(n913), .B(n912), .C(n911), .CO(n1134), .S(n966) );
  XNOR2XL U1077 ( .A(n1004), .B(n947), .Y(n915) );
  XNOR2X1 U1078 ( .A(B[3]), .B(n974), .Y(n951) );
  OAI22X1 U1079 ( .A0(n1039), .A1(n951), .B0(n1037), .B1(n918), .Y(n971) );
  OAI22X1 U1080 ( .A0(n957), .A1(n955), .B0(n956), .B1(n926), .Y(n970) );
  OAI22XL U1081 ( .A0(n1027), .A1(n915), .B0(n6), .B1(n914), .Y(n921) );
  XNOR2XL U1082 ( .A(n995), .B(A[3]), .Y(n936) );
  OAI22XL U1083 ( .A0(n997), .A1(n936), .B0(n640), .B1(n916), .Y(n920) );
  CMPR32X1 U1084 ( .A(n921), .B(n920), .C(n919), .CO(n1142), .S(n964) );
  CMPR32X1 U1085 ( .A(n924), .B(n923), .C(n922), .CO(n1137), .S(n1141) );
  XNOR2X1 U1086 ( .A(B[7]), .B(n953), .Y(n932) );
  XNOR2XL U1087 ( .A(n975), .B(n928), .Y(n944) );
  OAI22XL U1088 ( .A0(n8), .A1(n931), .B0(n942), .B1(n930), .Y(n940) );
  XNOR2XL U1089 ( .A(B[13]), .B(n1020), .Y(n934) );
  CMPR32X1 U1090 ( .A(n939), .B(n938), .C(n937), .CO(n1140), .S(n984) );
  ADDHXL U1091 ( .A(n941), .B(n940), .CO(n937), .S(n991) );
  OAI22XL U1092 ( .A0(n1024), .A1(n976), .B0(n944), .B1(n1021), .Y(n981) );
  OAI22X1 U1093 ( .A0(n949), .A1(n994), .B0(n1029), .B1(n948), .Y(n1010) );
  CMPR32X1 U1094 ( .A(n963), .B(n962), .C(n961), .CO(mult_x_1_n711), .S(
        mult_x_1_n712) );
  CMPR32X1 U1095 ( .A(n966), .B(n965), .C(n964), .CO(n958), .S(n988) );
  CMPR32X1 U1096 ( .A(n969), .B(n968), .C(n967), .CO(n985), .S(n1013) );
  CMPR32X1 U1097 ( .A(n972), .B(n971), .C(n970), .CO(n965), .S(n1012) );
  XNOR2XL U1098 ( .A(n1004), .B(A[3]), .Y(n1005) );
  OAI22X1 U1099 ( .A0(n1024), .A1(n1022), .B0(n976), .B1(n1021), .Y(n1007) );
  OAI22X1 U1100 ( .A0(n997), .A1(n979), .B0(n978), .B1(n977), .Y(n1006) );
  CMPR32X1 U1101 ( .A(n982), .B(n981), .C(n980), .CO(n990), .S(n1017) );
  CMPR32X1 U1102 ( .A(n989), .B(n990), .C(n991), .CO(n983), .S(n1016) );
  XNOR2XL U1103 ( .A(n995), .B(n1020), .Y(n996) );
  OAI22XL U1104 ( .A0(n1027), .A1(n1025), .B0(n6), .B1(n1005), .Y(n1047) );
  CMPR32X1 U1105 ( .A(n1010), .B(n1009), .C(n1008), .CO(n989), .S(n1043) );
  CMPR32X1 U1106 ( .A(n1013), .B(n1012), .C(n1011), .CO(n987), .S(n1014) );
  CMPR32X1 U1107 ( .A(n1016), .B(n1015), .C(n1014), .CO(mult_x_1_n737), .S(
        mult_x_1_n738) );
  CMPR32X1 U1108 ( .A(n1019), .B(n1018), .C(n1017), .CO(n1011), .S(n1157) );
  CMPR32X1 U1109 ( .A(n1042), .B(n1041), .C(n1040), .CO(n1045), .S(n1057) );
  CMPR32X1 U1110 ( .A(n1048), .B(n1047), .C(n1046), .CO(n1044), .S(n1088) );
  CMPR22X1 U1111 ( .A(n1050), .B(n1049), .CO(n1097), .S(n1093) );
  CMPR32X1 U1112 ( .A(n1053), .B(n1052), .C(n1051), .CO(n1059), .S(n1096) );
  CMPR32X1 U1113 ( .A(n1056), .B(n1055), .C(n1054), .CO(n1095), .S(n1107) );
  CMPR32X1 U1114 ( .A(n1059), .B(n1058), .C(n1057), .CO(n1156), .S(n1086) );
  CMPR32X1 U1115 ( .A(n1062), .B(n1061), .C(n1060), .CO(n1079), .S(n1084) );
  XNOR2XL U1116 ( .A(n1064), .B(n1063), .Y(n1065) );
  CMPR32X1 U1117 ( .A(n1074), .B(n1073), .C(n1072), .CO(n1075), .S(n1060) );
  CMPR32X1 U1118 ( .A(n1077), .B(n1076), .C(n1075), .S(n1078) );
  CMPR32X1 U1119 ( .A(n1088), .B(n1087), .C(n1086), .CO(n1082), .S(n1099) );
  CMPR32X1 U1120 ( .A(n1091), .B(n1090), .C(n1089), .CO(n1058), .S(n1104) );
  CMPR32X1 U1121 ( .A(n1094), .B(n1093), .C(n1092), .CO(n1103), .S(n1105) );
  CMPR32X1 U1122 ( .A(n1097), .B(n1096), .C(n1095), .CO(n1087), .S(n1102) );
  CMPR32X1 U1123 ( .A(n1104), .B(n1103), .C(n1102), .CO(n1098), .S(n1109) );
  CMPR32X1 U1124 ( .A(n1107), .B(n1106), .C(n1105), .CO(n1108), .S(n438) );
  NAND2XL U1125 ( .A(n1111), .B(n1110), .Y(n1112) );
  OAI21XL U1126 ( .A0(n1178), .A1(n1175), .B0(n1176), .Y(n1118) );
  OAI21XL U1127 ( .A0(n1121), .A1(n1120), .B0(n1119), .Y(n1126) );
  INVXL U1128 ( .A(n1122), .Y(n1124) );
  NAND2XL U1129 ( .A(n1124), .B(n1123), .Y(n1125) );
  XNOR2X1 U1130 ( .A(n1126), .B(n1125), .Y(PRODUCT[16]) );
  OAI21XL U1131 ( .A0(n1171), .A1(n1130), .B0(n1129), .Y(n1133) );
  CMPR32X1 U1132 ( .A(n1136), .B(n1135), .C(n1134), .CO(n1145), .S(n959) );
  CMPR32X1 U1133 ( .A(n1139), .B(n1138), .C(n1137), .CO(n899), .S(n1144) );
  CMPR32X1 U1134 ( .A(n1142), .B(n1141), .C(n1140), .CO(n1143), .S(n963) );
  CMPR32X1 U1135 ( .A(n1145), .B(n1144), .C(n1143), .CO(mult_x_1_n699), .S(
        mult_x_1_n700) );
  INVXL U1136 ( .A(n1146), .Y(n1188) );
  AOI21XL U1137 ( .A0(n1188), .A1(n1186), .B0(n1147), .Y(n1151) );
  CMPR32X1 U1138 ( .A(n1154), .B(n1153), .C(n1152), .CO(n897), .S(
        mult_x_1_n702) );
  NAND2XL U1139 ( .A(n1165), .B(n1161), .Y(n1163) );
  OAI21XL U1140 ( .A0(n1225), .A1(n1228), .B0(n1226), .Y(n1166) );
  OAI21XL U1141 ( .A0(n1171), .A1(n1163), .B0(n1162), .Y(n1164) );
  OAI21XL U1142 ( .A0(n1171), .A1(n1170), .B0(n1169), .Y(n1174) );
  XOR2XL U1143 ( .A(n1239), .B(n1237), .Y(PRODUCT[9]) );
  INVXL U1144 ( .A(n1235), .Y(n1180) );
  NAND2XL U1145 ( .A(n1180), .B(n1236), .Y(n1181) );
  OAI21XL U1146 ( .A0(n1182), .A1(n1235), .B0(n1236), .Y(n1185) );
  INVXL U1147 ( .A(n1233), .Y(n1183) );
  CMPR32X1 U1148 ( .A(n1191), .B(n1190), .C(n1189), .CO(n1200), .S(n901) );
  CMPR32X1 U1149 ( .A(n1194), .B(n1193), .C(n1192), .CO(n1199), .S(n900) );
  CMPR32X1 U1150 ( .A(n1197), .B(n1196), .C(n1195), .CO(n843), .S(n1198) );
  CMPR32X1 U1151 ( .A(n1200), .B(n1199), .C(n1198), .CO(mult_x_1_n669), .S(
        mult_x_1_n670) );
endmodule


module FFT2048_DW02_mult_2_stage_J1_11 ( A, B, TC, CLK, PRODUCT );
  input [25:0] A;
  input [16:0] B;
  output [42:0] PRODUCT;
  input TC, CLK;
  wire   n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         mult_x_1_n725, mult_x_1_n712, mult_x_1_n711, mult_x_1_n699,
         mult_x_1_n698, mult_x_1_n697, mult_x_1_n686, mult_x_1_n684,
         mult_x_1_n683, mult_x_1_n670, mult_x_1_n669, mult_x_1_n668,
         mult_x_1_n667, mult_x_1_n653, mult_x_1_n652, mult_x_1_n651,
         mult_x_1_n637, mult_x_1_n636, mult_x_1_n635, mult_x_1_n621,
         mult_x_1_n620, mult_x_1_n619, mult_x_1_n605, mult_x_1_n604,
         mult_x_1_n603, mult_x_1_n589, mult_x_1_n588, mult_x_1_n587,
         mult_x_1_n573, mult_x_1_n572, mult_x_1_n571, mult_x_1_n557,
         mult_x_1_n556, mult_x_1_n555, mult_x_1_n540, mult_x_1_n539,
         mult_x_1_n528, mult_x_1_n525, mult_x_1_n524, mult_x_1_n523,
         mult_x_1_n513, mult_x_1_n510, mult_x_1_n509, mult_x_1_n496,
         mult_x_1_n495, mult_x_1_n486, mult_x_1_n484, mult_x_1_n483,
         mult_x_1_n474, mult_x_1_n472, mult_x_1_n460, mult_x_1_n459,
         mult_x_1_n450, mult_x_1_n449, mult_x_1_n442, mult_x_1_n338,
         mult_x_1_n331, mult_x_1_n329, mult_x_1_n328, mult_x_1_n326,
         mult_x_1_n325, mult_x_1_n320, mult_x_1_n319, mult_x_1_n315,
         mult_x_1_n314, mult_x_1_n307, mult_x_1_n306, mult_x_1_n152,
         mult_x_1_n151, mult_x_1_n137, mult_x_1_n136, mult_x_1_n130,
         mult_x_1_n129, mult_x_1_n121, mult_x_1_n120, mult_x_1_n89,
         mult_x_1_n59, n6, n8, n9, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308;

  DFFHQXL mult_x_1_clk_r_REG24_S1 ( .D(mult_x_1_n151), .CK(CLK), .Q(n1239) );
  DFFHQX4 mult_x_1_clk_r_REG63_S1 ( .D(mult_x_1_n725), .CK(CLK), .Q(n1308) );
  DFFHQX4 mult_x_1_clk_r_REG62_S1 ( .D(mult_x_1_n712), .CK(CLK), .Q(n1307) );
  DFFHQX2 mult_x_1_clk_r_REG59_S1 ( .D(mult_x_1_n683), .CK(CLK), .Q(n1300) );
  DFFHQX2 mult_x_1_clk_r_REG50_S1 ( .D(mult_x_1_n667), .CK(CLK), .Q(n1296) );
  DFFHQX1 mult_x_1_clk_r_REG36_S1 ( .D(mult_x_1_n588), .CK(CLK), .Q(n1282) );
  DFFHQX4 mult_x_1_clk_r_REG32_S1 ( .D(mult_x_1_n571), .CK(CLK), .Q(n1278) );
  DFFHQXL mult_x_1_clk_r_REG25_S1 ( .D(mult_x_1_n137), .CK(CLK), .Q(n1238) );
  DFFHQXL mult_x_1_clk_r_REG20_S1 ( .D(mult_x_1_n449), .CK(CLK), .Q(n1255) );
  DFFHQXL mult_x_1_clk_r_REG11_S1 ( .D(mult_x_1_n495), .CK(CLK), .Q(n1264) );
  DFFHQXL mult_x_1_clk_r_REG21_S1 ( .D(mult_x_1_n450), .CK(CLK), .Q(n1256) );
  DFFHQXL mult_x_1_clk_r_REG3_S1 ( .D(mult_x_1_n540), .CK(CLK), .Q(n1274) );
  DFFHQXL mult_x_1_clk_r_REG8_S1 ( .D(mult_x_1_n509), .CK(CLK), .Q(n1266) );
  DFFHQXL mult_x_1_clk_r_REG22_S1 ( .D(mult_x_1_n442), .CK(CLK), .Q(n1254) );
  DFFHQXL mult_x_1_clk_r_REG61_S1 ( .D(mult_x_1_n711), .CK(CLK), .Q(n1306) );
  DFFHQXL mult_x_1_clk_r_REG17_S1 ( .D(mult_x_1_n459), .CK(CLK), .Q(n1257) );
  DFFHQXL mult_x_1_clk_r_REG9_S1 ( .D(mult_x_1_n510), .CK(CLK), .Q(n1267) );
  DFFHQXL mult_x_1_clk_r_REG33_S1 ( .D(mult_x_1_n572), .CK(CLK), .Q(n1279) );
  DFFHQXL mult_x_1_clk_r_REG45_S1 ( .D(mult_x_1_n636), .CK(CLK), .Q(n1291) );
  DFFHQXL mult_x_1_clk_r_REG23_S1 ( .D(mult_x_1_n152), .CK(CLK), .Q(n1240) );
  DFFHQXL mult_x_1_clk_r_REG64_S1 ( .D(mult_x_1_n307), .CK(CLK), .Q(n1242) );
  DFFHQXL mult_x_1_clk_r_REG57_S1 ( .D(mult_x_1_n697), .CK(CLK), .Q(n1303) );
  DFFHQXL clk_r_REG76_S1 ( .D(n1321), .CK(CLK), .Q(PRODUCT[8]) );
  DFFHQXL mult_x_1_clk_r_REG58_S1 ( .D(mult_x_1_n698), .CK(CLK), .Q(n1304) );
  DFFHQXL mult_x_1_clk_r_REG28_S1 ( .D(mult_x_1_n129), .CK(CLK), .Q(n1235) );
  DFFHQXL mult_x_1_clk_r_REG26_S1 ( .D(mult_x_1_n136), .CK(CLK), .Q(n1237) );
  DFFHQX1 mult_x_1_clk_r_REG39_S1 ( .D(mult_x_1_n604), .CK(CLK), .Q(n1285) );
  DFFHQX1 mult_x_1_clk_r_REG48_S1 ( .D(mult_x_1_n652), .CK(CLK), .Q(n1294) );
  DFFHQXL mult_x_1_clk_r_REG1_S1 ( .D(mult_x_1_n556), .CK(CLK), .Q(n1276) );
  DFFHQXL clk_r_REG78_S1 ( .D(n1322), .CK(CLK), .Q(PRODUCT[7]) );
  DFFHQXL clk_r_REG79_S1 ( .D(n1323), .CK(CLK), .Q(PRODUCT[6]) );
  DFFHQXL clk_r_REG80_S1 ( .D(n1324), .CK(CLK), .Q(PRODUCT[5]) );
  DFFHQXL clk_r_REG81_S1 ( .D(n1325), .CK(CLK), .Q(PRODUCT[4]) );
  DFFHQXL clk_r_REG82_S1 ( .D(n1326), .CK(CLK), .Q(PRODUCT[3]) );
  DFFHQXL clk_r_REG83_S1 ( .D(n1327), .CK(CLK), .Q(PRODUCT[2]) );
  DFFHQXL clk_r_REG84_S1 ( .D(n1328), .CK(CLK), .Q(PRODUCT[1]) );
  DFFHQXL clk_r_REG85_S1 ( .D(n1329), .CK(CLK), .Q(PRODUCT[0]) );
  DFFHQXL mult_x_1_clk_r_REG65_S1 ( .D(mult_x_1_n306), .CK(CLK), .Q(n1241) );
  DFFHQXL mult_x_1_clk_r_REG60_S1 ( .D(mult_x_1_n684), .CK(CLK), .Q(n1301) );
  DFFHQX2 mult_x_1_clk_r_REG54_S1 ( .D(mult_x_1_n669), .CK(CLK), .Q(n1298) );
  DFFHQX1 mult_x_1_clk_r_REG52_S1 ( .D(mult_x_1_n653), .CK(CLK), .Q(n1295) );
  DFFHQX2 mult_x_1_clk_r_REG49_S1 ( .D(mult_x_1_n637), .CK(CLK), .Q(n1292) );
  DFFHQX1 mult_x_1_clk_r_REG44_S1 ( .D(mult_x_1_n635), .CK(CLK), .Q(n1290) );
  DFFHQX2 mult_x_1_clk_r_REG46_S1 ( .D(mult_x_1_n621), .CK(CLK), .Q(n1289) );
  DFFHQXL mult_x_1_clk_r_REG42_S1 ( .D(mult_x_1_n620), .CK(CLK), .Q(n1288) );
  DFFHQX1 mult_x_1_clk_r_REG41_S1 ( .D(mult_x_1_n619), .CK(CLK), .Q(n1287) );
  DFFHQX1 mult_x_1_clk_r_REG38_S1 ( .D(mult_x_1_n603), .CK(CLK), .Q(n1284) );
  DFFHQX1 mult_x_1_clk_r_REG40_S1 ( .D(mult_x_1_n589), .CK(CLK), .Q(n1283) );
  DFFHQX1 mult_x_1_clk_r_REG35_S1 ( .D(mult_x_1_n587), .CK(CLK), .Q(n1281) );
  DFFHQX2 mult_x_1_clk_r_REG37_S1 ( .D(mult_x_1_n573), .CK(CLK), .Q(n1280) );
  DFFHQX1 mult_x_1_clk_r_REG34_S1 ( .D(mult_x_1_n557), .CK(CLK), .Q(n1277) );
  DFFHQX1 mult_x_1_clk_r_REG0_S1 ( .D(mult_x_1_n555), .CK(CLK), .Q(n1275) );
  DFFHQX1 mult_x_1_clk_r_REG2_S1 ( .D(mult_x_1_n539), .CK(CLK), .Q(n1273) );
  DFFHQX1 mult_x_1_clk_r_REG7_S1 ( .D(mult_x_1_n528), .CK(CLK), .Q(n1272) );
  DFFHQX1 mult_x_1_clk_r_REG6_S1 ( .D(mult_x_1_n525), .CK(CLK), .Q(n1271) );
  DFFHQXL mult_x_1_clk_r_REG5_S1 ( .D(mult_x_1_n524), .CK(CLK), .Q(n1270) );
  DFFHQXL mult_x_1_clk_r_REG4_S1 ( .D(mult_x_1_n523), .CK(CLK), .Q(n1269) );
  DFFHQX1 mult_x_1_clk_r_REG10_S1 ( .D(mult_x_1_n513), .CK(CLK), .Q(n1268) );
  DFFHQX1 mult_x_1_clk_r_REG15_S1 ( .D(mult_x_1_n486), .CK(CLK), .Q(n1263) );
  DFFHQXL mult_x_1_clk_r_REG16_S1 ( .D(mult_x_1_n472), .CK(CLK), .Q(n1259) );
  DFFHQXL mult_x_1_clk_r_REG18_S1 ( .D(mult_x_1_n460), .CK(CLK), .Q(n1258) );
  DFFHQXL mult_x_1_clk_r_REG77_S1 ( .D(mult_x_1_n338), .CK(CLK), .Q(n1253) );
  DFFHQXL mult_x_1_clk_r_REG75_S1 ( .D(mult_x_1_n331), .CK(CLK), .Q(n1252) );
  DFFHQXL mult_x_1_clk_r_REG74_S1 ( .D(mult_x_1_n89), .CK(CLK), .Q(n1251) );
  DFFHQX1 mult_x_1_clk_r_REG72_S1 ( .D(mult_x_1_n329), .CK(CLK), .Q(n1250) );
  DFFHQX1 mult_x_1_clk_r_REG73_S1 ( .D(mult_x_1_n328), .CK(CLK), .Q(n1249) );
  DFFHQX1 mult_x_1_clk_r_REG71_S1 ( .D(mult_x_1_n325), .CK(CLK), .Q(n1247) );
  DFFHQXL mult_x_1_clk_r_REG68_S1 ( .D(mult_x_1_n320), .CK(CLK), .Q(n1246) );
  DFFHQXL mult_x_1_clk_r_REG66_S1 ( .D(mult_x_1_n315), .CK(CLK), .Q(n1244) );
  DFFHQXL mult_x_1_clk_r_REG27_S1 ( .D(mult_x_1_n130), .CK(CLK), .Q(n1236) );
  DFFHQXL mult_x_1_clk_r_REG29_S1 ( .D(mult_x_1_n121), .CK(CLK), .Q(n1234) );
  DFFHQXL mult_x_1_clk_r_REG30_S1 ( .D(mult_x_1_n120), .CK(CLK), .Q(n1233) );
  DFFHQXL mult_x_1_clk_r_REG31_S1 ( .D(mult_x_1_n59), .CK(CLK), .Q(n1232) );
  DFFHQXL mult_x_1_clk_r_REG19_S1 ( .D(mult_x_1_n474), .CK(CLK), .Q(n1260) );
  DFFHQXL mult_x_1_clk_r_REG13_S1 ( .D(mult_x_1_n483), .CK(CLK), .Q(n1261) );
  DFFHQXL mult_x_1_clk_r_REG69_S1 ( .D(mult_x_1_n319), .CK(CLK), .Q(n1245) );
  DFFHQX1 mult_x_1_clk_r_REG47_S1 ( .D(mult_x_1_n651), .CK(CLK), .Q(n1293) );
  DFFHQXL mult_x_1_clk_r_REG51_S1 ( .D(mult_x_1_n668), .CK(CLK), .Q(n1297) );
  DFFHQXL mult_x_1_clk_r_REG70_S1 ( .D(mult_x_1_n326), .CK(CLK), .Q(n1248) );
  DFFHQXL mult_x_1_clk_r_REG67_S1 ( .D(mult_x_1_n314), .CK(CLK), .Q(n1243) );
  DFFHQX1 mult_x_1_clk_r_REG43_S1 ( .D(mult_x_1_n605), .CK(CLK), .Q(n1286) );
  DFFHQX1 mult_x_1_clk_r_REG53_S1 ( .D(mult_x_1_n686), .CK(CLK), .Q(n1302) );
  DFFHQX1 mult_x_1_clk_r_REG56_S1 ( .D(mult_x_1_n699), .CK(CLK), .Q(n1305) );
  DFFHQX2 mult_x_1_clk_r_REG55_S1 ( .D(mult_x_1_n670), .CK(CLK), .Q(n1299) );
  DFFHQX1 mult_x_1_clk_r_REG14_S1 ( .D(mult_x_1_n484), .CK(CLK), .Q(n1262) );
  DFFHQX1 mult_x_1_clk_r_REG12_S1 ( .D(mult_x_1_n496), .CK(CLK), .Q(n1265) );
  ADDFHX1 U1 ( .A(n987), .B(n986), .CI(n985), .CO(mult_x_1_n697), .S(
        mult_x_1_n698) );
  ADDFHX1 U2 ( .A(n990), .B(n989), .CI(n988), .CO(mult_x_1_n699), .S(n985) );
  ADDFHX1 U3 ( .A(n999), .B(n998), .CI(n997), .CO(n986), .S(n1000) );
  ADDFHX1 U4 ( .A(n996), .B(n995), .CI(n994), .CO(n1001), .S(n1003) );
  CMPR32X1 U5 ( .A(n532), .B(n531), .C(n530), .CO(n94), .S(n533) );
  NAND2X4 U6 ( .A(n66), .B(n974), .Y(n832) );
  BUFX4 U7 ( .A(n71), .Y(n1054) );
  NAND2X1 U8 ( .A(n65), .B(n335), .Y(n1011) );
  BUFX3 U9 ( .A(n901), .Y(n934) );
  NAND2X4 U10 ( .A(n68), .B(n901), .Y(n828) );
  INVX1 U11 ( .A(B[12]), .Y(n61) );
  XOR2X1 U12 ( .A(B[14]), .B(B[15]), .Y(n70) );
  NAND2X1 U13 ( .A(n543), .B(n40), .Y(n970) );
  BUFX3 U14 ( .A(n410), .Y(n8) );
  INVX1 U15 ( .A(B[9]), .Y(n471) );
  CLKBUFX3 U16 ( .A(B[1]), .Y(n612) );
  XNOR2X1 U17 ( .A(B[6]), .B(B[5]), .Y(n901) );
  OAI21XL U18 ( .A0(n203), .A1(n154), .B0(n153), .Y(n1177) );
  XNOR2X2 U19 ( .A(n231), .B(n230), .Y(PRODUCT[30]) );
  NAND2X1 U20 ( .A(n116), .B(n115), .Y(n297) );
  ADDFHX2 U21 ( .A(n1295), .B(n1293), .CI(n1291), .CO(n115), .S(n110) );
  ADDFHX1 U22 ( .A(n1298), .B(n1296), .CI(n1294), .CO(n109), .S(n108) );
  ADDFHX1 U23 ( .A(n1299), .B(n1300), .CI(n1297), .CO(n107), .S(n106) );
  OAI22X1 U24 ( .A0(n951), .A1(n949), .B0(n882), .B1(n1006), .Y(n966) );
  OAI21XL U25 ( .A0(n304), .A1(n310), .B0(n305), .Y(n111) );
  ADDFX2 U26 ( .A(n1260), .B(n1261), .CI(n1259), .CO(n146), .S(n145) );
  XOR2XL U27 ( .A(n313), .B(n312), .Y(PRODUCT[19]) );
  XNOR2XL U28 ( .A(n329), .B(n328), .Y(PRODUCT[15]) );
  XOR2XL U29 ( .A(n6), .B(n888), .Y(n34) );
  XNOR2XL U30 ( .A(n9), .B(n905), .Y(n369) );
  INVX1 U31 ( .A(n1054), .Y(n30) );
  XNOR2XL U32 ( .A(B[16]), .B(n884), .Y(n676) );
  XNOR2XL U33 ( .A(n9), .B(n898), .Y(n784) );
  XNOR2XL U34 ( .A(n9), .B(n1051), .Y(n1009) );
  XNOR2XL U35 ( .A(n900), .B(n889), .Y(n391) );
  XNOR2XL U36 ( .A(n9), .B(n850), .Y(n648) );
  XNOR2XL U37 ( .A(B[16]), .B(n889), .Y(n765) );
  CLKINVX2 U38 ( .A(B[15]), .Y(n953) );
  XNOR2XL U39 ( .A(n9), .B(n888), .Y(n339) );
  XNOR2XL U40 ( .A(n1049), .B(n850), .Y(n503) );
  XNOR2XL U41 ( .A(n1049), .B(n893), .Y(n569) );
  XNOR2XL U42 ( .A(n1027), .B(n852), .Y(n679) );
  XOR2X1 U43 ( .A(B[7]), .B(n41), .Y(n543) );
  XNOR2X2 U44 ( .A(B[2]), .B(B[1]), .Y(n926) );
  XNOR2XL U45 ( .A(n1151), .B(n1150), .Y(n1322) );
  XNOR2X1 U46 ( .A(n1228), .B(n55), .Y(n1321) );
  NAND2X1 U47 ( .A(n499), .B(n1227), .Y(n55) );
  INVXL U48 ( .A(n498), .Y(n1228) );
  OAI21XL U49 ( .A0(n37), .A1(n36), .B0(n35), .Y(mult_x_1_n449) );
  NAND2X1 U50 ( .A(n94), .B(n95), .Y(n35) );
  NOR2X1 U51 ( .A(n94), .B(n95), .Y(n37) );
  XNOR2X1 U52 ( .A(n93), .B(n39), .Y(n38) );
  INVX1 U53 ( .A(n93), .Y(n36) );
  INVXL U54 ( .A(n491), .Y(n56) );
  NAND2XL U55 ( .A(n25), .B(n24), .Y(n1043) );
  NAND2XL U56 ( .A(n29), .B(n27), .Y(n1107) );
  OR2XL U57 ( .A(n629), .B(n628), .Y(n601) );
  OAI21XL U58 ( .A0(n904), .A1(n74), .B0(n22), .Y(n83) );
  INVXL U59 ( .A(n52), .Y(n50) );
  NAND2BXL U60 ( .AN(n1024), .B(n30), .Y(n26) );
  NAND2XL U61 ( .A(n32), .B(n34), .Y(n31) );
  NAND2BXL U62 ( .AN(n85), .B(n30), .Y(n22) );
  NAND2BXL U63 ( .AN(n180), .B(n28), .Y(n18) );
  NAND2BX1 U64 ( .AN(n174), .B(n30), .Y(n21) );
  NAND2BX1 U65 ( .AN(n85), .B(n28), .Y(n20) );
  NOR2X1 U66 ( .A(n519), .B(n906), .Y(n1194) );
  NAND2BXL U67 ( .AN(n913), .B(n34), .Y(n33) );
  NAND2BXL U68 ( .AN(n1040), .B(n28), .Y(n27) );
  NAND2BXL U69 ( .AN(n1055), .B(n30), .Y(n29) );
  NAND2BXL U70 ( .AN(n1024), .B(n28), .Y(n24) );
  NAND2BXL U71 ( .AN(n1040), .B(n30), .Y(n25) );
  INVX1 U72 ( .A(n968), .Y(n32) );
  XNOR2X1 U73 ( .A(n308), .B(n307), .Y(PRODUCT[20]) );
  INVXL U74 ( .A(n901), .Y(n54) );
  XOR2X1 U75 ( .A(n320), .B(n319), .Y(PRODUCT[18]) );
  NOR2BXL U76 ( .AN(n402), .B(n901), .Y(n414) );
  XNOR2X1 U77 ( .A(n1128), .B(n1127), .Y(PRODUCT[16]) );
  NOR2X1 U78 ( .A(n204), .B(n205), .Y(n195) );
  BUFX2 U79 ( .A(A[4]), .Y(n889) );
  NOR2X1 U80 ( .A(n204), .B(n154), .Y(n1174) );
  AOI21XL U81 ( .A0(n134), .A1(n241), .B0(n133), .Y(n135) );
  NAND2X1 U82 ( .A(n234), .B(n233), .Y(n235) );
  NAND2X1 U83 ( .A(n257), .B(n256), .Y(n258) );
  NAND2X1 U84 ( .A(n266), .B(n265), .Y(n267) );
  NOR2X1 U85 ( .A(n146), .B(n1258), .Y(n215) );
  NAND2X1 U86 ( .A(n126), .B(n125), .Y(n271) );
  INVX1 U87 ( .A(n1243), .Y(n1143) );
  ADDFHX1 U88 ( .A(n1283), .B(n1281), .CI(n1279), .CO(n125), .S(n122) );
  ADDFHX1 U89 ( .A(n1292), .B(n1290), .CI(n1288), .CO(n117), .S(n116) );
  INVX1 U90 ( .A(n499), .Y(n1226) );
  XOR2X1 U91 ( .A(n38), .B(n94), .Y(mult_x_1_n450) );
  NOR2X1 U92 ( .A(n455), .B(n454), .Y(n1147) );
  NAND2X1 U93 ( .A(n453), .B(n452), .Y(n1163) );
  NOR2X1 U94 ( .A(n453), .B(n452), .Y(n1162) );
  XOR2X1 U95 ( .A(n480), .B(n51), .Y(n488) );
  XNOR2X1 U96 ( .A(n158), .B(n157), .Y(PRODUCT[36]) );
  XNOR2X1 U97 ( .A(n1161), .B(n1160), .Y(PRODUCT[37]) );
  NAND2X1 U98 ( .A(n21), .B(n20), .Y(n170) );
  OAI21XL U99 ( .A0(n343), .A1(n968), .B0(n33), .Y(n388) );
  XNOR2X1 U100 ( .A(n283), .B(n282), .Y(PRODUCT[24]) );
  NAND2BX1 U101 ( .AN(n972), .B(n28), .Y(n12) );
  NOR2X1 U102 ( .A(n519), .B(n616), .Y(n673) );
  NOR2X1 U103 ( .A(n519), .B(n765), .Y(n792) );
  NAND2BX1 U104 ( .AN(n767), .B(n28), .Y(n14) );
  NOR2X1 U105 ( .A(n519), .B(n676), .Y(n702) );
  NOR2X1 U106 ( .A(n519), .B(n705), .Y(n731) );
  NOR2X1 U107 ( .A(n519), .B(n614), .Y(n626) );
  NOR2X1 U108 ( .A(n519), .B(n796), .Y(n821) );
  NAND2BXL U109 ( .AN(n1055), .B(n28), .Y(n19) );
  NOR2X1 U110 ( .A(n519), .B(n862), .Y(n914) );
  NOR2X1 U111 ( .A(n519), .B(n826), .Y(n858) );
  OR2XL U112 ( .A(n426), .B(n425), .Y(n1219) );
  NAND2X1 U113 ( .A(n332), .B(n333), .Y(n410) );
  CLKINVX8 U114 ( .A(n471), .Y(n6) );
  BUFX2 U115 ( .A(A[5]), .Y(n896) );
  NAND2XL U116 ( .A(n269), .B(n272), .Y(n263) );
  BUFX2 U117 ( .A(A[19]), .Y(n763) );
  BUFX2 U118 ( .A(A[16]), .Y(n860) );
  BUFX2 U119 ( .A(A[21]), .Y(n1025) );
  BUFX2 U120 ( .A(A[18]), .Y(n794) );
  BUFX2 U121 ( .A(A[20]), .Y(n1007) );
  INVXL U122 ( .A(n402), .Y(n47) );
  BUFX2 U123 ( .A(A[23]), .Y(n1048) );
  BUFX2 U124 ( .A(A[13]), .Y(n885) );
  BUFX3 U125 ( .A(A[0]), .Y(n402) );
  NOR2X1 U126 ( .A(n128), .B(n127), .Y(n264) );
  NOR2X1 U127 ( .A(n130), .B(n129), .Y(n237) );
  NOR2X1 U128 ( .A(n122), .B(n121), .Y(n279) );
  NOR2X1 U129 ( .A(n143), .B(n142), .Y(n227) );
  NOR2X1 U130 ( .A(n1257), .B(n1256), .Y(n205) );
  ADDFHX1 U131 ( .A(n1272), .B(n1273), .CI(n1270), .CO(n131), .S(n130) );
  ADDFHX1 U132 ( .A(n1277), .B(n1275), .CI(n1274), .CO(n129), .S(n128) );
  OR2X2 U133 ( .A(n494), .B(n493), .Y(n484) );
  NAND2BX1 U134 ( .AN(n492), .B(n56), .Y(n1227) );
  NAND2XL U135 ( .A(n58), .B(n57), .Y(mult_x_1_n725) );
  OR2XL U136 ( .A(n1064), .B(n1063), .Y(n1066) );
  INVX1 U137 ( .A(n95), .Y(n39) );
  OAI2BB1XL U138 ( .A0N(n480), .A1N(n52), .B0(n48), .Y(n486) );
  OAI2BB1XL U139 ( .A0N(n43), .A1N(n965), .B0(n42), .Y(n1134) );
  NAND2XL U140 ( .A(n49), .B(n479), .Y(n48) );
  NAND2BXL U141 ( .AN(n480), .B(n50), .Y(n49) );
  XOR2X1 U142 ( .A(n965), .B(n45), .Y(n1130) );
  XOR2X1 U143 ( .A(n966), .B(n46), .Y(n45) );
  XOR2X1 U144 ( .A(n479), .B(n52), .Y(n51) );
  OAI21XL U145 ( .A0(n904), .A1(n1014), .B0(n26), .Y(n1030) );
  OAI21XL U146 ( .A0(n390), .A1(n970), .B0(n31), .Y(n1071) );
  NAND2BX1 U147 ( .AN(n570), .B(n28), .Y(n11) );
  AND2XL U148 ( .A(n1225), .B(n1224), .Y(n1328) );
  OR2X2 U149 ( .A(n442), .B(n441), .Y(n440) );
  XNOR2XL U150 ( .A(n1049), .B(n1048), .Y(n1050) );
  OR2XL U151 ( .A(n1223), .B(n1222), .Y(n1225) );
  XNOR2XL U152 ( .A(n1049), .B(A[22]), .Y(n1044) );
  NAND2BX1 U153 ( .AN(n475), .B(n54), .Y(n53) );
  XNOR2XL U154 ( .A(n1049), .B(n1007), .Y(n1008) );
  NAND2BXL U155 ( .AN(A[0]), .B(n1052), .Y(n952) );
  XNOR2XL U156 ( .A(n1052), .B(n1051), .Y(n1053) );
  CLKINVX8 U157 ( .A(n345), .Y(n9) );
  INVX1 U158 ( .A(B[8]), .Y(n41) );
  XNOR2X1 U159 ( .A(B[4]), .B(B[3]), .Y(n333) );
  BUFX2 U160 ( .A(A[25]), .Y(n1051) );
  BUFX2 U161 ( .A(A[12]), .Y(n852) );
  BUFX2 U162 ( .A(A[11]), .Y(n893) );
  BUFX2 U163 ( .A(A[6]), .Y(n848) );
  BUFX2 U164 ( .A(A[9]), .Y(n898) );
  BUFX2 U165 ( .A(A[10]), .Y(n899) );
  BUFX2 U166 ( .A(A[1]), .Y(n905) );
  BUFX2 U167 ( .A(A[14]), .Y(n850) );
  BUFX2 U168 ( .A(A[7]), .Y(n884) );
  BUFX2 U169 ( .A(A[15]), .Y(n881) );
  INVXL U170 ( .A(n246), .Y(n248) );
  INVXL U171 ( .A(n309), .Y(n311) );
  NAND2XL U172 ( .A(n207), .B(n206), .Y(n208) );
  INVXL U173 ( .A(n327), .Y(n62) );
  AND2XL U174 ( .A(n1176), .B(n1181), .Y(n1170) );
  ADDFHX2 U175 ( .A(n1302), .B(n1305), .CI(n1301), .CO(n105), .S(n104) );
  OAI21XL U176 ( .A0(n971), .A1(n1054), .B0(n12), .Y(n980) );
  OAI22X1 U177 ( .A0(n928), .A1(n408), .B0(n926), .B1(n462), .Y(n480) );
  XOR2X1 U178 ( .A(B[2]), .B(B[3]), .Y(n331) );
  AOI21X1 U179 ( .A0(n484), .A1(n1226), .B0(n495), .Y(n496) );
  NAND2X1 U180 ( .A(n492), .B(n491), .Y(n499) );
  CLKBUFX8 U181 ( .A(B[16]), .Y(n1049) );
  CLKINVX2 U182 ( .A(B[11]), .Y(n345) );
  NOR2X1 U183 ( .A(n519), .B(n520), .Y(n554) );
  OAI22X1 U184 ( .A0(n932), .A1(n929), .B0(n930), .B1(n897), .Y(n941) );
  OAI22X1 U185 ( .A0(n952), .A1(n1054), .B0(n904), .B1(n953), .Y(n963) );
  OAI22X1 U186 ( .A0(n548), .A1(n904), .B0(n1054), .B1(n522), .Y(n557) );
  OAI21XL U187 ( .A0(n1054), .A1(n548), .B0(n11), .Y(n572) );
  OAI22X1 U188 ( .A0(n514), .A1(n1054), .B0(n904), .B1(n522), .Y(n528) );
  OAI21XL U189 ( .A0(n707), .A1(n1054), .B0(n13), .Y(n739) );
  NAND2BX1 U190 ( .AN(n736), .B(n28), .Y(n13) );
  OAI21XL U191 ( .A0(n736), .A1(n1054), .B0(n14), .Y(n770) );
  OAI22X1 U192 ( .A0(n678), .A1(n904), .B0(n631), .B1(n1054), .Y(n681) );
  OAI21XL U193 ( .A0(n767), .A1(n1054), .B0(n15), .Y(n801) );
  NAND2BX1 U194 ( .AN(n798), .B(n28), .Y(n15) );
  OAI22X1 U195 ( .A0(n798), .A1(n1054), .B0(n829), .B1(n904), .Y(n834) );
  OAI21XL U196 ( .A0(n678), .A1(n1054), .B0(n16), .Y(n710) );
  NAND2BX1 U197 ( .AN(n707), .B(n28), .Y(n16) );
  OAI21XL U198 ( .A0(n74), .A1(n1054), .B0(n17), .Y(n508) );
  NAND2BX1 U199 ( .AN(n514), .B(n28), .Y(n17) );
  OAI21XL U200 ( .A0(n1014), .A1(n1054), .B0(n18), .Y(n1017) );
  OAI21XL U201 ( .A0(n1054), .A1(n1053), .B0(n19), .Y(n1056) );
  OAI21XL U202 ( .A0(n1054), .A1(n180), .B0(n23), .Y(n189) );
  NAND2BX1 U203 ( .AN(n174), .B(n28), .Y(n23) );
  CLKINVX3 U204 ( .A(n904), .Y(n28) );
  XOR2X1 U205 ( .A(B[9]), .B(B[8]), .Y(n40) );
  XNOR2X2 U206 ( .A(B[15]), .B(B[16]), .Y(n519) );
  NAND2XL U207 ( .A(n966), .B(n46), .Y(n42) );
  NAND2BX1 U208 ( .AN(n966), .B(n44), .Y(n43) );
  INVXL U209 ( .A(n46), .Y(n44) );
  NOR2X1 U210 ( .A(n519), .B(n47), .Y(n46) );
  OAI21XL U211 ( .A0(n406), .A1(n828), .B0(n53), .Y(n52) );
  NOR2X1 U212 ( .A(n275), .B(n279), .Y(n124) );
  INVX1 U213 ( .A(n238), .Y(n269) );
  NAND2X1 U214 ( .A(n124), .B(n284), .Y(n238) );
  NAND2XL U215 ( .A(n1004), .B(n1005), .Y(n57) );
  OAI21XL U216 ( .A0(n1004), .A1(n1005), .B0(n1003), .Y(n58) );
  XOR3X2 U217 ( .A(n1005), .B(n1003), .C(n1004), .Y(n382) );
  NOR2X1 U218 ( .A(n118), .B(n117), .Y(n292) );
  XNOR2X1 U219 ( .A(n1052), .B(n881), .Y(n522) );
  XNOR2X1 U220 ( .A(n1052), .B(n850), .Y(n548) );
  INVX2 U221 ( .A(n239), .Y(n300) );
  INVX1 U222 ( .A(n324), .Y(n301) );
  INVXL U223 ( .A(n1141), .Y(n1192) );
  XNOR2XL U224 ( .A(n1012), .B(n860), .Y(n551) );
  XNOR2X2 U225 ( .A(B[14]), .B(B[13]), .Y(n71) );
  OAI21XL U226 ( .A0(n227), .A1(n233), .B0(n228), .Y(n211) );
  XNOR2XL U227 ( .A(n612), .B(n899), .Y(n389) );
  XNOR2XL U228 ( .A(n612), .B(n898), .Y(n469) );
  INVXL U229 ( .A(n1241), .Y(n1119) );
  XNOR2XL U230 ( .A(n9), .B(A[24]), .Y(n182) );
  XNOR2XL U231 ( .A(n6), .B(n1051), .Y(n172) );
  XNOR2XL U232 ( .A(n9), .B(n1048), .Y(n176) );
  XNOR2XL U233 ( .A(n1052), .B(n763), .Y(n174) );
  XNOR2XL U234 ( .A(n900), .B(n883), .Y(n474) );
  XNOR2XL U235 ( .A(n900), .B(n1051), .Y(n77) );
  XNOR2XL U236 ( .A(n6), .B(A[24]), .Y(n87) );
  XNOR2XL U237 ( .A(n755), .B(A[24]), .Y(n547) );
  INVXL U238 ( .A(B[13]), .Y(n67) );
  XNOR2XL U239 ( .A(B[3]), .B(A[22]), .Y(n649) );
  XNOR2XL U240 ( .A(B[3]), .B(n1025), .Y(n667) );
  XNOR2XL U241 ( .A(B[3]), .B(n1007), .Y(n696) );
  XNOR2XL U242 ( .A(B[3]), .B(n763), .Y(n725) );
  XNOR2XL U243 ( .A(B[3]), .B(n794), .Y(n754) );
  XNOR2XL U244 ( .A(B[3]), .B(n823), .Y(n785) );
  XNOR2XL U245 ( .A(n612), .B(n860), .Y(n882) );
  XNOR2XL U246 ( .A(n612), .B(n881), .Y(n949) );
  XNOR2XL U247 ( .A(n1012), .B(n1048), .Y(n1013) );
  XNOR2XL U248 ( .A(n886), .B(n883), .Y(n436) );
  XNOR2XL U249 ( .A(n894), .B(n905), .Y(n419) );
  NAND2XL U250 ( .A(n294), .B(n293), .Y(n295) );
  AOI21XL U251 ( .A0(n239), .A1(n298), .B0(n60), .Y(n59) );
  XNOR2X1 U252 ( .A(n291), .B(n290), .Y(PRODUCT[23]) );
  NAND2XL U253 ( .A(n289), .B(n288), .Y(n290) );
  NAND2XL U254 ( .A(n272), .B(n271), .Y(n273) );
  NAND2XL U255 ( .A(n200), .B(n199), .Y(n201) );
  NAND2XL U256 ( .A(n162), .B(n1240), .Y(n163) );
  OAI21XL U257 ( .A0(n1180), .A1(n161), .B0(n160), .Y(n164) );
  INVXL U258 ( .A(n1177), .Y(n155) );
  INVXL U259 ( .A(n1238), .Y(n1155) );
  NAND2XL U260 ( .A(n327), .B(n326), .Y(n328) );
  XOR2XL U261 ( .A(n1145), .B(n1144), .Y(PRODUCT[13]) );
  NAND2XL U262 ( .A(n1143), .B(n1244), .Y(n1144) );
  INVXL U263 ( .A(n1059), .Y(n1041) );
  NOR2XL U264 ( .A(n519), .B(n1026), .Y(n1042) );
  XNOR2XL U265 ( .A(n6), .B(n1007), .Y(n550) );
  XNOR2XL U266 ( .A(n6), .B(n1025), .Y(n542) );
  NAND2X1 U267 ( .A(B[1]), .B(n330), .Y(n825) );
  NAND2X1 U268 ( .A(n331), .B(n926), .Y(n786) );
  BUFX3 U269 ( .A(n970), .Y(n913) );
  BUFX3 U270 ( .A(n333), .Y(n947) );
  NOR2XL U271 ( .A(n519), .B(n1044), .Y(n1058) );
  OAI2BB1XL U272 ( .A0N(n974), .A1N(n832), .B0(n1046), .Y(n1057) );
  NOR2X2 U273 ( .A(n110), .B(n109), .Y(n304) );
  NOR2XL U274 ( .A(n145), .B(n144), .Y(n210) );
  NOR2X1 U275 ( .A(n316), .B(n314), .Y(n303) );
  NOR2X1 U276 ( .A(n104), .B(n1303), .Y(n314) );
  NOR2X2 U277 ( .A(n106), .B(n105), .Y(n316) );
  INVXL U278 ( .A(n1252), .Y(n1186) );
  XNOR2XL U279 ( .A(n886), .B(n898), .Y(n371) );
  XNOR2XL U280 ( .A(n900), .B(n896), .Y(n368) );
  XNOR2XL U281 ( .A(n894), .B(n883), .Y(n407) );
  NOR2X1 U282 ( .A(n108), .B(n107), .Y(n309) );
  NAND2X1 U283 ( .A(n108), .B(n107), .Y(n310) );
  INVXL U284 ( .A(n227), .Y(n229) );
  NOR2X1 U285 ( .A(n141), .B(n140), .Y(n232) );
  NAND2X1 U286 ( .A(n141), .B(n140), .Y(n233) );
  INVXL U287 ( .A(n210), .Y(n224) );
  NAND2XL U288 ( .A(n220), .B(n148), .Y(n204) );
  NOR2XL U289 ( .A(n1237), .B(n1235), .Y(n1176) );
  INVXL U290 ( .A(n314), .Y(n322) );
  NAND2X1 U291 ( .A(n106), .B(n105), .Y(n317) );
  XNOR2XL U292 ( .A(n894), .B(n884), .Y(n372) );
  XNOR2XL U293 ( .A(n886), .B(A[8]), .Y(n393) );
  XNOR2XL U294 ( .A(n886), .B(n896), .Y(n462) );
  XNOR2XL U295 ( .A(n894), .B(n888), .Y(n464) );
  XNOR2XL U296 ( .A(n6), .B(n402), .Y(n460) );
  XNOR2XL U297 ( .A(n894), .B(n889), .Y(n463) );
  XNOR2XL U298 ( .A(n894), .B(n896), .Y(n461) );
  XNOR2XL U299 ( .A(n900), .B(n888), .Y(n458) );
  XNOR2XL U300 ( .A(n6), .B(n905), .Y(n459) );
  XNOR2XL U301 ( .A(n886), .B(n848), .Y(n468) );
  XNOR2XL U302 ( .A(n886), .B(n884), .Y(n467) );
  NAND2BXL U303 ( .AN(n402), .B(n6), .Y(n470) );
  OAI22XL U304 ( .A0(n951), .A1(n473), .B0(n472), .B1(n1006), .Y(n477) );
  NOR2BXL U305 ( .AN(n402), .B(n968), .Y(n478) );
  XNOR2XL U306 ( .A(n1052), .B(n794), .Y(n85) );
  XNOR2XL U307 ( .A(n612), .B(n1051), .Y(n613) );
  CLKINVX2 U308 ( .A(n504), .Y(n755) );
  XNOR2XL U309 ( .A(n755), .B(n1007), .Y(n650) );
  XNOR2XL U310 ( .A(n755), .B(n763), .Y(n668) );
  XNOR2XL U311 ( .A(n755), .B(n794), .Y(n697) );
  XNOR2XL U312 ( .A(n755), .B(n823), .Y(n726) );
  XNOR2XL U313 ( .A(n755), .B(n860), .Y(n756) );
  XNOR2XL U314 ( .A(n755), .B(n881), .Y(n787) );
  XNOR2XL U315 ( .A(n886), .B(n850), .Y(n887) );
  XNOR2XL U316 ( .A(n886), .B(n885), .Y(n925) );
  XNOR2X1 U317 ( .A(n1052), .B(n905), .Y(n971) );
  XNOR2XL U318 ( .A(n6), .B(n884), .Y(n967) );
  XNOR2XL U319 ( .A(n9), .B(n889), .Y(n931) );
  XNOR2XL U320 ( .A(n886), .B(n852), .Y(n927) );
  XNOR2XL U321 ( .A(n6), .B(n848), .Y(n969) );
  XNOR2XL U322 ( .A(n6), .B(n896), .Y(n334) );
  XNOR2XL U323 ( .A(n886), .B(n899), .Y(n363) );
  XNOR2XL U324 ( .A(n894), .B(A[8]), .Y(n364) );
  XNOR2XL U325 ( .A(n900), .B(n848), .Y(n362) );
  XNOR2XL U326 ( .A(n900), .B(A[8]), .Y(n935) );
  XNOR2XL U327 ( .A(n900), .B(n884), .Y(n352) );
  XNOR2XL U328 ( .A(n894), .B(n898), .Y(n351) );
  XNOR2XL U329 ( .A(n6), .B(n889), .Y(n343) );
  OAI22XL U330 ( .A0(n951), .A1(n389), .B0(n346), .B1(n1006), .Y(n374) );
  NAND2BXL U331 ( .AN(n402), .B(n9), .Y(n344) );
  OAI22XL U332 ( .A0(n951), .A1(n346), .B0(n354), .B1(n1006), .Y(n360) );
  NOR2BXL U333 ( .AN(n402), .B(n974), .Y(n361) );
  NAND2BXL U334 ( .AN(n402), .B(n1027), .Y(n355) );
  XNOR2XL U335 ( .A(n886), .B(n905), .Y(n437) );
  XNOR2XL U336 ( .A(n612), .B(n888), .Y(n435) );
  XNOR2XL U337 ( .A(n612), .B(n889), .Y(n434) );
  INVXL U338 ( .A(n900), .Y(n404) );
  INVXL U339 ( .A(n1174), .Y(n156) );
  INVXL U340 ( .A(n1237), .Y(n1156) );
  NAND2XL U341 ( .A(n1174), .B(n1156), .Y(n1158) );
  INVXL U342 ( .A(n1235), .Y(n1159) );
  INVXL U343 ( .A(n1168), .Y(n1169) );
  AOI21XL U344 ( .A0(n1175), .A1(n1181), .B0(n1167), .Y(n1168) );
  INVXL U345 ( .A(n1234), .Y(n1167) );
  INVXL U346 ( .A(n152), .Y(n153) );
  AOI21XL U347 ( .A0(n159), .A1(n162), .B0(n149), .Y(n150) );
  NAND2XL U348 ( .A(n1174), .B(n1176), .Y(n1179) );
  INVXL U349 ( .A(n1233), .Y(n1181) );
  NAND2XL U350 ( .A(n1126), .B(n1125), .Y(n1127) );
  XNOR2XL U351 ( .A(n1192), .B(n1191), .Y(PRODUCT[12]) );
  OAI22XL U352 ( .A0(n932), .A1(n176), .B0(n930), .B1(n182), .Y(n187) );
  OAI2BB1XL U353 ( .A0N(n968), .A1N(n913), .B0(n173), .Y(n184) );
  INVXL U354 ( .A(n172), .Y(n173) );
  XNOR2XL U355 ( .A(n9), .B(A[22]), .Y(n86) );
  XNOR2XL U356 ( .A(n6), .B(n1048), .Y(n73) );
  XNOR2XL U357 ( .A(n9), .B(n1025), .Y(n72) );
  OAI22XL U358 ( .A0(n832), .A1(n1013), .B0(n974), .B1(n1028), .Y(n1031) );
  CMPR32X1 U359 ( .A(n92), .B(n91), .C(n90), .CO(n165), .S(n531) );
  NOR2XL U360 ( .A(n519), .B(n76), .Y(n92) );
  INVXL U361 ( .A(n77), .Y(n78) );
  XNOR2XL U362 ( .A(n9), .B(n1007), .Y(n516) );
  XNOR2XL U363 ( .A(n900), .B(A[22]), .Y(n549) );
  XNOR2XL U364 ( .A(n9), .B(n794), .Y(n552) );
  XNOR2XL U365 ( .A(n9), .B(n763), .Y(n523) );
  XNOR2XL U366 ( .A(n900), .B(A[24]), .Y(n513) );
  XNOR2XL U367 ( .A(n6), .B(A[22]), .Y(n515) );
  XNOR2XL U368 ( .A(n886), .B(n1051), .Y(n545) );
  XNOR2X1 U369 ( .A(n1052), .B(n885), .Y(n570) );
  XNOR2XL U370 ( .A(n900), .B(n1025), .Y(n568) );
  XNOR2XL U371 ( .A(n900), .B(n1007), .Y(n590) );
  XNOR2XL U372 ( .A(n6), .B(n823), .Y(n625) );
  XNOR2XL U373 ( .A(n755), .B(n1025), .Y(n618) );
  INVXL U374 ( .A(n613), .Y(n584) );
  XNOR2XL U375 ( .A(B[3]), .B(n1048), .Y(n608) );
  XNOR2XL U376 ( .A(n755), .B(A[22]), .Y(n617) );
  XNOR2XL U377 ( .A(n755), .B(n1048), .Y(n586) );
  OAI22XL U378 ( .A0(n828), .A1(n630), .B0(n934), .B1(n590), .Y(n629) );
  XNOR2XL U379 ( .A(n9), .B(n860), .Y(n589) );
  XNOR2XL U380 ( .A(n6), .B(n794), .Y(n624) );
  XNOR2XL U381 ( .A(n6), .B(n763), .Y(n587) );
  XNOR2XL U382 ( .A(n900), .B(n763), .Y(n630) );
  XNOR2XL U383 ( .A(n6), .B(n860), .Y(n672) );
  XNOR2XL U384 ( .A(n6), .B(n881), .Y(n701) );
  OAI22XL U385 ( .A0(n951), .A1(n704), .B0(n675), .B1(n1006), .Y(n703) );
  XNOR2XL U386 ( .A(n900), .B(n794), .Y(n677) );
  XNOR2X1 U387 ( .A(n1052), .B(n899), .Y(n678) );
  XNOR2XL U388 ( .A(n6), .B(n850), .Y(n730) );
  XNOR2XL U389 ( .A(n900), .B(n823), .Y(n706) );
  XNOR2X1 U390 ( .A(n1052), .B(n898), .Y(n707) );
  XNOR2XL U391 ( .A(n6), .B(n885), .Y(n760) );
  OAI22XL U392 ( .A0(n825), .A1(n764), .B0(n733), .B1(n1006), .Y(n762) );
  XNOR2XL U393 ( .A(n900), .B(n860), .Y(n735) );
  XNOR2X1 U394 ( .A(n1052), .B(A[8]), .Y(n736) );
  XNOR2XL U395 ( .A(n6), .B(n852), .Y(n791) );
  XNOR2XL U396 ( .A(n900), .B(n881), .Y(n766) );
  XNOR2X1 U397 ( .A(n1052), .B(n884), .Y(n767) );
  XNOR2XL U398 ( .A(n6), .B(n893), .Y(n820) );
  OAI22XL U399 ( .A0(n825), .A1(n824), .B0(n795), .B1(n1006), .Y(n822) );
  XNOR2XL U400 ( .A(n900), .B(n850), .Y(n797) );
  XNOR2X1 U401 ( .A(n1052), .B(n848), .Y(n798) );
  XNOR2XL U402 ( .A(n6), .B(n899), .Y(n853) );
  XNOR2XL U403 ( .A(n894), .B(n850), .Y(n854) );
  XNOR2XL U404 ( .A(n894), .B(n885), .Y(n855) );
  XNOR2X1 U405 ( .A(n1052), .B(n896), .Y(n829) );
  XNOR2XL U406 ( .A(n900), .B(n885), .Y(n827) );
  XNOR2XL U407 ( .A(n900), .B(n852), .Y(n857) );
  XNOR2XL U408 ( .A(B[3]), .B(n860), .Y(n816) );
  XNOR2XL U409 ( .A(B[3]), .B(n881), .Y(n851) );
  XNOR2X1 U410 ( .A(n1052), .B(n889), .Y(n830) );
  XNOR2XL U411 ( .A(n894), .B(n852), .Y(n895) );
  XNOR2XL U412 ( .A(n900), .B(n898), .Y(n933) );
  BUFX3 U413 ( .A(n1011), .Y(n932) );
  XNOR2XL U414 ( .A(n900), .B(n893), .Y(n909) );
  XNOR2XL U415 ( .A(n6), .B(n898), .Y(n911) );
  XNOR2XL U416 ( .A(n6), .B(A[8]), .Y(n912) );
  XNOR2XL U417 ( .A(n900), .B(n899), .Y(n910) );
  BUFX3 U418 ( .A(n543), .Y(n968) );
  OAI22XL U419 ( .A0(n951), .A1(n882), .B0(n861), .B1(n1006), .Y(n915) );
  NAND2BXL U420 ( .AN(n402), .B(B[16]), .Y(n862) );
  XNOR2XL U421 ( .A(n894), .B(n893), .Y(n946) );
  XNOR2XL U422 ( .A(n894), .B(n899), .Y(n948) );
  OAI22XL U423 ( .A0(n951), .A1(n353), .B0(n950), .B1(n1006), .Y(n955) );
  NOR2BXL U424 ( .AN(n402), .B(n1054), .Y(n956) );
  OAI22XL U425 ( .A0(n832), .A1(n337), .B0(n974), .B1(n975), .Y(n954) );
  INVXL U426 ( .A(B[0]), .Y(n330) );
  XNOR2XL U427 ( .A(n612), .B(n905), .Y(n423) );
  BUFX3 U428 ( .A(n825), .Y(n951) );
  OAI22XL U429 ( .A0(n8), .A1(n420), .B0(n947), .B1(n419), .Y(n445) );
  OAI22XL U430 ( .A0(n928), .A1(n436), .B0(n926), .B1(n418), .Y(n446) );
  XNOR2XL U431 ( .A(n894), .B(n402), .Y(n420) );
  OAI22XL U432 ( .A0(n928), .A1(n418), .B0(n926), .B1(n408), .Y(n417) );
  ADDFX2 U433 ( .A(n81), .B(n80), .CI(n79), .CO(n95), .S(n530) );
  OAI22XL U434 ( .A0(n932), .A1(n72), .B0(n930), .B1(n86), .Y(n81) );
  INVXL U435 ( .A(n1056), .Y(n1061) );
  NOR2XL U436 ( .A(n519), .B(n1050), .Y(n1062) );
  NAND2XL U437 ( .A(n494), .B(n493), .Y(n1108) );
  OAI22XL U438 ( .A0(n913), .A1(n550), .B0(n543), .B1(n542), .Y(n567) );
  OAI22XL U439 ( .A0(n951), .A1(n402), .B0(n423), .B1(n1006), .Y(n1223) );
  NAND2XL U440 ( .A(n424), .B(n951), .Y(n1222) );
  NAND2BXL U441 ( .AN(n402), .B(n612), .Y(n424) );
  NAND2XL U442 ( .A(n1223), .B(n1222), .Y(n1224) );
  INVXL U443 ( .A(n1146), .Y(n1165) );
  NOR2XL U444 ( .A(n116), .B(n115), .Y(n296) );
  NOR2XL U445 ( .A(n120), .B(n119), .Y(n275) );
  AOI21XL U446 ( .A0(n270), .A1(n243), .B0(n242), .Y(n244) );
  OAI21X1 U447 ( .A0(n292), .A1(n297), .B0(n293), .Y(n285) );
  NOR2X1 U448 ( .A(n296), .B(n292), .Y(n284) );
  NOR2X1 U449 ( .A(n304), .B(n309), .Y(n112) );
  AOI21XL U450 ( .A0(n1252), .A1(n97), .B0(n96), .Y(n1141) );
  NOR2XL U451 ( .A(n1247), .B(n1249), .Y(n97) );
  XNOR2XL U452 ( .A(n612), .B(A[8]), .Y(n472) );
  XNOR2XL U453 ( .A(n612), .B(n893), .Y(n346) );
  XNOR2XL U454 ( .A(n612), .B(n852), .Y(n354) );
  NAND2BXL U455 ( .AN(n402), .B(n900), .Y(n403) );
  XNOR2XL U456 ( .A(n612), .B(n884), .Y(n473) );
  OAI21XL U457 ( .A0(n313), .A1(n309), .B0(n310), .Y(n308) );
  INVXL U458 ( .A(n304), .Y(n306) );
  INVXL U459 ( .A(n297), .Y(n60) );
  NAND2XL U460 ( .A(n118), .B(n117), .Y(n293) );
  INVXL U461 ( .A(n296), .Y(n298) );
  AOI21XL U462 ( .A0(n270), .A1(n272), .B0(n261), .Y(n262) );
  INVXL U463 ( .A(n220), .Y(n222) );
  INVXL U464 ( .A(n223), .Y(n212) );
  NAND2XL U465 ( .A(n220), .B(n224), .Y(n214) );
  INVXL U466 ( .A(n215), .Y(n217) );
  INVXL U467 ( .A(n205), .Y(n207) );
  NAND2XL U468 ( .A(n1255), .B(n1254), .Y(n199) );
  INVXL U469 ( .A(n199), .Y(n159) );
  INVXL U470 ( .A(n1240), .Y(n149) );
  NAND2XL U471 ( .A(n200), .B(n162), .Y(n151) );
  INVXL U472 ( .A(n1239), .Y(n162) );
  NAND2XL U473 ( .A(n1257), .B(n1256), .Y(n206) );
  NAND2XL U474 ( .A(n236), .B(n134), .Y(n136) );
  NAND2XL U475 ( .A(n327), .B(n1119), .Y(n1122) );
  NAND2BX1 U476 ( .AN(n1308), .B(n63), .Y(n327) );
  INVX1 U477 ( .A(n1307), .Y(n63) );
  XNOR2XL U478 ( .A(n1189), .B(n1188), .Y(PRODUCT[11]) );
  NAND2XL U479 ( .A(n1187), .B(n1248), .Y(n1188) );
  XNOR2XL U480 ( .A(n1049), .B(n794), .Y(n171) );
  XNOR2XL U481 ( .A(n1027), .B(n1051), .Y(n1045) );
  XNOR2XL U482 ( .A(n1049), .B(n1025), .Y(n1026) );
  XNOR2XL U483 ( .A(n1012), .B(A[24]), .Y(n1028) );
  XNOR2XL U484 ( .A(n1052), .B(A[22]), .Y(n1024) );
  XNOR2XL U485 ( .A(n1049), .B(n860), .Y(n76) );
  XNOR2XL U486 ( .A(n1049), .B(n885), .Y(n520) );
  XNOR2XL U487 ( .A(n612), .B(A[24]), .Y(n615) );
  XNOR2XL U488 ( .A(n612), .B(n1048), .Y(n675) );
  XNOR2XL U489 ( .A(n612), .B(A[22]), .Y(n704) );
  XNOR2XL U490 ( .A(n612), .B(n1025), .Y(n733) );
  XNOR2XL U491 ( .A(n612), .B(n1007), .Y(n764) );
  XNOR2XL U492 ( .A(n612), .B(n763), .Y(n795) );
  XNOR2XL U493 ( .A(n612), .B(n794), .Y(n824) );
  XNOR2XL U494 ( .A(n612), .B(n823), .Y(n861) );
  XNOR2XL U495 ( .A(n612), .B(n850), .Y(n950) );
  XNOR2XL U496 ( .A(n612), .B(n885), .Y(n353) );
  XNOR2XL U497 ( .A(n1027), .B(n905), .Y(n337) );
  XNOR2XL U498 ( .A(n1027), .B(n402), .Y(n338) );
  XNOR2XL U499 ( .A(n9), .B(n883), .Y(n347) );
  OAI22XL U500 ( .A0(n951), .A1(n469), .B0(n389), .B1(n1006), .Y(n1076) );
  OAI22XL U501 ( .A0(n913), .A1(n459), .B0(n968), .B1(n390), .Y(n1075) );
  OAI22XL U502 ( .A0(n928), .A1(n393), .B0(n926), .B1(n371), .Y(n394) );
  OAI22XL U503 ( .A0(n932), .A1(n370), .B0(n930), .B1(n369), .Y(n395) );
  OAI22XL U504 ( .A0(n8), .A1(n372), .B0(n947), .B1(n364), .Y(n375) );
  OAI22XL U505 ( .A0(n828), .A1(n368), .B0(n934), .B1(n362), .Y(n377) );
  OAI22XL U506 ( .A0(n928), .A1(n371), .B0(n926), .B1(n363), .Y(n376) );
  XNOR2XL U507 ( .A(n612), .B(n883), .Y(n428) );
  OAI22XL U508 ( .A0(n8), .A1(n407), .B0(n947), .B1(n464), .Y(n479) );
  XNOR2XL U509 ( .A(n886), .B(n889), .Y(n408) );
  XNOR2XL U510 ( .A(n886), .B(n888), .Y(n418) );
  NAND2BXL U511 ( .AN(n402), .B(n894), .Y(n411) );
  OAI22XL U512 ( .A0(n8), .A1(n419), .B0(n947), .B1(n407), .Y(n412) );
  XOR2X1 U513 ( .A(n300), .B(n299), .Y(PRODUCT[21]) );
  NAND2XL U514 ( .A(n298), .B(n297), .Y(n299) );
  XOR2X2 U515 ( .A(n1180), .B(n235), .Y(PRODUCT[29]) );
  INVXL U516 ( .A(n232), .Y(n234) );
  OAI21X2 U517 ( .A0(n1180), .A1(n232), .B0(n233), .Y(n231) );
  XNOR2X1 U518 ( .A(n324), .B(n323), .Y(PRODUCT[17]) );
  XOR2XL U519 ( .A(n1123), .B(n1120), .Y(PRODUCT[14]) );
  NAND2XL U520 ( .A(n1119), .B(n1242), .Y(n1120) );
  INVXL U521 ( .A(n185), .Y(n168) );
  OAI22XL U522 ( .A0(n1011), .A1(n86), .B0(n930), .B1(n176), .Y(n169) );
  INVXL U523 ( .A(n1045), .Y(n1046) );
  XNOR2XL U524 ( .A(n1052), .B(n1048), .Y(n1040) );
  XNOR2XL U525 ( .A(n1052), .B(A[24]), .Y(n1055) );
  OAI2BB1XL U526 ( .A0N(n335), .A1N(n1011), .B0(n1010), .Y(n1021) );
  NOR2XL U527 ( .A(n519), .B(n1008), .Y(n1023) );
  INVXL U528 ( .A(n1009), .Y(n1010) );
  OAI22XL U529 ( .A0(n8), .A1(n392), .B0(n947), .B1(n372), .Y(n1072) );
  OAI22XL U530 ( .A0(n928), .A1(n467), .B0(n926), .B1(n393), .Y(n1091) );
  OAI22XL U531 ( .A0(n8), .A1(n464), .B0(n947), .B1(n463), .Y(n482) );
  OAI22XL U532 ( .A0(n928), .A1(n462), .B0(n926), .B1(n468), .Y(n483) );
  OAI22XL U533 ( .A0(n8), .A1(n463), .B0(n947), .B1(n461), .Y(n1078) );
  OAI22XL U534 ( .A0(n913), .A1(n460), .B0(n968), .B1(n459), .Y(n1079) );
  OAI22XL U535 ( .A0(n828), .A1(n474), .B0(n934), .B1(n458), .Y(n1080) );
  OAI22XL U536 ( .A0(n928), .A1(n468), .B0(n926), .B1(n467), .Y(n1096) );
  OAI22XL U537 ( .A0(n913), .A1(n73), .B0(n968), .B1(n87), .Y(n84) );
  OAI22XL U538 ( .A0(n832), .A1(n75), .B0(n974), .B1(n88), .Y(n82) );
  OAI22XL U539 ( .A0(n8), .A1(n586), .B0(n947), .B1(n547), .Y(n573) );
  OAI22XL U540 ( .A0(n828), .A1(n568), .B0(n934), .B1(n549), .Y(n571) );
  OAI22XL U541 ( .A0(n932), .A1(n588), .B0(n930), .B1(n552), .Y(n574) );
  OAI22XL U542 ( .A0(n913), .A1(n587), .B0(n968), .B1(n550), .Y(n576) );
  OAI22XL U543 ( .A0(n832), .A1(n585), .B0(n974), .B1(n551), .Y(n575) );
  OAI22XL U544 ( .A0(n913), .A1(n672), .B0(n968), .B1(n625), .Y(n656) );
  OAI22XL U545 ( .A0(n8), .A1(n650), .B0(n947), .B1(n618), .Y(n651) );
  OAI22XL U546 ( .A0(n786), .A1(n649), .B0(n926), .B1(n608), .Y(n652) );
  OAI22XL U547 ( .A0(n932), .A1(n648), .B0(n930), .B1(n607), .Y(n653) );
  OAI22XL U548 ( .A0(n8), .A1(n668), .B0(n947), .B1(n650), .Y(n669) );
  OAI22XL U549 ( .A0(n1011), .A1(n666), .B0(n930), .B1(n648), .Y(n671) );
  OAI22XL U550 ( .A0(n928), .A1(n667), .B0(n926), .B1(n649), .Y(n670) );
  OAI22XL U551 ( .A0(n8), .A1(n697), .B0(n947), .B1(n668), .Y(n698) );
  OAI22XL U552 ( .A0(n932), .A1(n695), .B0(n930), .B1(n666), .Y(n700) );
  OAI22XL U553 ( .A0(n928), .A1(n696), .B0(n926), .B1(n667), .Y(n699) );
  OAI22XL U554 ( .A0(n8), .A1(n726), .B0(n947), .B1(n697), .Y(n727) );
  OAI22XL U555 ( .A0(n932), .A1(n724), .B0(n930), .B1(n695), .Y(n729) );
  OAI22XL U556 ( .A0(n928), .A1(n725), .B0(n926), .B1(n696), .Y(n728) );
  OAI22XL U557 ( .A0(n8), .A1(n756), .B0(n947), .B1(n726), .Y(n757) );
  OAI22XL U558 ( .A0(n932), .A1(n753), .B0(n930), .B1(n724), .Y(n759) );
  OAI22XL U559 ( .A0(n928), .A1(n754), .B0(n926), .B1(n725), .Y(n758) );
  OAI22XL U560 ( .A0(n8), .A1(n787), .B0(n947), .B1(n756), .Y(n788) );
  OAI22XL U561 ( .A0(n786), .A1(n785), .B0(n926), .B1(n754), .Y(n789) );
  OAI22XL U562 ( .A0(n932), .A1(n784), .B0(n930), .B1(n753), .Y(n790) );
  OAI22XL U563 ( .A0(n8), .A1(n854), .B0(n947), .B1(n787), .Y(n817) );
  OAI22XL U564 ( .A0(n786), .A1(n816), .B0(n926), .B1(n785), .Y(n818) );
  OAI22XL U565 ( .A0(n932), .A1(n815), .B0(n930), .B1(n784), .Y(n819) );
  OAI22XL U566 ( .A0(n8), .A1(n895), .B0(n947), .B1(n855), .Y(n890) );
  OAI22XL U567 ( .A0(n932), .A1(n897), .B0(n930), .B1(n849), .Y(n892) );
  OAI22XL U568 ( .A0(n928), .A1(n887), .B0(n926), .B1(n851), .Y(n891) );
  OAI22XL U569 ( .A0(n970), .A1(n967), .B0(n968), .B1(n912), .Y(n939) );
  OAI22XL U570 ( .A0(n832), .A1(n973), .B0(n974), .B1(n908), .Y(n937) );
  OAI22XL U571 ( .A0(n928), .A1(n925), .B0(n926), .B1(n887), .Y(n938) );
  OAI22XL U572 ( .A0(n904), .A1(n971), .B0(n1054), .B1(n903), .Y(n965) );
  OAI22XL U573 ( .A0(n828), .A1(n935), .B0(n934), .B1(n933), .Y(n943) );
  OAI22XL U574 ( .A0(n928), .A1(n927), .B0(n926), .B1(n925), .Y(n945) );
  OAI22XL U575 ( .A0(n970), .A1(n969), .B0(n968), .B1(n967), .Y(n981) );
  OAI22XL U576 ( .A0(n832), .A1(n975), .B0(n974), .B1(n973), .Y(n979) );
  OAI22XL U577 ( .A0(n928), .A1(n336), .B0(n926), .B1(n927), .Y(n976) );
  OAI22XL U578 ( .A0(n970), .A1(n334), .B0(n968), .B1(n969), .Y(n978) );
  OAI22XL U579 ( .A0(n932), .A1(n339), .B0(n930), .B1(n931), .Y(n977) );
  OAI22XL U580 ( .A0(n8), .A1(n364), .B0(n947), .B1(n351), .Y(n340) );
  OAI22XL U581 ( .A0(n913), .A1(n343), .B0(n968), .B1(n334), .Y(n342) );
  OAI22XL U582 ( .A0(n8), .A1(n351), .B0(n947), .B1(n948), .Y(n984) );
  OAI22XL U583 ( .A0(n828), .A1(n352), .B0(n934), .B1(n935), .Y(n983) );
  INVXL U584 ( .A(n1022), .Y(n1015) );
  NOR2XL U585 ( .A(n519), .B(n181), .Y(n1016) );
  OAI22XL U586 ( .A0(n832), .A1(n183), .B0(n974), .B1(n1013), .Y(n1020) );
  ADDFX2 U587 ( .A(n388), .B(n386), .CI(n387), .CO(n378), .S(n1069) );
  OAI22XL U588 ( .A0(n951), .A1(n423), .B0(n428), .B1(n1006), .Y(n426) );
  NOR2BXL U589 ( .AN(n402), .B(n926), .Y(n425) );
  OAI22XL U590 ( .A0(n928), .A1(n431), .B0(n926), .B1(n430), .Y(n432) );
  NAND2BXL U591 ( .AN(n402), .B(n886), .Y(n430) );
  OAI22XL U592 ( .A0(n951), .A1(n435), .B0(n434), .B1(n1006), .Y(n448) );
  NOR2BXL U593 ( .AN(n402), .B(n947), .Y(n449) );
  OAI22XL U594 ( .A0(n928), .A1(n437), .B0(n926), .B1(n436), .Y(n447) );
  ADDFX2 U595 ( .A(n490), .B(n489), .CI(n488), .CO(n491), .S(n455) );
  NAND2XL U596 ( .A(n1156), .B(n1238), .Y(n157) );
  NAND2XL U597 ( .A(n1159), .B(n1236), .Y(n1160) );
  XNOR2XL U598 ( .A(n1173), .B(n1232), .Y(PRODUCT[39]) );
  NAND2XL U599 ( .A(n1174), .B(n1170), .Y(n1172) );
  XNOR2XL U600 ( .A(n1183), .B(n1182), .Y(PRODUCT[38]) );
  NAND2XL U601 ( .A(n1181), .B(n1234), .Y(n1182) );
  NOR2XL U602 ( .A(n519), .B(n89), .Y(n166) );
  OAI22XL U603 ( .A0(n832), .A1(n88), .B0(n974), .B1(n175), .Y(n167) );
  XNOR2XL U604 ( .A(n1049), .B(n823), .Y(n89) );
  ADDFX2 U605 ( .A(n179), .B(n178), .CI(n177), .CO(n500), .S(n93) );
  OAI22XL U606 ( .A0(n913), .A1(n515), .B0(n968), .B1(n73), .Y(n511) );
  INVXL U607 ( .A(n91), .Y(n510) );
  OAI22XL U608 ( .A0(n932), .A1(n516), .B0(n930), .B1(n72), .Y(n507) );
  NOR2XL U609 ( .A(n519), .B(n69), .Y(n509) );
  OAI22XL U610 ( .A0(n932), .A1(n523), .B0(n930), .B1(n516), .Y(n541) );
  OAI22XL U611 ( .A0(n832), .A1(n518), .B0(n974), .B1(n517), .Y(n540) );
  OAI22XL U612 ( .A0(n932), .A1(n552), .B0(n930), .B1(n523), .Y(n556) );
  OAI22XL U613 ( .A0(n828), .A1(n549), .B0(n934), .B1(n521), .Y(n558) );
  OAI2BB1XL U614 ( .A0N(n947), .A1N(n8), .B0(n506), .Y(n524) );
  INVXL U615 ( .A(n505), .Y(n506) );
  OAI22XL U616 ( .A0(n913), .A1(n542), .B0(n968), .B1(n515), .Y(n527) );
  OAI22XL U617 ( .A0(n828), .A1(n521), .B0(n934), .B1(n513), .Y(n529) );
  ADDFX2 U618 ( .A(n579), .B(n578), .CI(n577), .CO(n559), .S(n580) );
  OAI2BB1XL U619 ( .A0N(n926), .A1N(n786), .B0(n546), .Y(n598) );
  INVXL U620 ( .A(n545), .Y(n546) );
  OAI22XL U621 ( .A0(n904), .A1(n591), .B0(n1054), .B1(n570), .Y(n621) );
  OAI22XL U622 ( .A0(n828), .A1(n590), .B0(n934), .B1(n568), .Y(n623) );
  OAI22XL U623 ( .A0(n913), .A1(n625), .B0(n968), .B1(n624), .Y(n638) );
  XNOR2XL U624 ( .A(n629), .B(n628), .Y(n636) );
  OAI22XL U625 ( .A0(n8), .A1(n618), .B0(n947), .B1(n617), .Y(n635) );
  OAI22XL U626 ( .A0(n832), .A1(n632), .B0(n974), .B1(n620), .Y(n633) );
  OAI2BB1XL U627 ( .A0N(n1006), .A1N(n825), .B0(n584), .Y(n609) );
  OAI22XL U628 ( .A0(n932), .A1(n607), .B0(n930), .B1(n589), .Y(n611) );
  OAI22XL U629 ( .A0(n786), .A1(n608), .B0(n926), .B1(n583), .Y(n610) );
  OAI22XL U630 ( .A0(n8), .A1(n617), .B0(n947), .B1(n586), .Y(n596) );
  OAI22XL U631 ( .A0(n913), .A1(n624), .B0(n968), .B1(n587), .Y(n603) );
  OAI22XL U632 ( .A0(n932), .A1(n589), .B0(n930), .B1(n588), .Y(n602) );
  ADDFX2 U633 ( .A(n688), .B(n687), .CI(n686), .CO(n665), .S(n689) );
  OAI22XL U634 ( .A0(n832), .A1(n679), .B0(n974), .B1(n632), .Y(n680) );
  OAI22XL U635 ( .A0(n828), .A1(n677), .B0(n934), .B1(n630), .Y(n682) );
  OAI22XL U636 ( .A0(n913), .A1(n701), .B0(n968), .B1(n672), .Y(n685) );
  ADDFX2 U637 ( .A(n717), .B(n716), .CI(n715), .CO(n691), .S(n718) );
  OAI22XL U638 ( .A0(n913), .A1(n730), .B0(n968), .B1(n701), .Y(n714) );
  OAI22XL U639 ( .A0(n832), .A1(n708), .B0(n974), .B1(n679), .Y(n709) );
  OAI22XL U640 ( .A0(n828), .A1(n706), .B0(n934), .B1(n677), .Y(n711) );
  ADDFX2 U641 ( .A(n746), .B(n745), .CI(n744), .CO(n720), .S(n747) );
  OAI22XL U642 ( .A0(n913), .A1(n760), .B0(n968), .B1(n730), .Y(n743) );
  OAI22XL U643 ( .A0(n832), .A1(n737), .B0(n974), .B1(n708), .Y(n738) );
  OAI22XL U644 ( .A0(n828), .A1(n735), .B0(n934), .B1(n706), .Y(n740) );
  OAI22XL U645 ( .A0(n913), .A1(n791), .B0(n968), .B1(n760), .Y(n774) );
  OAI22XL U646 ( .A0(n832), .A1(n768), .B0(n974), .B1(n737), .Y(n769) );
  OAI22XL U647 ( .A0(n828), .A1(n766), .B0(n934), .B1(n735), .Y(n771) );
  OAI22XL U648 ( .A0(n913), .A1(n820), .B0(n968), .B1(n791), .Y(n805) );
  OAI22XL U649 ( .A0(n828), .A1(n797), .B0(n934), .B1(n766), .Y(n802) );
  OAI22XL U650 ( .A0(n913), .A1(n853), .B0(n968), .B1(n820), .Y(n838) );
  OAI22XL U651 ( .A0(n832), .A1(n831), .B0(n974), .B1(n799), .Y(n833) );
  OAI22XL U652 ( .A0(n828), .A1(n827), .B0(n934), .B1(n797), .Y(n835) );
  OAI22XL U653 ( .A0(n828), .A1(n909), .B0(n934), .B1(n857), .Y(n871) );
  OAI22XL U654 ( .A0(n8), .A1(n855), .B0(n947), .B1(n854), .Y(n864) );
  OAI22XL U655 ( .A0(n913), .A1(n911), .B0(n968), .B1(n853), .Y(n865) );
  OAI22XL U656 ( .A0(n832), .A1(n907), .B0(n974), .B1(n856), .Y(n863) );
  OAI22XL U657 ( .A0(n828), .A1(n857), .B0(n934), .B1(n827), .Y(n868) );
  OAI22XL U658 ( .A0(n832), .A1(n856), .B0(n974), .B1(n831), .Y(n866) );
  OAI22X1 U659 ( .A0(n904), .A1(n830), .B0(n1054), .B1(n829), .Y(n867) );
  OAI22XL U660 ( .A0(n928), .A1(n851), .B0(n926), .B1(n816), .Y(n1199) );
  OAI22XL U661 ( .A0(n932), .A1(n849), .B0(n930), .B1(n815), .Y(n1201) );
  OAI22XL U662 ( .A0(n904), .A1(n902), .B0(n1054), .B1(n830), .Y(n1200) );
  OAI22XL U663 ( .A0(n828), .A1(n933), .B0(n901), .B1(n910), .Y(n940) );
  OAI22XL U664 ( .A0(n8), .A1(n946), .B0(n947), .B1(n895), .Y(n942) );
  OAI22XL U665 ( .A0(n832), .A1(n908), .B0(n974), .B1(n907), .Y(n1193) );
  OAI22XL U666 ( .A0(n913), .A1(n912), .B0(n968), .B1(n911), .Y(n1197) );
  OAI22XL U667 ( .A0(n828), .A1(n910), .B0(n934), .B1(n909), .Y(n1198) );
  OAI22XL U668 ( .A0(n8), .A1(n948), .B0(n947), .B1(n946), .Y(n962) );
  ADDFX2 U669 ( .A(n1131), .B(n1130), .CI(n1129), .CO(n1140), .S(n989) );
  ADDFX2 U670 ( .A(n993), .B(n992), .CI(n991), .CO(n988), .S(n1002) );
  ADDFX2 U671 ( .A(n380), .B(n379), .CI(n378), .CO(n1004), .S(n383) );
  NAND2XL U672 ( .A(n426), .B(n425), .Y(n1218) );
  INVXL U673 ( .A(n1224), .Y(n1220) );
  NOR2XL U674 ( .A(n433), .B(n432), .Y(n1213) );
  NAND2XL U675 ( .A(n433), .B(n432), .Y(n1214) );
  AOI21XL U676 ( .A0(n1219), .A1(n1220), .B0(n427), .Y(n1216) );
  INVXL U677 ( .A(n1218), .Y(n427) );
  NAND2XL U678 ( .A(n442), .B(n441), .Y(n1210) );
  AOI21XL U679 ( .A0(n1211), .A1(n440), .B0(n443), .Y(n1208) );
  INVXL U680 ( .A(n1210), .Y(n443) );
  NOR2XL U681 ( .A(n451), .B(n450), .Y(n1205) );
  NAND2XL U682 ( .A(n451), .B(n450), .Y(n1206) );
  NOR2XL U683 ( .A(n1087), .B(n1086), .Y(mult_x_1_n136) );
  NOR2XL U684 ( .A(n1033), .B(n1032), .Y(mult_x_1_n129) );
  NAND2XL U685 ( .A(n1087), .B(n1086), .Y(mult_x_1_n137) );
  NOR2XL U686 ( .A(n1085), .B(n1084), .Y(mult_x_1_n319) );
  NAND2XL U687 ( .A(n1066), .B(n1065), .Y(mult_x_1_n59) );
  NAND2XL U688 ( .A(n1064), .B(n1063), .Y(n1065) );
  NOR2XL U689 ( .A(n1110), .B(n1109), .Y(mult_x_1_n120) );
  NAND2XL U690 ( .A(n1110), .B(n1109), .Y(mult_x_1_n121) );
  NAND2XL U691 ( .A(n1033), .B(n1032), .Y(mult_x_1_n130) );
  NAND2XL U692 ( .A(n1085), .B(n1084), .Y(mult_x_1_n320) );
  NOR2XL U693 ( .A(n1101), .B(n1100), .Y(mult_x_1_n325) );
  NAND2XL U694 ( .A(n1101), .B(n1100), .Y(mult_x_1_n326) );
  NOR2XL U695 ( .A(n1118), .B(n1117), .Y(mult_x_1_n328) );
  NAND2XL U696 ( .A(n1118), .B(n1117), .Y(mult_x_1_n329) );
  NAND2XL U697 ( .A(n484), .B(n1108), .Y(mult_x_1_n89) );
  INVXL U698 ( .A(n1108), .Y(n495) );
  ADDFX2 U699 ( .A(n535), .B(n534), .CI(n533), .CO(mult_x_1_n459), .S(
        mult_x_1_n460) );
  ADDFX2 U700 ( .A(n921), .B(n920), .CI(n919), .CO(mult_x_1_n667), .S(
        mult_x_1_n668) );
  NOR2BXL U701 ( .AN(n402), .B(n1006), .Y(n1329) );
  XNOR2XL U702 ( .A(n1221), .B(n1220), .Y(n1327) );
  NAND2XL U703 ( .A(n1219), .B(n1218), .Y(n1221) );
  XOR2XL U704 ( .A(n1217), .B(n1216), .Y(n1326) );
  NAND2XL U705 ( .A(n1215), .B(n1214), .Y(n1217) );
  INVXL U706 ( .A(n1213), .Y(n1215) );
  XNOR2XL U707 ( .A(n1212), .B(n1211), .Y(n1325) );
  NAND2XL U708 ( .A(n440), .B(n1210), .Y(n1212) );
  XOR2XL U709 ( .A(n1209), .B(n1208), .Y(n1324) );
  NAND2XL U710 ( .A(n1207), .B(n1206), .Y(n1209) );
  INVXL U711 ( .A(n1205), .Y(n1207) );
  XOR2XL U712 ( .A(n1166), .B(n1165), .Y(n1323) );
  NAND2XL U713 ( .A(n1164), .B(n1163), .Y(n1166) );
  INVXL U714 ( .A(n1162), .Y(n1164) );
  NAND2XL U715 ( .A(n1149), .B(n1148), .Y(n1150) );
  INVXL U716 ( .A(n1147), .Y(n1149) );
  INVX1 U717 ( .A(n240), .Y(n270) );
  CMPR22X1 U718 ( .A(n466), .B(n465), .CO(n481), .S(n490) );
  OAI22X1 U719 ( .A0(n828), .A1(n404), .B0(n934), .B1(n403), .Y(n465) );
  CMPR22X1 U720 ( .A(n674), .B(n673), .CO(n654), .S(n684) );
  CMPR22X1 U721 ( .A(n732), .B(n731), .CO(n712), .S(n742) );
  CMPR22X1 U722 ( .A(n793), .B(n792), .CO(n772), .S(n804) );
  CMPR22X1 U723 ( .A(n859), .B(n858), .CO(n836), .S(n870) );
  OAI22X1 U724 ( .A0(n928), .A1(n583), .B0(n926), .B1(n545), .Y(n599) );
  BUFX3 U725 ( .A(n786), .Y(n928) );
  CMPR22X1 U726 ( .A(n358), .B(n357), .CO(n982), .S(n367) );
  OAI22X1 U727 ( .A0(n951), .A1(n950), .B0(n949), .B1(n1006), .Y(n964) );
  OAI22X1 U728 ( .A0(n8), .A1(n547), .B0(n947), .B1(n505), .Y(n525) );
  XNOR2X1 U729 ( .A(n894), .B(n1051), .Y(n505) );
  CMPR22X1 U730 ( .A(n627), .B(n626), .CO(n637), .S(n655) );
  CMPR22X1 U731 ( .A(n422), .B(n421), .CO(n416), .S(n444) );
  OAI22X1 U732 ( .A0(n904), .A1(n631), .B0(n1054), .B1(n591), .Y(n628) );
  CMPR22X1 U733 ( .A(n964), .B(n963), .CO(n1131), .S(n961) );
  XOR2X1 U734 ( .A(n59), .B(n295), .Y(PRODUCT[22]) );
  XNOR2X1 U735 ( .A(n274), .B(n273), .Y(PRODUCT[25]) );
  CLKINVX3 U736 ( .A(n431), .Y(n886) );
  AOI2BB1X2 U737 ( .A0N(n62), .A1N(n1242), .B0(n101), .Y(n1121) );
  OAI21X4 U738 ( .A0(n114), .A1(n301), .B0(n113), .Y(n239) );
  XOR2X4 U739 ( .A(B[11]), .B(n61), .Y(n974) );
  AOI21X1 U740 ( .A0(n324), .A1(n303), .B0(n302), .Y(n313) );
  OAI21X2 U741 ( .A0(n316), .A1(n321), .B0(n317), .Y(n302) );
  NAND2X1 U742 ( .A(n104), .B(n1303), .Y(n321) );
  NAND2BX2 U743 ( .AN(n102), .B(n64), .Y(n324) );
  NAND2X1 U744 ( .A(n325), .B(n103), .Y(n64) );
  OAI21XL U745 ( .A0(n1180), .A1(n204), .B0(n203), .Y(n209) );
  XNOR2X1 U746 ( .A(n209), .B(n208), .Y(PRODUCT[33]) );
  XNOR2X1 U747 ( .A(n202), .B(n201), .Y(PRODUCT[34]) );
  XNOR2X1 U748 ( .A(n250), .B(n249), .Y(PRODUCT[28]) );
  OAI21XL U749 ( .A0(n245), .A1(n300), .B0(n244), .Y(n250) );
  XNOR2X1 U750 ( .A(n259), .B(n258), .Y(PRODUCT[27]) );
  XNOR2X1 U751 ( .A(n164), .B(n163), .Y(PRODUCT[35]) );
  AOI21X2 U752 ( .A0(n124), .A1(n285), .B0(n123), .Y(n240) );
  NOR2X1 U753 ( .A(n237), .B(n246), .Y(n134) );
  XNOR2XL U754 ( .A(n886), .B(n402), .Y(n429) );
  XNOR2XL U755 ( .A(n1049), .B(n898), .Y(n614) );
  XNOR2XL U756 ( .A(n1049), .B(n896), .Y(n734) );
  XNOR2XL U757 ( .A(n1049), .B(n883), .Y(n826) );
  XNOR2XL U758 ( .A(n1012), .B(n1007), .Y(n88) );
  XNOR2XL U759 ( .A(n9), .B(n823), .Y(n588) );
  XNOR2XL U760 ( .A(n9), .B(n881), .Y(n607) );
  XOR2X1 U761 ( .A(B[10]), .B(B[11]), .Y(n65) );
  XNOR2X1 U762 ( .A(B[10]), .B(B[9]), .Y(n335) );
  XOR2X1 U763 ( .A(B[12]), .B(B[13]), .Y(n66) );
  CLKINVX3 U764 ( .A(n67), .Y(n1012) );
  XNOR2X1 U765 ( .A(n1012), .B(n794), .Y(n517) );
  XNOR2X1 U766 ( .A(n1012), .B(n763), .Y(n75) );
  OAI22X1 U767 ( .A0(n832), .A1(n517), .B0(n974), .B1(n75), .Y(n512) );
  XOR2X1 U768 ( .A(B[6]), .B(B[7]), .Y(n68) );
  BUFX4 U769 ( .A(B[7]), .Y(n900) );
  OAI22X1 U770 ( .A0(n828), .A1(n513), .B0(n934), .B1(n77), .Y(n91) );
  XNOR2X1 U771 ( .A(n1049), .B(n881), .Y(n69) );
  NAND2X4 U772 ( .A(n70), .B(n71), .Y(n904) );
  INVX8 U773 ( .A(n953), .Y(n1052) );
  XNOR2X1 U774 ( .A(n1052), .B(n860), .Y(n514) );
  BUFX1 U775 ( .A(A[17]), .Y(n823) );
  XNOR2X1 U776 ( .A(n1052), .B(n823), .Y(n74) );
  OAI2BB1X1 U777 ( .A0N(n934), .A1N(n828), .B0(n78), .Y(n90) );
  CMPR32X1 U778 ( .A(n84), .B(n83), .C(n82), .CO(n179), .S(n532) );
  OAI22X1 U779 ( .A0(n913), .A1(n87), .B0(n968), .B1(n172), .Y(n185) );
  XNOR2XL U780 ( .A(n1012), .B(n1025), .Y(n175) );
  ADDFHX1 U781 ( .A(n1289), .B(n1287), .CI(n1285), .CO(n119), .S(n118) );
  ADDFHX1 U782 ( .A(n1286), .B(n1284), .CI(n1282), .CO(n121), .S(n120) );
  NOR2XL U783 ( .A(n126), .B(n125), .Y(n260) );
  CMPR32X1 U784 ( .A(n1280), .B(n1278), .C(n1276), .CO(n127), .S(n126) );
  NOR2XL U785 ( .A(n260), .B(n264), .Y(n236) );
  NOR2X1 U786 ( .A(n132), .B(n131), .Y(n246) );
  NOR2X1 U787 ( .A(n238), .B(n136), .Y(n138) );
  NAND2X1 U788 ( .A(n112), .B(n303), .Y(n114) );
  NOR2XL U789 ( .A(n1304), .B(n1306), .Y(n1124) );
  NOR2XL U790 ( .A(n1122), .B(n1124), .Y(n103) );
  OAI21XL U791 ( .A0(n1247), .A1(n1250), .B0(n1248), .Y(n96) );
  INVX1 U792 ( .A(n1245), .Y(n1190) );
  NAND2XL U793 ( .A(n1143), .B(n1190), .Y(n100) );
  INVXL U794 ( .A(n1246), .Y(n1142) );
  INVXL U795 ( .A(n1244), .Y(n98) );
  AOI21XL U796 ( .A0(n1143), .A1(n1142), .B0(n98), .Y(n99) );
  OAI21XL U797 ( .A0(n1141), .A1(n100), .B0(n99), .Y(n325) );
  NAND2XL U798 ( .A(n1307), .B(n1308), .Y(n326) );
  INVXL U799 ( .A(n326), .Y(n101) );
  NAND2XL U800 ( .A(n1304), .B(n1306), .Y(n1125) );
  OAI21XL U801 ( .A0(n1121), .A1(n1124), .B0(n1125), .Y(n102) );
  NAND2XL U802 ( .A(n110), .B(n109), .Y(n305) );
  AOI21X2 U803 ( .A0(n112), .A1(n302), .B0(n111), .Y(n113) );
  NAND2XL U804 ( .A(n120), .B(n119), .Y(n288) );
  NAND2XL U805 ( .A(n122), .B(n121), .Y(n280) );
  OAI21XL U806 ( .A0(n279), .A1(n288), .B0(n280), .Y(n123) );
  NAND2XL U807 ( .A(n128), .B(n127), .Y(n265) );
  OAI21XL U808 ( .A0(n264), .A1(n271), .B0(n265), .Y(n241) );
  NAND2X1 U809 ( .A(n130), .B(n129), .Y(n256) );
  NAND2XL U810 ( .A(n132), .B(n131), .Y(n247) );
  OAI21XL U811 ( .A0(n246), .A1(n256), .B0(n247), .Y(n133) );
  OAI21X1 U812 ( .A0(n240), .A1(n136), .B0(n135), .Y(n137) );
  AOI21X2 U813 ( .A0(n138), .A1(n239), .B0(n137), .Y(n139) );
  BUFX8 U814 ( .A(n139), .Y(n1180) );
  ADDFHX1 U815 ( .A(n1271), .B(n1269), .CI(n1267), .CO(n141), .S(n132) );
  CMPR32X1 U816 ( .A(n1268), .B(n1265), .C(n1266), .CO(n143), .S(n140) );
  NOR2XL U817 ( .A(n232), .B(n227), .Y(n220) );
  CMPR32X1 U818 ( .A(n1263), .B(n1262), .C(n1264), .CO(n144), .S(n142) );
  NOR2XL U819 ( .A(n210), .B(n215), .Y(n148) );
  OR2X2 U820 ( .A(n1255), .B(n1254), .Y(n200) );
  OR2X2 U821 ( .A(n151), .B(n205), .Y(n154) );
  NAND2XL U822 ( .A(n143), .B(n142), .Y(n228) );
  NAND2XL U823 ( .A(n145), .B(n144), .Y(n223) );
  NAND2XL U824 ( .A(n146), .B(n1258), .Y(n216) );
  OAI21XL U825 ( .A0(n215), .A1(n223), .B0(n216), .Y(n147) );
  AOI21X1 U826 ( .A0(n211), .A1(n148), .B0(n147), .Y(n203) );
  OAI21XL U827 ( .A0(n151), .A1(n206), .B0(n150), .Y(n152) );
  OAI21XL U828 ( .A0(n1180), .A1(n156), .B0(n155), .Y(n158) );
  NAND2XL U829 ( .A(n195), .B(n200), .Y(n161) );
  OAI21XL U830 ( .A0(n203), .A1(n205), .B0(n206), .Y(n196) );
  AOI21XL U831 ( .A0(n196), .A1(n200), .B0(n159), .Y(n160) );
  CMPR32X1 U832 ( .A(n167), .B(n166), .C(n165), .CO(n502), .S(n177) );
  CMPR32X1 U833 ( .A(n170), .B(n169), .C(n168), .CO(n192), .S(n178) );
  NOR2XL U834 ( .A(n519), .B(n171), .Y(n186) );
  XNOR2X1 U835 ( .A(n1052), .B(n1007), .Y(n180) );
  XNOR2XL U836 ( .A(n1012), .B(A[22]), .Y(n183) );
  OAI22XL U837 ( .A0(n832), .A1(n175), .B0(n974), .B1(n183), .Y(n188) );
  XNOR2X1 U838 ( .A(n1052), .B(n1025), .Y(n1014) );
  XNOR2X1 U839 ( .A(n1049), .B(n763), .Y(n181) );
  OAI22X1 U840 ( .A0(n1011), .A1(n182), .B0(n930), .B1(n1009), .Y(n1022) );
  CMPR32X1 U841 ( .A(n186), .B(n185), .C(n184), .CO(n1019), .S(n191) );
  CMPR32X1 U842 ( .A(n189), .B(n188), .C(n187), .CO(n1018), .S(n190) );
  CMPR32X1 U843 ( .A(n192), .B(n191), .C(n190), .CO(n1034), .S(n501) );
  NOR2XL U844 ( .A(n194), .B(n193), .Y(mult_x_1_n151) );
  NAND2XL U845 ( .A(n194), .B(n193), .Y(mult_x_1_n152) );
  INVXL U846 ( .A(n195), .Y(n198) );
  INVXL U847 ( .A(n196), .Y(n197) );
  OAI21XL U848 ( .A0(n1180), .A1(n198), .B0(n197), .Y(n202) );
  AOI21XL U849 ( .A0(n211), .A1(n224), .B0(n212), .Y(n213) );
  OAI21X4 U850 ( .A0(n1180), .A1(n214), .B0(n213), .Y(n219) );
  NAND2X1 U851 ( .A(n217), .B(n216), .Y(n218) );
  XNOR2X2 U852 ( .A(n219), .B(n218), .Y(PRODUCT[32]) );
  INVXL U853 ( .A(n211), .Y(n221) );
  OAI21X4 U854 ( .A0(n1180), .A1(n222), .B0(n221), .Y(n226) );
  NAND2X1 U855 ( .A(n224), .B(n223), .Y(n225) );
  XNOR2X4 U856 ( .A(n226), .B(n225), .Y(PRODUCT[31]) );
  NAND2X1 U857 ( .A(n229), .B(n228), .Y(n230) );
  INVXL U858 ( .A(n236), .Y(n251) );
  INVXL U859 ( .A(n237), .Y(n257) );
  NOR2XL U860 ( .A(n251), .B(n237), .Y(n243) );
  NAND2XL U861 ( .A(n243), .B(n269), .Y(n245) );
  INVXL U862 ( .A(n241), .Y(n252) );
  OAI21XL U863 ( .A0(n252), .A1(n237), .B0(n256), .Y(n242) );
  NAND2XL U864 ( .A(n248), .B(n247), .Y(n249) );
  INVXL U865 ( .A(n251), .Y(n253) );
  NAND2XL U866 ( .A(n269), .B(n253), .Y(n255) );
  AOI21XL U867 ( .A0(n270), .A1(n253), .B0(n241), .Y(n254) );
  OAI21XL U868 ( .A0(n300), .A1(n255), .B0(n254), .Y(n259) );
  INVXL U869 ( .A(n260), .Y(n272) );
  INVXL U870 ( .A(n271), .Y(n261) );
  OAI21XL U871 ( .A0(n300), .A1(n263), .B0(n262), .Y(n268) );
  INVXL U872 ( .A(n264), .Y(n266) );
  XNOR2X1 U873 ( .A(n268), .B(n267), .Y(PRODUCT[26]) );
  OAI21XL U874 ( .A0(n300), .A1(n238), .B0(n240), .Y(n274) );
  INVXL U875 ( .A(n275), .Y(n289) );
  NAND2XL U876 ( .A(n284), .B(n289), .Y(n278) );
  INVXL U877 ( .A(n288), .Y(n276) );
  AOI21XL U878 ( .A0(n285), .A1(n289), .B0(n276), .Y(n277) );
  OAI21XL U879 ( .A0(n300), .A1(n278), .B0(n277), .Y(n283) );
  INVXL U880 ( .A(n279), .Y(n281) );
  NAND2X1 U881 ( .A(n281), .B(n280), .Y(n282) );
  INVXL U882 ( .A(n284), .Y(n287) );
  INVXL U883 ( .A(n285), .Y(n286) );
  OAI21XL U884 ( .A0(n300), .A1(n287), .B0(n286), .Y(n291) );
  INVXL U885 ( .A(n292), .Y(n294) );
  NAND2XL U886 ( .A(n306), .B(n305), .Y(n307) );
  NAND2XL U887 ( .A(n311), .B(n310), .Y(n312) );
  INVXL U888 ( .A(n321), .Y(n315) );
  AOI21XL U889 ( .A0(n324), .A1(n322), .B0(n315), .Y(n320) );
  INVXL U890 ( .A(n316), .Y(n318) );
  NAND2XL U891 ( .A(n318), .B(n317), .Y(n319) );
  NAND2XL U892 ( .A(n322), .B(n321), .Y(n323) );
  INVXL U893 ( .A(n325), .Y(n1123) );
  OAI21XL U894 ( .A0(n1123), .A1(n1241), .B0(n1242), .Y(n329) );
  BUFX3 U895 ( .A(n330), .Y(n1006) );
  INVX1 U896 ( .A(B[13]), .Y(n356) );
  CLKINVX3 U897 ( .A(n356), .Y(n1027) );
  BUFX1 U898 ( .A(A[2]), .Y(n883) );
  XNOR2X1 U899 ( .A(n1027), .B(n883), .Y(n975) );
  INVX1 U900 ( .A(B[3]), .Y(n431) );
  XNOR2XL U901 ( .A(n886), .B(n893), .Y(n336) );
  OAI22XL U902 ( .A0(n928), .A1(n363), .B0(n926), .B1(n336), .Y(n341) );
  XOR2X1 U903 ( .A(B[4]), .B(B[5]), .Y(n332) );
  CLKINVX3 U904 ( .A(B[5]), .Y(n504) );
  CLKINVX3 U905 ( .A(n504), .Y(n894) );
  BUFX1 U906 ( .A(A[3]), .Y(n888) );
  BUFX3 U907 ( .A(n335), .Y(n930) );
  OAI22X1 U908 ( .A0(n828), .A1(n362), .B0(n934), .B1(n352), .Y(n350) );
  OAI22X1 U909 ( .A0(n832), .A1(n338), .B0(n974), .B1(n337), .Y(n349) );
  OAI22XL U910 ( .A0(n932), .A1(n347), .B0(n930), .B1(n339), .Y(n348) );
  CMPR32X1 U911 ( .A(n342), .B(n341), .C(n340), .CO(n958), .S(n379) );
  OAI22XL U912 ( .A0(n1011), .A1(n345), .B0(n335), .B1(n344), .Y(n373) );
  OAI22XL U913 ( .A0(n932), .A1(n369), .B0(n930), .B1(n347), .Y(n359) );
  CMPR32X1 U914 ( .A(n350), .B(n349), .C(n348), .CO(n996), .S(n380) );
  OAI22X1 U915 ( .A0(n951), .A1(n354), .B0(n353), .B1(n1006), .Y(n358) );
  OAI22X1 U916 ( .A0(n832), .A1(n356), .B0(n974), .B1(n355), .Y(n357) );
  CMPR32X1 U917 ( .A(n361), .B(n360), .C(n359), .CO(n366), .S(n386) );
  CMPR32X1 U918 ( .A(n367), .B(n366), .C(n365), .CO(n994), .S(n385) );
  OAI22XL U919 ( .A0(n828), .A1(n391), .B0(n934), .B1(n368), .Y(n396) );
  XNOR2X1 U920 ( .A(n9), .B(n402), .Y(n370) );
  XNOR2XL U921 ( .A(n894), .B(n848), .Y(n392) );
  XNOR2XL U922 ( .A(n6), .B(n883), .Y(n390) );
  ADDHXL U923 ( .A(n374), .B(n373), .CO(n387), .S(n1070) );
  CMPR32X1 U924 ( .A(n377), .B(n376), .C(n375), .CO(n365), .S(n397) );
  NOR2XL U925 ( .A(n382), .B(n381), .Y(mult_x_1_n306) );
  NAND2XL U926 ( .A(n382), .B(n381), .Y(mult_x_1_n307) );
  CMPR32X1 U927 ( .A(n385), .B(n384), .C(n383), .CO(n381), .S(n401) );
  NOR2BX1 U928 ( .AN(n402), .B(n930), .Y(n1077) );
  OAI22XL U929 ( .A0(n828), .A1(n458), .B0(n934), .B1(n391), .Y(n1093) );
  OAI22XL U930 ( .A0(n8), .A1(n461), .B0(n947), .B1(n392), .Y(n1092) );
  CMPR32X1 U931 ( .A(n396), .B(n395), .C(n394), .CO(n399), .S(n1081) );
  CMPR32X1 U932 ( .A(n399), .B(n398), .C(n397), .CO(n384), .S(n1067) );
  NOR2XL U933 ( .A(n401), .B(n400), .Y(mult_x_1_n314) );
  NAND2XL U934 ( .A(n401), .B(n400), .Y(mult_x_1_n315) );
  XNOR2XL U935 ( .A(n612), .B(n848), .Y(n405) );
  OAI22X1 U936 ( .A0(n951), .A1(n405), .B0(n473), .B1(n1006), .Y(n466) );
  XNOR2XL U937 ( .A(n612), .B(n896), .Y(n409) );
  OAI22XL U938 ( .A0(n951), .A1(n409), .B0(n405), .B1(n1006), .Y(n413) );
  XNOR2XL U939 ( .A(n900), .B(n402), .Y(n406) );
  XNOR2X1 U940 ( .A(n900), .B(n905), .Y(n475) );
  OAI22X1 U941 ( .A0(n951), .A1(n434), .B0(n409), .B1(n1006), .Y(n422) );
  OAI22X1 U942 ( .A0(n8), .A1(n504), .B0(n947), .B1(n411), .Y(n421) );
  CMPR32X1 U943 ( .A(n414), .B(n413), .C(n412), .CO(n489), .S(n415) );
  CMPR32X1 U944 ( .A(n417), .B(n416), .C(n415), .CO(n454), .S(n453) );
  NOR2XL U945 ( .A(n1147), .B(n1162), .Y(n457) );
  OAI22X1 U946 ( .A0(n951), .A1(n428), .B0(n435), .B1(n1006), .Y(n439) );
  OAI22X1 U947 ( .A0(n928), .A1(n429), .B0(n926), .B1(n437), .Y(n438) );
  OAI21XL U948 ( .A0(n1216), .A1(n1213), .B0(n1214), .Y(n1211) );
  CMPR22X1 U949 ( .A(n439), .B(n438), .CO(n441), .S(n433) );
  CMPR32X1 U950 ( .A(n446), .B(n445), .C(n444), .CO(n452), .S(n451) );
  CMPR32X1 U951 ( .A(n449), .B(n448), .C(n447), .CO(n450), .S(n442) );
  OAI21XL U952 ( .A0(n1208), .A1(n1205), .B0(n1206), .Y(n1146) );
  NAND2XL U953 ( .A(n455), .B(n454), .Y(n1148) );
  OAI21XL U954 ( .A0(n1147), .A1(n1163), .B0(n1148), .Y(n456) );
  AOI21XL U955 ( .A0(n457), .A1(n1146), .B0(n456), .Y(n498) );
  OAI22X1 U956 ( .A0(n951), .A1(n472), .B0(n469), .B1(n1006), .Y(n1074) );
  OAI22X1 U957 ( .A0(n913), .A1(n471), .B0(n968), .B1(n470), .Y(n1073) );
  OAI22XL U958 ( .A0(n828), .A1(n475), .B0(n934), .B1(n474), .Y(n476) );
  CMPR32X1 U959 ( .A(n478), .B(n477), .C(n476), .CO(n1094), .S(n487) );
  CMPR32X1 U960 ( .A(n483), .B(n482), .C(n481), .CO(n1115), .S(n485) );
  CMPR32X1 U961 ( .A(n487), .B(n486), .C(n485), .CO(n493), .S(n492) );
  NAND2XL U962 ( .A(n484), .B(n1227), .Y(n497) );
  OAI21XL U963 ( .A0(n498), .A1(n497), .B0(n496), .Y(mult_x_1_n331) );
  CMPR32X1 U964 ( .A(n502), .B(n501), .C(n500), .CO(n194), .S(mult_x_1_n442)
         );
  NOR2XL U965 ( .A(n519), .B(n503), .Y(n526) );
  CMPR32X1 U966 ( .A(n509), .B(n508), .C(n507), .CO(n79), .S(n1230) );
  CMPR32X1 U967 ( .A(n512), .B(n511), .C(n510), .CO(n80), .S(n1229) );
  XNOR2X1 U968 ( .A(n900), .B(n1048), .Y(n521) );
  XNOR2X1 U969 ( .A(n1012), .B(n823), .Y(n518) );
  OAI22X1 U970 ( .A0(n832), .A1(n551), .B0(n974), .B1(n518), .Y(n555) );
  INVXL U971 ( .A(n525), .Y(n553) );
  CMPR32X1 U972 ( .A(n526), .B(n525), .C(n524), .CO(n1231), .S(n563) );
  CMPR32X1 U973 ( .A(n529), .B(n528), .C(n527), .CO(n538), .S(n562) );
  ADDFHX1 U974 ( .A(n538), .B(n537), .CI(n536), .CO(n534), .S(mult_x_1_n472)
         );
  CMPR32X1 U975 ( .A(n541), .B(n540), .C(n539), .CO(n537), .S(n561) );
  XNOR2X1 U976 ( .A(n1049), .B(n852), .Y(n544) );
  NOR2XL U977 ( .A(n519), .B(n544), .Y(n600) );
  XNOR2XL U978 ( .A(n886), .B(A[24]), .Y(n583) );
  XNOR2XL U979 ( .A(n1012), .B(n881), .Y(n585) );
  CMPR32X1 U980 ( .A(n555), .B(n554), .C(n553), .CO(n539), .S(n578) );
  CMPR32X1 U981 ( .A(n558), .B(n557), .C(n556), .CO(n564), .S(n577) );
  CMPR32X1 U982 ( .A(n561), .B(n560), .C(n559), .CO(mult_x_1_n483), .S(
        mult_x_1_n484) );
  CMPR32X1 U983 ( .A(n564), .B(n563), .C(n562), .CO(n536), .S(mult_x_1_n486)
         );
  CMPR32X1 U984 ( .A(n567), .B(n566), .C(n565), .CO(n560), .S(n582) );
  NOR2XL U985 ( .A(n519), .B(n569), .Y(n622) );
  XNOR2X1 U986 ( .A(n1052), .B(n852), .Y(n591) );
  CMPR32X1 U987 ( .A(n573), .B(n572), .C(n571), .CO(n565), .S(n593) );
  CMPR32X1 U988 ( .A(n576), .B(n575), .C(n574), .CO(n579), .S(n592) );
  CMPR32X1 U989 ( .A(n582), .B(n581), .C(n580), .CO(mult_x_1_n495), .S(
        mult_x_1_n496) );
  XNOR2XL U990 ( .A(n1027), .B(n850), .Y(n620) );
  OAI22XL U991 ( .A0(n832), .A1(n620), .B0(n974), .B1(n585), .Y(n597) );
  INVXL U992 ( .A(n599), .Y(n595) );
  XNOR2X1 U993 ( .A(n1052), .B(n893), .Y(n631) );
  CMPR32X1 U994 ( .A(n594), .B(n593), .C(n592), .CO(n581), .S(n605) );
  CMPR32X1 U995 ( .A(n597), .B(n596), .C(n595), .CO(n1154), .S(n646) );
  CMPR32X1 U996 ( .A(n600), .B(n599), .C(n598), .CO(n566), .S(n1153) );
  CMPR32X1 U997 ( .A(n603), .B(n602), .C(n601), .CO(n1152), .S(n645) );
  CMPR32X1 U998 ( .A(n606), .B(n605), .C(n604), .CO(mult_x_1_n509), .S(
        mult_x_1_n510) );
  CMPR32X1 U999 ( .A(n611), .B(n610), .C(n609), .CO(n647), .S(n658) );
  OAI22X1 U1000 ( .A0(n951), .A1(n615), .B0(n613), .B1(n1006), .Y(n627) );
  OAI22X1 U1001 ( .A0(n951), .A1(n675), .B0(n615), .B1(n1006), .Y(n674) );
  XNOR2X1 U1002 ( .A(n1049), .B(A[8]), .Y(n616) );
  XNOR2X1 U1003 ( .A(B[16]), .B(n899), .Y(n619) );
  NOR2XL U1004 ( .A(n519), .B(n619), .Y(n634) );
  XNOR2X1 U1005 ( .A(n1027), .B(n885), .Y(n632) );
  CMPR32X1 U1006 ( .A(n623), .B(n622), .C(n621), .CO(n594), .S(n643) );
  CMPR32X1 U1007 ( .A(n635), .B(n634), .C(n633), .CO(n644), .S(n661) );
  CMPR32X1 U1008 ( .A(n638), .B(n637), .C(n636), .CO(n642), .S(n660) );
  CMPR32X1 U1009 ( .A(n641), .B(n640), .C(n639), .CO(mult_x_1_n523), .S(
        mult_x_1_n524) );
  CMPR32X1 U1010 ( .A(n644), .B(n643), .C(n642), .CO(mult_x_1_n525), .S(n640)
         );
  CMPR32X1 U1011 ( .A(n647), .B(n646), .C(n645), .CO(n606), .S(mult_x_1_n528)
         );
  XNOR2X1 U1012 ( .A(n9), .B(n885), .Y(n666) );
  CMPR32X1 U1013 ( .A(n653), .B(n652), .C(n651), .CO(n659), .S(n687) );
  CMPR32X1 U1014 ( .A(n656), .B(n655), .C(n654), .CO(n657), .S(n686) );
  CMPR32X1 U1015 ( .A(n659), .B(n658), .C(n657), .CO(n641), .S(n664) );
  CMPR32X1 U1016 ( .A(n662), .B(n661), .C(n660), .CO(n639), .S(n663) );
  CMPR32X1 U1017 ( .A(n665), .B(n664), .C(n663), .CO(mult_x_1_n539), .S(
        mult_x_1_n540) );
  XNOR2X1 U1018 ( .A(n9), .B(n852), .Y(n695) );
  CMPR32X1 U1019 ( .A(n671), .B(n670), .C(n669), .CO(n688), .S(n716) );
  XNOR2X1 U1020 ( .A(n1027), .B(n893), .Y(n708) );
  CMPR32X1 U1021 ( .A(n682), .B(n681), .C(n680), .CO(n662), .S(n693) );
  CMPR32X1 U1022 ( .A(n685), .B(n684), .C(n683), .CO(n692), .S(n715) );
  CMPR32X1 U1023 ( .A(n691), .B(n690), .C(n689), .CO(mult_x_1_n555), .S(
        mult_x_1_n556) );
  CMPR32X1 U1024 ( .A(n694), .B(n693), .C(n692), .CO(mult_x_1_n557), .S(n690)
         );
  XNOR2X1 U1025 ( .A(n9), .B(n893), .Y(n724) );
  CMPR32X1 U1026 ( .A(n700), .B(n699), .C(n698), .CO(n717), .S(n745) );
  ADDHXL U1027 ( .A(n703), .B(n702), .CO(n683), .S(n713) );
  OAI22X1 U1028 ( .A0(n951), .A1(n733), .B0(n704), .B1(n1006), .Y(n732) );
  XNOR2X1 U1029 ( .A(B[16]), .B(n848), .Y(n705) );
  XNOR2X1 U1030 ( .A(n1027), .B(n899), .Y(n737) );
  CMPR32X1 U1031 ( .A(n711), .B(n710), .C(n709), .CO(n694), .S(n722) );
  CMPR32X1 U1032 ( .A(n714), .B(n712), .C(n713), .CO(n721), .S(n744) );
  CMPR32X1 U1033 ( .A(n720), .B(n719), .C(n718), .CO(mult_x_1_n571), .S(
        mult_x_1_n572) );
  CMPR32X1 U1034 ( .A(n723), .B(n722), .C(n721), .CO(mult_x_1_n573), .S(n719)
         );
  XNOR2X1 U1035 ( .A(n9), .B(n899), .Y(n753) );
  CMPR32X1 U1036 ( .A(n729), .B(n728), .C(n727), .CO(n746), .S(n776) );
  NOR2XL U1037 ( .A(n519), .B(n734), .Y(n761) );
  XNOR2X1 U1038 ( .A(n1027), .B(n898), .Y(n768) );
  CMPR32X1 U1039 ( .A(n740), .B(n739), .C(n738), .CO(n723), .S(n751) );
  CMPR32X1 U1040 ( .A(n743), .B(n742), .C(n741), .CO(n750), .S(n775) );
  CMPR32X1 U1041 ( .A(n749), .B(n748), .C(n747), .CO(mult_x_1_n587), .S(
        mult_x_1_n588) );
  CMPR32X1 U1042 ( .A(n752), .B(n751), .C(n750), .CO(mult_x_1_n589), .S(n748)
         );
  CMPR32X1 U1043 ( .A(n759), .B(n758), .C(n757), .CO(n777), .S(n807) );
  ADDHXL U1044 ( .A(n762), .B(n761), .CO(n741), .S(n773) );
  OAI22X1 U1045 ( .A0(n825), .A1(n795), .B0(n764), .B1(n1006), .Y(n793) );
  XNOR2X1 U1046 ( .A(n1027), .B(A[8]), .Y(n799) );
  OAI22XL U1047 ( .A0(n832), .A1(n799), .B0(n974), .B1(n768), .Y(n800) );
  CMPR32X1 U1048 ( .A(n771), .B(n770), .C(n769), .CO(n752), .S(n782) );
  CMPR32X1 U1049 ( .A(n774), .B(n772), .C(n773), .CO(n781), .S(n806) );
  CMPR32X1 U1050 ( .A(n777), .B(n776), .C(n775), .CO(n749), .S(n778) );
  CMPR32X1 U1051 ( .A(n780), .B(n779), .C(n778), .CO(mult_x_1_n603), .S(
        mult_x_1_n604) );
  CMPR32X1 U1052 ( .A(n783), .B(n782), .C(n781), .CO(mult_x_1_n605), .S(n779)
         );
  XNOR2X1 U1053 ( .A(n9), .B(A[8]), .Y(n815) );
  CMPR32X1 U1054 ( .A(n790), .B(n789), .C(n788), .CO(n808), .S(n840) );
  XNOR2X1 U1055 ( .A(B[16]), .B(n888), .Y(n796) );
  XNOR2X1 U1056 ( .A(n1027), .B(n884), .Y(n831) );
  CMPR32X1 U1057 ( .A(n802), .B(n801), .C(n800), .CO(n783), .S(n813) );
  CMPR32X1 U1058 ( .A(n805), .B(n804), .C(n803), .CO(n812), .S(n839) );
  CMPR32X1 U1059 ( .A(n808), .B(n807), .C(n806), .CO(n780), .S(n809) );
  CMPR32X1 U1060 ( .A(n811), .B(n810), .C(n809), .CO(mult_x_1_n619), .S(
        mult_x_1_n620) );
  CMPR32X1 U1061 ( .A(n814), .B(n813), .C(n812), .CO(mult_x_1_n621), .S(n810)
         );
  XNOR2X1 U1062 ( .A(n9), .B(n884), .Y(n849) );
  XNOR2X1 U1063 ( .A(n1052), .B(n888), .Y(n902) );
  CMPR32X1 U1064 ( .A(n819), .B(n818), .C(n817), .CO(n841), .S(n873) );
  ADDHXL U1065 ( .A(n822), .B(n821), .CO(n803), .S(n837) );
  OAI22X1 U1066 ( .A0(n825), .A1(n861), .B0(n824), .B1(n1006), .Y(n859) );
  XNOR2X1 U1067 ( .A(n1027), .B(n848), .Y(n856) );
  CMPR32X1 U1068 ( .A(n835), .B(n834), .C(n833), .CO(n814), .S(n846) );
  CMPR32X1 U1069 ( .A(n838), .B(n836), .C(n837), .CO(n845), .S(n872) );
  CMPR32X1 U1070 ( .A(n841), .B(n840), .C(n839), .CO(n811), .S(n842) );
  CMPR32X1 U1071 ( .A(n844), .B(n843), .C(n842), .CO(mult_x_1_n635), .S(
        mult_x_1_n636) );
  CMPR32X1 U1072 ( .A(n847), .B(n846), .C(n845), .CO(mult_x_1_n637), .S(n843)
         );
  XNOR2X1 U1073 ( .A(n9), .B(n848), .Y(n897) );
  XNOR2X1 U1074 ( .A(n1027), .B(n896), .Y(n907) );
  CMPR32X1 U1075 ( .A(n865), .B(n864), .C(n863), .CO(n880), .S(n917) );
  CMPR32X1 U1076 ( .A(n868), .B(n867), .C(n866), .CO(n847), .S(n879) );
  CMPR32X1 U1077 ( .A(n871), .B(n870), .C(n869), .CO(n878), .S(n916) );
  CMPR32X1 U1078 ( .A(n874), .B(n873), .C(n872), .CO(n844), .S(n875) );
  CMPR32X1 U1079 ( .A(n877), .B(n876), .C(n875), .CO(mult_x_1_n651), .S(
        mult_x_1_n652) );
  CMPR32X1 U1080 ( .A(n880), .B(n879), .C(n878), .CO(mult_x_1_n653), .S(n876)
         );
  XNOR2X1 U1081 ( .A(n1052), .B(n883), .Y(n903) );
  XNOR2X1 U1082 ( .A(n1027), .B(n888), .Y(n973) );
  XNOR2X1 U1083 ( .A(n1027), .B(n889), .Y(n908) );
  CMPR32X1 U1084 ( .A(n892), .B(n891), .C(n890), .CO(n918), .S(n1132) );
  XNOR2XL U1085 ( .A(n9), .B(n896), .Y(n929) );
  OAI22XL U1086 ( .A0(n904), .A1(n903), .B0(n1054), .B1(n902), .Y(n1195) );
  XNOR2X1 U1087 ( .A(B[16]), .B(n905), .Y(n906) );
  ADDHXL U1088 ( .A(n915), .B(n914), .CO(n869), .S(n1196) );
  CMPR32X1 U1089 ( .A(n918), .B(n917), .C(n916), .CO(n877), .S(n919) );
  CMPR32X1 U1090 ( .A(n924), .B(n923), .C(n922), .CO(n920), .S(mult_x_1_n686)
         );
  OAI22XL U1091 ( .A0(n932), .A1(n931), .B0(n930), .B1(n929), .Y(n944) );
  CMPR32X1 U1092 ( .A(n939), .B(n938), .C(n937), .CO(n1133), .S(n1136) );
  CMPR32X1 U1093 ( .A(n942), .B(n941), .C(n940), .CO(n924), .S(n1135) );
  CMPR32X1 U1094 ( .A(n945), .B(n944), .C(n943), .CO(n1137), .S(n999) );
  CMPR32X1 U1095 ( .A(n956), .B(n955), .C(n954), .CO(n960), .S(n959) );
  CMPR32X1 U1096 ( .A(n959), .B(n958), .C(n957), .CO(n997), .S(n1005) );
  CMPR32X1 U1097 ( .A(n962), .B(n961), .C(n960), .CO(n990), .S(n998) );
  XNOR2X1 U1098 ( .A(n1052), .B(n402), .Y(n972) );
  CMPR32X1 U1099 ( .A(n978), .B(n977), .C(n976), .CO(n993), .S(n957) );
  CMPR32X1 U1100 ( .A(n981), .B(n980), .C(n979), .CO(n1129), .S(n992) );
  CMPR32X1 U1101 ( .A(n984), .B(n983), .C(n982), .CO(n991), .S(n995) );
  CMPR32X1 U1102 ( .A(n1002), .B(n1001), .C(n1000), .CO(mult_x_1_n711), .S(
        mult_x_1_n712) );
  CMPR32X1 U1103 ( .A(n1017), .B(n1016), .C(n1015), .CO(n1029), .S(n1036) );
  CMPR32X1 U1104 ( .A(n1020), .B(n1019), .C(n1018), .CO(n1037), .S(n1035) );
  CMPR32X1 U1105 ( .A(n1023), .B(n1022), .C(n1021), .CO(n1104), .S(n1039) );
  OAI22X1 U1106 ( .A0(n832), .A1(n1028), .B0(n974), .B1(n1045), .Y(n1059) );
  CMPR32X1 U1107 ( .A(n1031), .B(n1030), .C(n1029), .CO(n1102), .S(n1038) );
  CMPR32X1 U1108 ( .A(n1036), .B(n1035), .C(n1034), .CO(n1087), .S(n193) );
  CMPR32X1 U1109 ( .A(n1039), .B(n1038), .C(n1037), .CO(n1033), .S(n1086) );
  CMPR32X1 U1110 ( .A(n1043), .B(n1042), .C(n1041), .CO(n1106), .S(n1103) );
  CMPR32X1 U1111 ( .A(n1059), .B(n1058), .C(n1057), .CO(n1060), .S(n1105) );
  CMPR32X1 U1112 ( .A(n1062), .B(n1061), .C(n1060), .S(n1063) );
  CMPR32X1 U1113 ( .A(n1069), .B(n1068), .C(n1067), .CO(n400), .S(n1085) );
  CMPR32X1 U1114 ( .A(n1072), .B(n1071), .C(n1070), .CO(n398), .S(n1090) );
  CMPR22X1 U1115 ( .A(n1074), .B(n1073), .CO(n1099), .S(n1095) );
  CMPR32X1 U1116 ( .A(n1077), .B(n1076), .C(n1075), .CO(n1083), .S(n1098) );
  CMPR32X1 U1117 ( .A(n1080), .B(n1079), .C(n1078), .CO(n1097), .S(n1116) );
  CMPR32X1 U1118 ( .A(n1083), .B(n1082), .C(n1081), .CO(n1068), .S(n1088) );
  CMPR32X1 U1119 ( .A(n1090), .B(n1089), .C(n1088), .CO(n1084), .S(n1101) );
  CMPR32X1 U1120 ( .A(n1093), .B(n1092), .C(n1091), .CO(n1082), .S(n1113) );
  CMPR32X1 U1121 ( .A(n1096), .B(n1095), .C(n1094), .CO(n1112), .S(n1114) );
  CMPR32X1 U1122 ( .A(n1099), .B(n1098), .C(n1097), .CO(n1089), .S(n1111) );
  CMPR32X1 U1123 ( .A(n1104), .B(n1103), .C(n1102), .CO(n1110), .S(n1032) );
  CMPR32X1 U1124 ( .A(n1107), .B(n1106), .C(n1105), .CO(n1064), .S(n1109) );
  CMPR32X1 U1125 ( .A(n1113), .B(n1112), .C(n1111), .CO(n1100), .S(n1118) );
  CMPR32X1 U1126 ( .A(n1116), .B(n1115), .C(n1114), .CO(n1117), .S(n494) );
  OAI21XL U1127 ( .A0(n1123), .A1(n1122), .B0(n1121), .Y(n1128) );
  INVXL U1128 ( .A(n1124), .Y(n1126) );
  CMPR32X1 U1129 ( .A(n1134), .B(n1133), .C(n1132), .CO(n921), .S(n1139) );
  CMPR32X1 U1130 ( .A(n1137), .B(n1136), .C(n1135), .CO(n1138), .S(n987) );
  CMPR32X1 U1131 ( .A(n1140), .B(n1139), .C(n1138), .CO(mult_x_1_n683), .S(
        mult_x_1_n684) );
  AOI21XL U1132 ( .A0(n1192), .A1(n1190), .B0(n1142), .Y(n1145) );
  OAI21XL U1133 ( .A0(n1165), .A1(n1162), .B0(n1163), .Y(n1151) );
  CMPR32X1 U1134 ( .A(n1154), .B(n1153), .C(n1152), .CO(mult_x_1_n513), .S(
        n604) );
  AOI21XL U1135 ( .A0(n1177), .A1(n1156), .B0(n1155), .Y(n1157) );
  OAI21XL U1136 ( .A0(n1180), .A1(n1158), .B0(n1157), .Y(n1161) );
  OAI21XL U1137 ( .A0(n1235), .A1(n1238), .B0(n1236), .Y(n1175) );
  AOI21XL U1138 ( .A0(n1177), .A1(n1170), .B0(n1169), .Y(n1171) );
  OAI21XL U1139 ( .A0(n1180), .A1(n1172), .B0(n1171), .Y(n1173) );
  AOI21XL U1140 ( .A0(n1177), .A1(n1176), .B0(n1175), .Y(n1178) );
  OAI21XL U1141 ( .A0(n1180), .A1(n1179), .B0(n1178), .Y(n1183) );
  XOR2XL U1142 ( .A(n1253), .B(n1251), .Y(PRODUCT[9]) );
  INVXL U1143 ( .A(n1249), .Y(n1184) );
  NAND2XL U1144 ( .A(n1184), .B(n1250), .Y(n1185) );
  XOR2XL U1145 ( .A(n1186), .B(n1185), .Y(PRODUCT[10]) );
  OAI21XL U1146 ( .A0(n1186), .A1(n1249), .B0(n1250), .Y(n1189) );
  INVXL U1147 ( .A(n1247), .Y(n1187) );
  NAND2XL U1148 ( .A(n1190), .B(n1246), .Y(n1191) );
  CMPR32X1 U1149 ( .A(n1195), .B(n1194), .C(n1193), .CO(n1204), .S(n923) );
  CMPR32X1 U1150 ( .A(n1198), .B(n1197), .C(n1196), .CO(n1203), .S(n922) );
  CMPR32X1 U1151 ( .A(n1201), .B(n1200), .C(n1199), .CO(n874), .S(n1202) );
  CMPR32X1 U1152 ( .A(n1204), .B(n1203), .C(n1202), .CO(mult_x_1_n669), .S(
        mult_x_1_n670) );
  AOI21XL U1153 ( .A0(n1228), .A1(n1227), .B0(n1226), .Y(mult_x_1_n338) );
  CMPR32X1 U1154 ( .A(n1231), .B(n1230), .C(n1229), .CO(n535), .S(
        mult_x_1_n474) );
endmodule


module FFT2048_DW02_mult_2_stage_J1_10 ( A, B, TC, CLK, PRODUCT );
  input [25:0] A;
  input [16:0] B;
  output [42:0] PRODUCT;
  input TC, CLK;
  wire   n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, mult_x_1_n601, mult_x_1_n586, mult_x_1_n321,
         mult_x_1_n316, mult_x_1_n309, mult_x_1_n307, mult_x_1_n306,
         mult_x_1_n296, mult_x_1_n295, mult_x_1_n293, mult_x_1_n292,
         mult_x_1_n287, mult_x_1_n286, mult_x_1_n282, mult_x_1_n281,
         mult_x_1_n277, mult_x_1_n276, mult_x_1_n274, mult_x_1_n273,
         mult_x_1_n266, mult_x_1_n265, mult_x_1_n263, mult_x_1_n262,
         mult_x_1_n245, mult_x_1_n244, mult_x_1_n234, mult_x_1_n233,
         mult_x_1_n227, mult_x_1_n226, mult_x_1_n216, mult_x_1_n215,
         mult_x_1_n207, mult_x_1_n206, mult_x_1_n198, mult_x_1_n197,
         mult_x_1_n195, mult_x_1_n194, mult_x_1_n184, mult_x_1_n183,
         mult_x_1_n177, mult_x_1_n176, mult_x_1_n170, mult_x_1_n169,
         mult_x_1_n161, mult_x_1_n160, mult_x_1_n152, mult_x_1_n151,
         mult_x_1_n137, mult_x_1_n136, mult_x_1_n130, mult_x_1_n129,
         mult_x_1_n121, mult_x_1_n120, mult_x_1_n110, mult_x_1_n109,
         mult_x_1_n86, mult_x_1_n85, mult_x_1_n84, mult_x_1_n83, mult_x_1_n58,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311;

  DFFHQXL mult_x_1_clk_r_REG11_S1 ( .D(mult_x_1_n194), .CK(CLK), .Q(n1274) );
  DFFHQXL mult_x_1_clk_r_REG15_S1 ( .D(mult_x_1_n176), .CK(CLK), .Q(n1270) );
  DFFHQXL mult_x_1_clk_r_REG13_S1 ( .D(mult_x_1_n183), .CK(CLK), .Q(n1272) );
  DFFHQX4 mult_x_1_clk_r_REG1_S1 ( .D(mult_x_1_n233), .CK(CLK), .Q(n1284) );
  DFFHQX4 mult_x_1_clk_r_REG34_S1 ( .D(mult_x_1_n601), .CK(CLK), .Q(n1311) );
  DFFHQX4 mult_x_1_clk_r_REG56_S1 ( .D(mult_x_1_n309), .CK(CLK), .Q(n1308) );
  DFFHQX4 mult_x_1_clk_r_REG50_S1 ( .D(mult_x_1_n296), .CK(CLK), .Q(n1307) );
  DFFHQX4 mult_x_1_clk_r_REG51_S1 ( .D(mult_x_1_n295), .CK(CLK), .Q(n1302) );
  DFFHQX4 mult_x_1_clk_r_REG48_S1 ( .D(mult_x_1_n292), .CK(CLK), .Q(n1300) );
  DFFHQX4 mult_x_1_clk_r_REG44_S1 ( .D(mult_x_1_n281), .CK(CLK), .Q(n1296) );
  DFFHQX4 mult_x_1_clk_r_REG37_S1 ( .D(mult_x_1_n266), .CK(CLK), .Q(n1291) );
  DFFHQXL mult_x_1_clk_r_REG6_S1 ( .D(mult_x_1_n207), .CK(CLK), .Q(n1279) );
  DFFHQX4 mult_x_1_clk_r_REG47_S1 ( .D(mult_x_1_n293), .CK(CLK), .Q(n1301) );
  DFFHQXL mult_x_1_clk_r_REG9_S1 ( .D(mult_x_1_n197), .CK(CLK), .Q(n1276) );
  DFFHQXL mult_x_1_clk_r_REG20_S1 ( .D(mult_x_1_n152), .CK(CLK), .Q(n1265) );
  DFFHQXL mult_x_1_clk_r_REG14_S1 ( .D(mult_x_1_n177), .CK(CLK), .Q(n1271) );
  DFFHQXL mult_x_1_clk_r_REG18_S1 ( .D(mult_x_1_n161), .CK(CLK), .Q(n1267) );
  DFFHQXL mult_x_1_clk_r_REG16_S1 ( .D(mult_x_1_n170), .CK(CLK), .Q(n1269) );
  DFFHQXL mult_x_1_clk_r_REG8_S1 ( .D(mult_x_1_n198), .CK(CLK), .Q(n1277) );
  DFFHQXL clk_r_REG62_S1 ( .D(n1326), .CK(CLK), .Q(PRODUCT[9]) );
  DFFHQXL clk_r_REG61_S1 ( .D(n1325), .CK(CLK), .Q(PRODUCT[10]) );
  DFFHQXL mult_x_1_clk_r_REG4_S1 ( .D(mult_x_1_n216), .CK(CLK), .Q(n1281) );
  DFFHQXL mult_x_1_clk_r_REG58_S1 ( .D(mult_x_1_n316), .CK(CLK), .Q(n1309) );
  DFFHQXL mult_x_1_clk_r_REG2_S1 ( .D(mult_x_1_n227), .CK(CLK), .Q(n1283) );
  DFFHQXL mult_x_1_clk_r_REG49_S1 ( .D(mult_x_1_n83), .CK(CLK), .Q(n1303) );
  DFFHQXL clk_r_REG59_S1 ( .D(n1324), .CK(CLK), .Q(PRODUCT[11]) );
  DFFHQXL clk_r_REG71_S1 ( .D(n1335), .CK(CLK), .Q(PRODUCT[0]) );
  DFFHQXL mult_x_1_clk_r_REG26_S1 ( .D(mult_x_1_n121), .CK(CLK), .Q(n1259) );
  DFFHQXL mult_x_1_clk_r_REG19_S1 ( .D(mult_x_1_n160), .CK(CLK), .Q(n1266) );
  DFFHQXL mult_x_1_clk_r_REG12_S1 ( .D(mult_x_1_n184), .CK(CLK), .Q(n1273) );
  DFFHQX4 mult_x_1_clk_r_REG36_S1 ( .D(mult_x_1_n262), .CK(CLK), .Q(n1288) );
  DFFHQXL mult_x_1_clk_r_REG60_S1 ( .D(mult_x_1_n321), .CK(CLK), .Q(n1254) );
  DFFHQX4 mult_x_1_clk_r_REG3_S1 ( .D(mult_x_1_n226), .CK(CLK), .Q(n1282) );
  DFFHQX4 mult_x_1_clk_r_REG32_S1 ( .D(mult_x_1_n244), .CK(CLK), .Q(n1286) );
  DFFHQX1 mult_x_1_clk_r_REG38_S1 ( .D(mult_x_1_n265), .CK(CLK), .Q(n1290) );
  DFFHQXL clk_r_REG63_S1 ( .D(n1327), .CK(CLK), .Q(PRODUCT[8]) );
  DFFHQXL clk_r_REG64_S1 ( .D(n1328), .CK(CLK), .Q(PRODUCT[7]) );
  DFFHQXL clk_r_REG65_S1 ( .D(n1329), .CK(CLK), .Q(PRODUCT[6]) );
  DFFHQXL clk_r_REG66_S1 ( .D(n1330), .CK(CLK), .Q(PRODUCT[5]) );
  DFFHQXL clk_r_REG67_S1 ( .D(n1331), .CK(CLK), .Q(PRODUCT[4]) );
  DFFHQXL clk_r_REG68_S1 ( .D(n1332), .CK(CLK), .Q(PRODUCT[3]) );
  DFFHQXL clk_r_REG69_S1 ( .D(n1333), .CK(CLK), .Q(PRODUCT[2]) );
  DFFHQXL clk_r_REG70_S1 ( .D(n1334), .CK(CLK), .Q(PRODUCT[1]) );
  DFFHQX1 mult_x_1_clk_r_REG5_S1 ( .D(mult_x_1_n215), .CK(CLK), .Q(n1280) );
  DFFHQXL mult_x_1_clk_r_REG57_S1 ( .D(mult_x_1_n86), .CK(CLK), .Q(n1306) );
  DFFHQX1 mult_x_1_clk_r_REG55_S1 ( .D(mult_x_1_n85), .CK(CLK), .Q(n1305) );
  DFFHQXL mult_x_1_clk_r_REG22_S1 ( .D(mult_x_1_n137), .CK(CLK), .Q(n1263) );
  DFFHQXL mult_x_1_clk_r_REG24_S1 ( .D(mult_x_1_n130), .CK(CLK), .Q(n1261) );
  DFFHQXL mult_x_1_clk_r_REG25_S1 ( .D(mult_x_1_n129), .CK(CLK), .Q(n1260) );
  DFFHQXL mult_x_1_clk_r_REG27_S1 ( .D(mult_x_1_n120), .CK(CLK), .Q(n1258) );
  DFFHQXL mult_x_1_clk_r_REG28_S1 ( .D(mult_x_1_n110), .CK(CLK), .Q(n1257) );
  DFFHQXL mult_x_1_clk_r_REG29_S1 ( .D(mult_x_1_n109), .CK(CLK), .Q(n1256) );
  DFFHQXL mult_x_1_clk_r_REG30_S1 ( .D(mult_x_1_n58), .CK(CLK), .Q(n1255) );
  DFFHQXL mult_x_1_clk_r_REG53_S1 ( .D(mult_x_1_n307), .CK(CLK), .Q(n1253) );
  DFFHQXL mult_x_1_clk_r_REG54_S1 ( .D(mult_x_1_n306), .CK(CLK), .Q(n1252) );
  DFFHQX1 mult_x_1_clk_r_REG39_S1 ( .D(mult_x_1_n274), .CK(CLK), .Q(n1293) );
  DFFHQXL mult_x_1_clk_r_REG23_S1 ( .D(mult_x_1_n136), .CK(CLK), .Q(n1262) );
  DFFHQXL mult_x_1_clk_r_REG21_S1 ( .D(mult_x_1_n151), .CK(CLK), .Q(n1264) );
  DFFHQXL mult_x_1_clk_r_REG10_S1 ( .D(mult_x_1_n195), .CK(CLK), .Q(n1275) );
  DFFHQXL mult_x_1_clk_r_REG17_S1 ( .D(mult_x_1_n169), .CK(CLK), .Q(n1268) );
  DFFHQXL mult_x_1_clk_r_REG31_S1 ( .D(mult_x_1_n245), .CK(CLK), .Q(n1287) );
  DFFHQX1 mult_x_1_clk_r_REG43_S1 ( .D(mult_x_1_n282), .CK(CLK), .Q(n1297) );
  DFFHQXL mult_x_1_clk_r_REG52_S1 ( .D(mult_x_1_n84), .CK(CLK), .Q(n1304) );
  DFFHQX1 mult_x_1_clk_r_REG46_S1 ( .D(mult_x_1_n286), .CK(CLK), .Q(n1298) );
  DFFHQX1 mult_x_1_clk_r_REG41_S1 ( .D(mult_x_1_n277), .CK(CLK), .Q(n1295) );
  DFFHQX2 mult_x_1_clk_r_REG42_S1 ( .D(mult_x_1_n276), .CK(CLK), .Q(n1294) );
  DFFHQX2 mult_x_1_clk_r_REG45_S1 ( .D(mult_x_1_n287), .CK(CLK), .Q(n1299) );
  DFFHQX2 mult_x_1_clk_r_REG40_S1 ( .D(mult_x_1_n273), .CK(CLK), .Q(n1292) );
  DFFHQX2 mult_x_1_clk_r_REG33_S1 ( .D(mult_x_1_n586), .CK(CLK), .Q(n1310) );
  DFFHQX1 mult_x_1_clk_r_REG7_S1 ( .D(mult_x_1_n206), .CK(CLK), .Q(n1278) );
  DFFHQX1 mult_x_1_clk_r_REG35_S1 ( .D(mult_x_1_n263), .CK(CLK), .Q(n1289) );
  DFFHQXL mult_x_1_clk_r_REG0_S1 ( .D(mult_x_1_n234), .CK(CLK), .Q(n1285) );
  ADDFHX2 U1 ( .A(n627), .B(n626), .CI(n625), .CO(n597), .S(n633) );
  ADDFHX1 U2 ( .A(n892), .B(n891), .CI(n890), .CO(n859), .S(n898) );
  ADDFHX1 U3 ( .A(n813), .B(n812), .CI(n811), .CO(n1083), .S(n818) );
  ADDFHX1 U4 ( .A(n785), .B(n784), .CI(n783), .CO(n1080), .S(n1082) );
  ADDFHX1 U5 ( .A(n850), .B(n849), .CI(n848), .CO(n819), .S(n858) );
  ADDFHX2 U6 ( .A(n807), .B(n806), .CI(n805), .CO(n820), .S(n849) );
  ADDFX2 U7 ( .A(n1055), .B(n1054), .CI(n1053), .CO(n1058), .S(n1057) );
  ADDFHX1 U8 ( .A(n782), .B(n781), .CI(n780), .CO(n785), .S(n811) );
  ADDFHX1 U9 ( .A(n624), .B(n623), .CI(n622), .CO(n627), .S(n664) );
  ADDFHX1 U10 ( .A(n499), .B(n498), .CI(n497), .CO(n485), .S(n545) );
  ADDFHX1 U11 ( .A(n663), .B(n662), .CI(n661), .CO(n666), .S(n704) );
  ADDFHX1 U12 ( .A(n844), .B(n843), .CI(n842), .CO(n860), .S(n891) );
  ADDFHX1 U13 ( .A(n779), .B(n778), .CI(n777), .CO(n1084), .S(n812) );
  ADDFHX1 U14 ( .A(n744), .B(n743), .CI(n742), .CO(n747), .S(n783) );
  ADDFHX1 U15 ( .A(n741), .B(n740), .CI(n739), .CO(n1081), .S(n784) );
  CMPR32X1 U16 ( .A(n568), .B(n567), .C(n566), .CO(n546), .S(n598) );
  ADDFHX2 U17 ( .A(n586), .B(n585), .CI(n584), .CO(n564), .S(n596) );
  ADDFX2 U18 ( .A(n1046), .B(n1045), .CI(n1044), .CO(n1051), .S(n1053) );
  ADDFX2 U19 ( .A(n947), .B(n946), .CI(n945), .CO(n934), .S(n991) );
  CMPR32X1 U20 ( .A(n773), .B(n772), .C(n771), .CO(n782), .S(n809) );
  ADDFHX1 U21 ( .A(n278), .B(n277), .CI(n276), .CO(n284), .S(n283) );
  ADDFHX1 U22 ( .A(n654), .B(n653), .CI(n652), .CO(n663), .S(n702) );
  ADDFHX1 U23 ( .A(n463), .B(n462), .CI(n461), .CO(n455), .S(n498) );
  ADDFHX1 U24 ( .A(n641), .B(n640), .CI(n639), .CO(n621), .S(n659) );
  ADDFHX1 U25 ( .A(n683), .B(n682), .CI(n681), .CO(n660), .S(n699) );
  ADDFX2 U26 ( .A(n694), .B(n693), .CI(n692), .CO(n703), .S(n743) );
  ADDFHX1 U27 ( .A(n724), .B(n723), .CI(n722), .CO(n700), .S(n740) );
  ADDFHX1 U28 ( .A(n735), .B(n734), .CI(n733), .CO(n744), .S(n781) );
  OAI22X1 U29 ( .A0(n966), .A1(n648), .B0(n964), .B1(n610), .Y(n654) );
  OAI22X1 U30 ( .A0(n730), .A1(n966), .B0(n964), .B1(n98), .Y(n735) );
  ADDFHX1 U31 ( .A(n580), .B(n579), .CI(n578), .CO(n586), .S(n626) );
  ADDFX2 U32 ( .A(n534), .B(n533), .CI(n532), .CO(n565), .S(n585) );
  ADDFHX1 U33 ( .A(n801), .B(n800), .CI(n799), .CO(n810), .S(n846) );
  CMPR32X1 U34 ( .A(n1026), .B(n1025), .C(n1024), .CO(n1046), .S(n1043) );
  CMPR32X1 U35 ( .A(n1009), .B(n1008), .C(n1007), .CO(n1023), .S(n1038) );
  XOR2X1 U36 ( .A(n922), .B(n99), .Y(n98) );
  XNOR2X1 U37 ( .A(n1138), .B(A[9]), .Y(n637) );
  ADDFHX1 U38 ( .A(n223), .B(n222), .CI(n221), .CO(n280), .S(n224) );
  ADDFHX1 U39 ( .A(n604), .B(n603), .CI(n602), .CO(n583), .S(n620) );
  CMPR32X1 U40 ( .A(n878), .B(n877), .C(n876), .CO(n889), .S(n916) );
  ADDFX2 U41 ( .A(n185), .B(n184), .CI(n183), .CO(n191), .S(n190) );
  ADDFX2 U42 ( .A(n973), .B(n972), .CI(n971), .CO(n957), .S(n1022) );
  CMPR32X1 U43 ( .A(n997), .B(n996), .C(n995), .CO(n994), .S(n1035) );
  OAI22X1 U44 ( .A0(n1161), .A1(n861), .B0(n8), .B1(n797), .Y(n869) );
  ADDFHX1 U45 ( .A(n929), .B(n928), .CI(n927), .CO(n917), .S(n993) );
  BUFX8 U46 ( .A(n1161), .Y(n7) );
  CLKBUFX8 U47 ( .A(n48), .Y(n8) );
  CLKBUFX8 U48 ( .A(B[13]), .Y(n1120) );
  BUFX4 U49 ( .A(n643), .Y(n962) );
  XOR2X1 U50 ( .A(B[12]), .B(B[13]), .Y(n75) );
  XNOR2X2 U51 ( .A(B[11]), .B(B[12]), .Y(n237) );
  CLKBUFX8 U52 ( .A(n979), .Y(n926) );
  BUFX3 U53 ( .A(n685), .Y(n960) );
  BUFX3 U54 ( .A(n921), .Y(n970) );
  BUFX3 U55 ( .A(n113), .Y(n9) );
  BUFX3 U56 ( .A(n835), .Y(n976) );
  XNOR2X1 U57 ( .A(n445), .B(n444), .Y(PRODUCT[31]) );
  CLKINVX4 U58 ( .A(n47), .Y(n1250) );
  XOR2X1 U59 ( .A(n30), .B(n857), .Y(PRODUCT[20]) );
  AOI21XL U60 ( .A0(n440), .A1(n298), .B0(n297), .Y(n1246) );
  AND2X1 U61 ( .A(n631), .B(n1283), .Y(n632) );
  BUFX3 U62 ( .A(B[5]), .Y(n650) );
  XNOR2XL U63 ( .A(n650), .B(A[1]), .Y(n122) );
  XNOR2XL U64 ( .A(n650), .B(A[7]), .Y(n244) );
  XNOR2X1 U65 ( .A(n1138), .B(A[11]), .Y(n536) );
  XNOR2XL U66 ( .A(n308), .B(n54), .Y(n314) );
  XNOR2XL U67 ( .A(n650), .B(A[13]), .Y(n834) );
  XNOR2XL U68 ( .A(n1138), .B(A[2]), .Y(n872) );
  XNOR2XL U69 ( .A(n924), .B(A[8]), .Y(n977) );
  XNOR2XL U70 ( .A(n1120), .B(A[11]), .Y(n638) );
  XNOR2XL U71 ( .A(n650), .B(A[25]), .Y(n370) );
  XNOR2XL U72 ( .A(n308), .B(n51), .Y(n487) );
  XNOR2XL U73 ( .A(n908), .B(A[13]), .Y(n725) );
  ADDFX2 U74 ( .A(n870), .B(n869), .CI(n868), .CO(n847), .S(n901) );
  XNOR2XL U75 ( .A(n1194), .B(n1193), .Y(n1328) );
  INVX4 U76 ( .A(B[11]), .Y(n308) );
  XOR2XL U77 ( .A(n897), .B(n896), .Y(PRODUCT[19]) );
  OR2X2 U78 ( .A(n283), .B(n282), .Y(n6) );
  XOR2X1 U79 ( .A(n1078), .B(n1077), .Y(n1326) );
  NAND2XL U80 ( .A(n814), .B(n815), .Y(mult_x_1_n263) );
  NAND2X1 U81 ( .A(n192), .B(n191), .Y(n1075) );
  XNOR2X1 U82 ( .A(n520), .B(n519), .Y(n541) );
  NOR2X1 U83 ( .A(n1158), .B(n346), .Y(n374) );
  OAI22XL U84 ( .A0(n962), .A1(n422), .B0(n685), .B1(n415), .Y(n457) );
  NOR2X1 U85 ( .A(n1158), .B(n301), .Y(n322) );
  NOR2X1 U86 ( .A(n1158), .B(n325), .Y(n1105) );
  NOR2X1 U87 ( .A(n1158), .B(n309), .Y(n330) );
  XNOR2X1 U88 ( .A(n1215), .B(n1214), .Y(PRODUCT[39]) );
  OAI22XL U89 ( .A0(n976), .A1(n770), .B0(n9), .B1(n732), .Y(n771) );
  NOR2BX1 U90 ( .AN(A[0]), .B(n960), .Y(n176) );
  NOR2BX1 U91 ( .AN(A[0]), .B(n757), .Y(n117) );
  OAI22X1 U92 ( .A0(n970), .A1(n769), .B0(n968), .B1(n731), .Y(n772) );
  XOR2X1 U93 ( .A(n19), .B(n632), .Y(PRODUCT[26]) );
  NAND2BXL U94 ( .AN(n28), .B(n29), .Y(n101) );
  OAI21XL U95 ( .A0(n1086), .A1(n20), .B0(n41), .Y(n19) );
  NAND2BX1 U96 ( .AN(n714), .B(n554), .Y(n29) );
  NAND2X1 U97 ( .A(n443), .B(n1273), .Y(n444) );
  AND2XL U98 ( .A(n715), .B(n1287), .Y(n65) );
  NAND2BX1 U99 ( .AN(n1252), .B(n1308), .Y(n32) );
  INVXL U100 ( .A(n1303), .Y(n33) );
  NAND2XL U101 ( .A(n551), .B(n550), .Y(mult_x_1_n198) );
  INVX1 U102 ( .A(n64), .Y(n1076) );
  NAND2X1 U103 ( .A(n1056), .B(n1057), .Y(mult_x_1_n307) );
  ADDFHX1 U104 ( .A(n1084), .B(n1083), .CI(n1082), .CO(mult_x_1_n601), .S(n815) );
  NOR2X1 U105 ( .A(n159), .B(n158), .Y(n1190) );
  INVX1 U106 ( .A(n1199), .Y(n85) );
  INVX1 U107 ( .A(n935), .Y(n89) );
  NAND2X1 U108 ( .A(n156), .B(n157), .Y(n1200) );
  ADDFHX1 U109 ( .A(n457), .B(n456), .CI(n455), .CO(n453), .S(n486) );
  AND2X1 U110 ( .A(n195), .B(n196), .Y(n223) );
  NOR2X1 U111 ( .A(n1158), .B(n1119), .Y(n1130) );
  NOR2X1 U112 ( .A(n1158), .B(n1097), .Y(n1117) );
  NOR2BX1 U113 ( .AN(A[0]), .B(n8), .Y(n1003) );
  XNOR2X1 U114 ( .A(n1181), .B(n1180), .Y(PRODUCT[36]) );
  OR2X2 U115 ( .A(n146), .B(n145), .Y(n144) );
  XNOR2X1 U116 ( .A(n1188), .B(n1187), .Y(PRODUCT[37]) );
  XNOR2X1 U117 ( .A(n368), .B(n367), .Y(PRODUCT[33]) );
  XNOR2X1 U118 ( .A(n1198), .B(n1197), .Y(PRODUCT[38]) );
  INVXL U119 ( .A(n976), .Y(n81) );
  OAI22XL U120 ( .A0(n834), .A1(n9), .B0(n835), .B1(n90), .Y(n876) );
  INVXL U121 ( .A(n1250), .Y(n43) );
  CLKINVX3 U122 ( .A(B[15]), .Y(n306) );
  OAI21XL U123 ( .A0(n1250), .A1(n340), .B0(n339), .Y(n342) );
  NAND3XL U124 ( .A(n47), .B(n337), .C(n1173), .Y(n46) );
  XOR2X1 U125 ( .A(n101), .B(n65), .Y(PRODUCT[24]) );
  OAI21XL U126 ( .A0(n1086), .A1(n559), .B0(n558), .Y(n562) );
  NAND2X1 U127 ( .A(n10), .B(n1291), .Y(n1089) );
  NAND2X1 U128 ( .A(n554), .B(n816), .Y(n10) );
  INVX1 U129 ( .A(n27), .Y(n853) );
  BUFX3 U130 ( .A(B[3]), .Y(n919) );
  INVXL U131 ( .A(n713), .Y(n28) );
  CLKINVX3 U132 ( .A(n21), .Y(n26) );
  NAND3X1 U133 ( .A(n21), .B(n17), .C(n855), .Y(n12) );
  INVX1 U134 ( .A(n25), .Y(n23) );
  XNOR2X1 U135 ( .A(n1017), .B(n1016), .Y(PRODUCT[16]) );
  NAND2X1 U136 ( .A(n32), .B(n1253), .Y(n31) );
  NAND2X1 U137 ( .A(n987), .B(n1299), .Y(n988) );
  NAND2X1 U138 ( .A(n895), .B(n1295), .Y(n896) );
  OAI21X1 U139 ( .A0(n1286), .A1(n752), .B0(n1287), .Y(n100) );
  NAND2XL U140 ( .A(n472), .B(n1275), .Y(n473) );
  INVXL U141 ( .A(A[16]), .Y(n51) );
  INVXL U142 ( .A(A[17]), .Y(n52) );
  BUFX2 U143 ( .A(A[14]), .Y(n904) );
  INVX1 U144 ( .A(n1290), .Y(n816) );
  ADDFHX1 U145 ( .A(n991), .B(n990), .CI(n989), .CO(n985), .S(n1014) );
  NAND2X1 U146 ( .A(n1074), .B(n1076), .Y(n95) );
  NAND2XL U147 ( .A(n73), .B(n942), .Y(n72) );
  INVXL U148 ( .A(n62), .Y(n61) );
  NAND2X1 U149 ( .A(n283), .B(n282), .Y(n1068) );
  NAND2XL U150 ( .A(n97), .B(n74), .Y(n73) );
  NAND2XL U151 ( .A(n564), .B(n565), .Y(n60) );
  NOR2X1 U152 ( .A(n1057), .B(n1056), .Y(mult_x_1_n306) );
  ADDFHX1 U153 ( .A(n549), .B(n548), .CI(n547), .CO(n507), .S(n550) );
  NOR2X1 U154 ( .A(n231), .B(n230), .Y(n1069) );
  INVXL U155 ( .A(n565), .Y(n63) );
  ADDFHX1 U156 ( .A(n1020), .B(n1019), .CI(n1018), .CO(n1013), .S(n1037) );
  NAND2BXL U157 ( .AN(n1011), .B(n70), .Y(n69) );
  NAND2XL U158 ( .A(n943), .B(n944), .Y(n96) );
  INVXL U159 ( .A(n943), .Y(n74) );
  INVXL U160 ( .A(n944), .Y(n97) );
  OR2XL U161 ( .A(n1166), .B(n1165), .Y(n1168) );
  INVXL U162 ( .A(n1012), .Y(n70) );
  NAND2XL U163 ( .A(n1011), .B(n1012), .Y(n68) );
  ADDFHX2 U164 ( .A(n889), .B(n888), .CI(n887), .CO(n892), .S(n933) );
  ADDFHX2 U165 ( .A(n703), .B(n702), .CI(n701), .CO(n706), .S(n745) );
  NAND2XL U166 ( .A(n847), .B(n846), .Y(n36) );
  ADDFHX2 U167 ( .A(n918), .B(n917), .CI(n916), .CO(n935), .S(n983) );
  XNOR2XL U168 ( .A(n1138), .B(A[25]), .Y(n1159) );
  NAND2BXL U169 ( .AN(n122), .B(n81), .Y(n80) );
  XNOR2X1 U170 ( .A(n308), .B(n52), .Y(n481) );
  XOR2X1 U171 ( .A(n44), .B(n299), .Y(PRODUCT[35]) );
  NAND2XL U172 ( .A(n40), .B(n38), .Y(n1181) );
  AND2XL U173 ( .A(n1223), .B(n1222), .Y(n1334) );
  NAND2XL U174 ( .A(n1204), .B(n43), .Y(n40) );
  INVXL U175 ( .A(n117), .Y(n78) );
  AOI21XL U176 ( .A0(n338), .A1(n1173), .B0(n45), .Y(n44) );
  OR2XL U177 ( .A(n1221), .B(n1220), .Y(n1223) );
  NAND2XL U178 ( .A(n46), .B(n1267), .Y(n45) );
  OAI2BB1XL U179 ( .A0N(n968), .A1N(n970), .B0(n418), .Y(n477) );
  XOR2X1 U180 ( .A(n562), .B(n561), .Y(PRODUCT[28]) );
  NAND2X1 U181 ( .A(n108), .B(n134), .Y(n921) );
  INVXL U182 ( .A(n1210), .Y(n38) );
  XOR2X1 U183 ( .A(n941), .B(n940), .Y(PRODUCT[18]) );
  CLKINVX3 U184 ( .A(n26), .Y(n27) );
  OR2XL U185 ( .A(n1239), .B(n1245), .Y(n1249) );
  NAND2BX1 U186 ( .AN(n553), .B(n672), .Y(n20) );
  INVXL U187 ( .A(n1246), .Y(n39) );
  XOR2X1 U188 ( .A(n33), .B(n31), .Y(PRODUCT[15]) );
  INVXL U189 ( .A(A[11]), .Y(n99) );
  NAND2BXL U190 ( .AN(n1266), .B(n1175), .Y(n1178) );
  AND2X2 U191 ( .A(n856), .B(n1293), .Y(n857) );
  NAND2XL U192 ( .A(n672), .B(n1285), .Y(n673) );
  AND2X2 U193 ( .A(n560), .B(n1279), .Y(n561) );
  INVXL U194 ( .A(A[12]), .Y(n91) );
  INVXL U195 ( .A(A[8]), .Y(n35) );
  INVXL U196 ( .A(A[24]), .Y(n59) );
  INVXL U197 ( .A(A[23]), .Y(n54) );
  INVXL U198 ( .A(n1266), .Y(n1173) );
  INVX1 U199 ( .A(n1284), .Y(n672) );
  INVXL U200 ( .A(A[19]), .Y(n56) );
  INVXL U201 ( .A(A[18]), .Y(n53) );
  INVXL U202 ( .A(A[22]), .Y(n55) );
  INVXL U203 ( .A(A[21]), .Y(n58) );
  INVXL U204 ( .A(A[20]), .Y(n57) );
  NOR2X1 U205 ( .A(n1284), .B(n1282), .Y(n552) );
  NAND2X2 U206 ( .A(n12), .B(n11), .Y(n554) );
  AOI21X4 U207 ( .A0(n854), .A1(n17), .B0(n16), .Y(n11) );
  INVX4 U208 ( .A(n13), .Y(n15) );
  OAI21X4 U209 ( .A0(n1307), .A1(n1300), .B0(n1301), .Y(n13) );
  NAND2X4 U210 ( .A(n15), .B(n14), .Y(n21) );
  NAND3BX4 U211 ( .AN(n1300), .B(n18), .C(n1308), .Y(n14) );
  OAI21X2 U212 ( .A0(n1292), .A1(n1295), .B0(n1293), .Y(n16) );
  NOR2X2 U213 ( .A(n1292), .B(n1294), .Y(n17) );
  OAI21X2 U214 ( .A0(n1299), .A1(n1296), .B0(n1297), .Y(n854) );
  CLKINVX3 U215 ( .A(n1302), .Y(n18) );
  INVX1 U216 ( .A(n553), .Y(n669) );
  CLKINVX3 U217 ( .A(n554), .Y(n1086) );
  AOI21X1 U218 ( .A0(n21), .A1(n987), .B0(n938), .Y(n941) );
  XOR2X1 U219 ( .A(n853), .B(n988), .Y(PRODUCT[17]) );
  NAND2X2 U220 ( .A(n296), .B(n22), .Y(n47) );
  AOI22X2 U221 ( .A0(n24), .A1(n554), .B0(n670), .B1(n23), .Y(n22) );
  NAND2BX2 U222 ( .AN(n100), .B(n42), .Y(n670) );
  NOR2X1 U223 ( .A(n25), .B(n553), .Y(n24) );
  NAND2X1 U224 ( .A(n295), .B(n552), .Y(n25) );
  AOI21X2 U225 ( .A0(n27), .A1(n855), .B0(n854), .Y(n897) );
  NOR2X1 U226 ( .A(n1298), .B(n1296), .Y(n855) );
  OAI21XL U227 ( .A0(n897), .A1(n1294), .B0(n1295), .Y(n30) );
  OAI22X1 U228 ( .A0(n1135), .A1(n638), .B0(n954), .B1(n601), .Y(n639) );
  NAND2X1 U229 ( .A(n708), .B(n707), .Y(mult_x_1_n234) );
  BUFX8 U230 ( .A(n307), .Y(n966) );
  XNOR2X1 U231 ( .A(n1138), .B(A[7]), .Y(n720) );
  XNOR2X4 U232 ( .A(B[14]), .B(B[13]), .Y(n48) );
  OAI22X1 U233 ( .A0(n768), .A1(n964), .B0(n966), .B1(n34), .Y(n801) );
  OAI22X1 U234 ( .A0(n832), .A1(n966), .B0(n964), .B1(n34), .Y(n870) );
  XOR2X1 U235 ( .A(n922), .B(n35), .Y(n34) );
  OAI2BB1X1 U236 ( .A0N(n37), .A1N(n845), .B0(n36), .Y(n850) );
  OR2X2 U237 ( .A(n847), .B(n846), .Y(n37) );
  XOR3X2 U238 ( .A(n846), .B(n847), .C(n845), .Y(n890) );
  OAI2BB1X1 U239 ( .A0N(n1238), .A1N(n39), .B0(n1179), .Y(n1210) );
  NAND2X1 U240 ( .A(n1311), .B(n1310), .Y(n752) );
  AOI21X1 U241 ( .A0(n670), .A1(n672), .B0(n630), .Y(n41) );
  NAND2X1 U242 ( .A(n710), .B(n71), .Y(n42) );
  NAND2X1 U243 ( .A(n750), .B(n71), .Y(n553) );
  NOR2X1 U244 ( .A(n709), .B(n1286), .Y(n71) );
  NOR2X1 U245 ( .A(n1310), .B(n1311), .Y(n709) );
  NOR2X1 U246 ( .A(n1290), .B(n1288), .Y(n750) );
  NOR2BX1 U247 ( .AN(n1238), .B(n1239), .Y(n1204) );
  NOR2X1 U248 ( .A(n1239), .B(n1268), .Y(n337) );
  OAI21XL U249 ( .A0(n1246), .A1(n1268), .B0(n1269), .Y(n338) );
  OAI21XL U250 ( .A0(n1282), .A1(n1285), .B0(n1283), .Y(n555) );
  OAI21XL U251 ( .A0(n1250), .A1(n1239), .B0(n1246), .Y(n368) );
  OAI22X1 U252 ( .A0(n907), .A1(n8), .B0(n306), .B1(n1161), .Y(n949) );
  NAND2X4 U253 ( .A(n48), .B(n49), .Y(n1161) );
  XOR2X2 U254 ( .A(B[14]), .B(B[15]), .Y(n49) );
  XNOR2X1 U255 ( .A(n308), .B(n50), .Y(n521) );
  INVX1 U256 ( .A(A[15]), .Y(n50) );
  XNOR2X1 U257 ( .A(n308), .B(n53), .Y(n424) );
  XNOR2X1 U258 ( .A(n308), .B(n55), .Y(n343) );
  XNOR2X1 U259 ( .A(n308), .B(n56), .Y(n388) );
  XNOR2X1 U260 ( .A(n308), .B(n57), .Y(n381) );
  XNOR2X1 U261 ( .A(n308), .B(n58), .Y(n348) );
  XNOR2X1 U262 ( .A(n308), .B(n59), .Y(n326) );
  OAI2BB1X1 U263 ( .A0N(n61), .A1N(n563), .B0(n60), .Y(n551) );
  NOR2XL U264 ( .A(n564), .B(n565), .Y(n62) );
  XNOR3X2 U265 ( .A(n63), .B(n564), .C(n563), .Y(n588) );
  NOR2X1 U266 ( .A(n192), .B(n191), .Y(n64) );
  XOR2X1 U267 ( .A(B[6]), .B(B[7]), .Y(n103) );
  OAI22X1 U268 ( .A0(n1100), .A1(n569), .B0(n1101), .B1(n521), .Y(n574) );
  OAI22X1 U269 ( .A0(n7), .A1(n758), .B0(n8), .B1(n720), .Y(n761) );
  OAI22X1 U270 ( .A0(n7), .A1(n536), .B0(n8), .B1(n483), .Y(n519) );
  XNOR2X1 U271 ( .A(n1138), .B(A[5]), .Y(n787) );
  XNOR2X1 U272 ( .A(n1138), .B(A[6]), .Y(n758) );
  OAI22X2 U273 ( .A0(n7), .A1(n720), .B0(n8), .B1(n679), .Y(n723) );
  NAND2X1 U274 ( .A(n107), .B(n113), .Y(n835) );
  OAI21XL U275 ( .A0(n1274), .A1(n1277), .B0(n1275), .Y(n440) );
  XNOR2XL U276 ( .A(n905), .B(A[9]), .Y(n198) );
  INVXL U277 ( .A(n1243), .Y(n1179) );
  INVXL U278 ( .A(n1237), .Y(n1209) );
  NOR2XL U279 ( .A(n1178), .B(n1268), .Y(n1238) );
  NOR2XL U280 ( .A(n1237), .B(n1256), .Y(n1242) );
  INVXL U281 ( .A(n1262), .Y(n1183) );
  XNOR2XL U282 ( .A(n1127), .B(A[19]), .Y(n312) );
  XNOR2X1 U283 ( .A(n908), .B(A[5]), .Y(n961) );
  NAND2BXL U284 ( .AN(A[0]), .B(n908), .Y(n168) );
  OAI22XL U285 ( .A0(n240), .A1(n170), .B0(n198), .B1(n1085), .Y(n196) );
  XNOR2XL U286 ( .A(n908), .B(A[24]), .Y(n315) );
  XNOR2XL U287 ( .A(n908), .B(A[23]), .Y(n345) );
  XNOR2XL U288 ( .A(n1120), .B(A[19]), .Y(n344) );
  XNOR2XL U289 ( .A(n1127), .B(A[16]), .Y(n379) );
  XNOR2XL U290 ( .A(n908), .B(A[22]), .Y(n380) );
  XNOR2XL U291 ( .A(n1120), .B(A[18]), .Y(n382) );
  XNOR2X2 U292 ( .A(B[8]), .B(B[7]), .Y(n685) );
  XNOR2XL U293 ( .A(n905), .B(A[5]), .Y(n112) );
  XNOR2XL U294 ( .A(n905), .B(A[6]), .Y(n106) );
  XNOR2XL U295 ( .A(n905), .B(A[8]), .Y(n170) );
  NAND2X1 U296 ( .A(n103), .B(n105), .Y(n979) );
  NAND2XL U297 ( .A(n1238), .B(n1242), .Y(n1245) );
  NAND2XL U298 ( .A(n366), .B(n1269), .Y(n367) );
  XNOR2X1 U299 ( .A(n408), .B(n407), .Y(PRODUCT[32]) );
  NAND2XL U300 ( .A(n406), .B(n1271), .Y(n407) );
  OAI21XL U301 ( .A0(n1250), .A1(n405), .B0(n404), .Y(n408) );
  XNOR2XL U302 ( .A(n1120), .B(A[21]), .Y(n313) );
  XNOR2XL U303 ( .A(n1120), .B(A[22]), .Y(n327) );
  XNOR2XL U304 ( .A(n1127), .B(A[21]), .Y(n1103) );
  XNOR2XL U305 ( .A(n1127), .B(A[22]), .Y(n1118) );
  BUFX3 U306 ( .A(n212), .Y(n1101) );
  NAND2BXL U307 ( .AN(A[0]), .B(n1138), .Y(n907) );
  OAI22XL U308 ( .A0(n240), .A1(n952), .B0(n951), .B1(n1085), .Y(n1002) );
  OAI22XL U309 ( .A0(n1135), .A1(n955), .B0(n954), .B1(n953), .Y(n1001) );
  XNOR2XL U310 ( .A(n905), .B(A[4]), .Y(n139) );
  XNOR2XL U311 ( .A(n1127), .B(A[24]), .Y(n1139) );
  OAI2BB1XL U312 ( .A0N(n1136), .A1N(n1135), .B0(n1134), .Y(n1140) );
  NOR2XL U313 ( .A(n1158), .B(n1132), .Y(n1141) );
  INVXL U314 ( .A(n1133), .Y(n1134) );
  XNOR2XL U315 ( .A(n1127), .B(A[23]), .Y(n1128) );
  NAND3X1 U316 ( .A(n86), .B(n1075), .C(n95), .Y(n289) );
  OAI22XL U317 ( .A0(n970), .A1(n141), .B0(n968), .B1(n121), .Y(n150) );
  ADDFX2 U318 ( .A(n120), .B(n67), .CI(n118), .CO(n158), .S(n157) );
  OAI22XL U319 ( .A0(n970), .A1(n121), .B0(n968), .B1(n111), .Y(n120) );
  XOR2XL U320 ( .A(n82), .B(n79), .Y(n118) );
  OAI22XL U321 ( .A0(n1161), .A1(n1139), .B0(n8), .B1(n1159), .Y(n1164) );
  INVXL U322 ( .A(n1224), .Y(n147) );
  NOR2XL U323 ( .A(n155), .B(n154), .Y(n1232) );
  NAND2XL U324 ( .A(n155), .B(n154), .Y(n1233) );
  NOR2X1 U325 ( .A(n157), .B(n156), .Y(n1199) );
  NAND2XL U326 ( .A(n159), .B(n158), .Y(n1191) );
  INVXL U327 ( .A(n1267), .Y(n1176) );
  XNOR2XL U328 ( .A(n905), .B(A[17]), .Y(n830) );
  XNOR2XL U329 ( .A(n905), .B(A[25]), .Y(n517) );
  XNOR2XL U330 ( .A(n919), .B(A[22]), .Y(n570) );
  NOR2XL U331 ( .A(n1276), .B(n1274), .Y(n439) );
  INVXL U332 ( .A(n1264), .Y(n1175) );
  NAND2XL U333 ( .A(n669), .B(n552), .Y(n592) );
  INVXL U334 ( .A(n1280), .Y(n593) );
  INVXL U335 ( .A(n1263), .Y(n1182) );
  NAND2XL U336 ( .A(n1204), .B(n1183), .Y(n1185) );
  INVXL U337 ( .A(n1260), .Y(n1186) );
  INVX1 U338 ( .A(n1298), .Y(n987) );
  XNOR2X1 U339 ( .A(n924), .B(A[3]), .Y(n207) );
  XNOR2XL U340 ( .A(n919), .B(A[8]), .Y(n214) );
  XNOR2XL U341 ( .A(n919), .B(A[9]), .Y(n243) );
  XNOR2XL U342 ( .A(n924), .B(A[5]), .Y(n242) );
  NAND2BXL U343 ( .AN(A[0]), .B(n1120), .Y(n236) );
  XNOR2XL U344 ( .A(n905), .B(A[12]), .Y(n238) );
  XNOR2XL U345 ( .A(n919), .B(A[10]), .Y(n248) );
  XNOR2XL U346 ( .A(n908), .B(A[17]), .Y(n527) );
  XNOR2X1 U347 ( .A(n924), .B(A[21]), .Y(n458) );
  XNOR2XL U348 ( .A(n1120), .B(A[6]), .Y(n823) );
  XNOR2XL U349 ( .A(n905), .B(A[13]), .Y(n952) );
  XNOR2X1 U350 ( .A(n1120), .B(A[1]), .Y(n955) );
  XNOR2XL U351 ( .A(n1120), .B(A[0]), .Y(n246) );
  XNOR2XL U352 ( .A(n924), .B(A[7]), .Y(n978) );
  XNOR2XL U353 ( .A(n908), .B(A[4]), .Y(n250) );
  XNOR2XL U354 ( .A(n908), .B(A[3]), .Y(n251) );
  XNOR2XL U355 ( .A(n650), .B(A[6]), .Y(n208) );
  NAND2BXL U356 ( .AN(A[0]), .B(n922), .Y(n194) );
  OAI22XL U357 ( .A0(n240), .A1(n198), .B0(n197), .B1(n1085), .Y(n205) );
  NOR2BXL U358 ( .AN(A[0]), .B(n212), .Y(n206) );
  XNOR2XL U359 ( .A(n905), .B(A[21]), .Y(n688) );
  XNOR2X1 U360 ( .A(n922), .B(A[13]), .Y(n610) );
  XNOR2XL U361 ( .A(n919), .B(A[21]), .Y(n611) );
  XNOR2XL U362 ( .A(n905), .B(A[20]), .Y(n728) );
  XNOR2XL U363 ( .A(n905), .B(A[18]), .Y(n795) );
  XNOR2XL U364 ( .A(n905), .B(A[19]), .Y(n766) );
  XNOR2XL U365 ( .A(n650), .B(n904), .Y(n822) );
  XNOR2XL U366 ( .A(n919), .B(A[17]), .Y(n769) );
  XNOR2XL U367 ( .A(n919), .B(A[18]), .Y(n731) );
  XNOR2XL U368 ( .A(n919), .B(A[19]), .Y(n690) );
  XNOR2XL U369 ( .A(n919), .B(A[20]), .Y(n649) );
  XNOR2XL U370 ( .A(n919), .B(A[24]), .Y(n488) );
  INVXL U371 ( .A(n517), .Y(n490) );
  XNOR2XL U372 ( .A(n1156), .B(n904), .Y(n369) );
  XNOR2XL U373 ( .A(n1127), .B(A[15]), .Y(n387) );
  XNOR2XL U374 ( .A(n1120), .B(n904), .Y(n512) );
  OAI22XL U375 ( .A0(n926), .A1(n535), .B0(n757), .B1(n482), .Y(n520) );
  XNOR2XL U376 ( .A(n908), .B(A[18]), .Y(n516) );
  XNOR2XL U377 ( .A(n919), .B(A[25]), .Y(n417) );
  OAI22X1 U378 ( .A0(n970), .A1(n488), .B0(n968), .B1(n417), .Y(n478) );
  CMPR32X1 U379 ( .A(n427), .B(n426), .C(n425), .CO(n412), .S(n468) );
  INVXL U380 ( .A(n390), .Y(n425) );
  OAI22XL U381 ( .A0(n1135), .A1(n423), .B0(n1136), .B1(n383), .Y(n427) );
  XNOR2XL U382 ( .A(B[9]), .B(A[21]), .Y(n415) );
  NAND2BXL U383 ( .AN(A[0]), .B(n650), .Y(n114) );
  XNOR2XL U384 ( .A(n919), .B(A[5]), .Y(n162) );
  XNOR2XL U385 ( .A(n905), .B(A[7]), .Y(n171) );
  NAND2XL U386 ( .A(n1204), .B(n1209), .Y(n1212) );
  INVXL U387 ( .A(n1240), .Y(n1208) );
  INVXL U388 ( .A(n1256), .Y(n1213) );
  AOI21XL U389 ( .A0(n1243), .A1(n1242), .B0(n1241), .Y(n1244) );
  INVXL U390 ( .A(n1276), .Y(n508) );
  NAND2XL U391 ( .A(n1183), .B(n1263), .Y(n1180) );
  NAND2XL U392 ( .A(n1206), .B(n1259), .Y(n1197) );
  XOR2X1 U393 ( .A(n1062), .B(n1304), .Y(PRODUCT[14]) );
  INVXL U394 ( .A(n1294), .Y(n895) );
  XOR2X1 U395 ( .A(n1086), .B(n817), .Y(PRODUCT[21]) );
  ADDFX2 U396 ( .A(n203), .B(n202), .CI(n201), .CO(n221), .S(n229) );
  OAI22XL U397 ( .A0(n835), .A1(n163), .B0(n9), .B1(n209), .Y(n201) );
  OAI22X1 U398 ( .A0(n962), .A1(n161), .B0(n960), .B1(n200), .Y(n202) );
  OAI22XL U399 ( .A0(n926), .A1(n172), .B0(n757), .B1(n207), .Y(n203) );
  OAI22XL U400 ( .A0(n921), .A1(n167), .B0(n968), .B1(n210), .Y(n220) );
  XOR2XL U401 ( .A(n195), .B(n196), .Y(n219) );
  XNOR2XL U402 ( .A(n1120), .B(A[20]), .Y(n317) );
  OAI2BB1XL U403 ( .A0N(n685), .A1N(n643), .B0(n311), .Y(n328) );
  INVXL U404 ( .A(n310), .Y(n311) );
  OAI22XL U405 ( .A0(n1100), .A1(n314), .B0(n1101), .B1(n326), .Y(n331) );
  OAI22XL U406 ( .A0(n1135), .A1(n313), .B0(n1136), .B1(n327), .Y(n332) );
  XNOR2XL U407 ( .A(n1120), .B(A[23]), .Y(n1102) );
  XNOR2XL U408 ( .A(n1156), .B(A[20]), .Y(n1097) );
  OAI22X1 U409 ( .A0(n966), .A1(n879), .B0(n964), .B1(n832), .Y(n878) );
  OAI22XL U410 ( .A0(n7), .A1(n872), .B0(n8), .B1(n861), .Y(n883) );
  OAI22XL U411 ( .A0(n1135), .A1(n912), .B0(n954), .B1(n875), .Y(n927) );
  OAI22X1 U412 ( .A0(n962), .A1(n909), .B0(n960), .B1(n873), .Y(n929) );
  ADDFX2 U413 ( .A(n932), .B(n931), .CI(n930), .CO(n947), .S(n992) );
  OAI22X1 U414 ( .A0(n948), .A1(n976), .B0(n9), .B1(n90), .Y(n932) );
  OAI22X1 U415 ( .A0(n966), .A1(n923), .B0(n964), .B1(n879), .Y(n931) );
  ADDFX2 U416 ( .A(n915), .B(n914), .CI(n913), .CO(n918), .S(n956) );
  OAI22XL U417 ( .A0(n240), .A1(n906), .B0(n871), .B1(n1085), .Y(n914) );
  NOR2BXL U418 ( .AN(A[0]), .B(n384), .Y(n915) );
  OAI22XL U419 ( .A0(n7), .A1(n910), .B0(n8), .B1(n872), .Y(n913) );
  OAI22X1 U420 ( .A0(n962), .A1(n959), .B0(n960), .B1(n909), .Y(n973) );
  OAI22X1 U421 ( .A0(n7), .A1(n911), .B0(n8), .B1(n910), .Y(n972) );
  OAI22XL U422 ( .A0(n970), .A1(n969), .B0(n968), .B1(n967), .Y(n1007) );
  OAI22XL U423 ( .A0(n962), .A1(n961), .B0(n960), .B1(n959), .Y(n1009) );
  OAI2BB1XL U424 ( .A0N(n757), .A1N(n926), .B0(n305), .Y(n352) );
  NOR2XL U425 ( .A(n1158), .B(n302), .Y(n354) );
  OAI22XL U426 ( .A0(n1100), .A1(n381), .B0(n1101), .B1(n348), .Y(n372) );
  OAI22XL U427 ( .A0(n7), .A1(n379), .B0(n8), .B1(n347), .Y(n373) );
  ADDFX2 U428 ( .A(n377), .B(n376), .CI(n375), .CO(n356), .S(n409) );
  OAI22XL U429 ( .A0(n962), .A1(n380), .B0(n960), .B1(n345), .Y(n376) );
  OAI22XL U430 ( .A0(n1135), .A1(n382), .B0(n1136), .B1(n344), .Y(n377) );
  XNOR2XL U431 ( .A(n919), .B(A[4]), .Y(n111) );
  ADDFX2 U432 ( .A(n229), .B(n228), .CI(n227), .CO(n230), .S(n192) );
  INVXL U433 ( .A(n1142), .Y(n1129) );
  INVXL U434 ( .A(n1116), .Y(n1104) );
  OAI22XL U435 ( .A0(n1161), .A1(n324), .B0(n8), .B1(n1103), .Y(n1106) );
  OAI22XL U436 ( .A0(n976), .A1(n974), .B0(n9), .B1(n948), .Y(n1000) );
  XNOR2XL U437 ( .A(n905), .B(A[1]), .Y(n126) );
  OAI22XL U438 ( .A0(n970), .A1(n136), .B0(n968), .B1(n135), .Y(n137) );
  INVXL U439 ( .A(n919), .Y(n136) );
  NAND2BXL U440 ( .AN(A[0]), .B(n919), .Y(n135) );
  XNOR2XL U441 ( .A(n919), .B(A[0]), .Y(n133) );
  OAI22XL U442 ( .A0(n240), .A1(n140), .B0(n139), .B1(n1085), .Y(n152) );
  NOR2BXL U443 ( .AN(A[0]), .B(n9), .Y(n153) );
  OAI21XL U444 ( .A0(n970), .A1(n93), .B0(n92), .Y(n151) );
  OAI21XL U445 ( .A0(n78), .A1(n77), .B0(n76), .Y(n187) );
  INVXL U446 ( .A(n116), .Y(n77) );
  OAI2BB1XL U447 ( .A0N(n8), .A1N(n1161), .B0(n1160), .Y(n1162) );
  INVXL U448 ( .A(n1159), .Y(n1160) );
  NOR2XL U449 ( .A(n1158), .B(n1157), .Y(n1163) );
  XNOR2XL U450 ( .A(n1156), .B(A[24]), .Y(n1157) );
  NOR2XL U451 ( .A(n1158), .B(n1137), .Y(n1155) );
  INVXL U452 ( .A(n1164), .Y(n1154) );
  XNOR2XL U453 ( .A(n1156), .B(A[23]), .Y(n1137) );
  OAI22XL U454 ( .A0(n240), .A1(A[0]), .B0(n126), .B1(n1085), .Y(n1221) );
  NAND2XL U455 ( .A(n128), .B(n240), .Y(n1220) );
  NAND2BXL U456 ( .AN(A[0]), .B(n905), .Y(n128) );
  NAND2XL U457 ( .A(n1221), .B(n1220), .Y(n1222) );
  INVXL U458 ( .A(n1222), .Y(n1218) );
  NOR2XL U459 ( .A(n138), .B(n137), .Y(n1227) );
  NAND2XL U460 ( .A(n138), .B(n137), .Y(n1228) );
  AOI21XL U461 ( .A0(n1217), .A1(n1218), .B0(n131), .Y(n1230) );
  INVXL U462 ( .A(n1216), .Y(n131) );
  NAND2XL U463 ( .A(n146), .B(n145), .Y(n1224) );
  OAI21XL U464 ( .A0(n1227), .A1(n1230), .B0(n1228), .Y(n1225) );
  INVXL U465 ( .A(n1189), .Y(n1201) );
  NAND3X2 U466 ( .A(n84), .B(n83), .C(n1191), .Y(n1172) );
  OR2X2 U467 ( .A(n1190), .B(n1200), .Y(n83) );
  NAND2XL U468 ( .A(n1203), .B(n1206), .Y(n1237) );
  INVXL U469 ( .A(n1285), .Y(n630) );
  NOR2XL U470 ( .A(n1262), .B(n1260), .Y(n1203) );
  XNOR2XL U471 ( .A(n905), .B(A[10]), .Y(n197) );
  XNOR2XL U472 ( .A(n905), .B(A[24]), .Y(n530) );
  XNOR2XL U473 ( .A(n905), .B(A[23]), .Y(n608) );
  XNOR2XL U474 ( .A(n905), .B(A[22]), .Y(n646) );
  AOI21XL U475 ( .A0(n1176), .A1(n1175), .B0(n1174), .Y(n1177) );
  INVXL U476 ( .A(n1265), .Y(n1174) );
  AOI21XL U477 ( .A0(n1207), .A1(n1206), .B0(n1205), .Y(n1240) );
  INVXL U478 ( .A(n1259), .Y(n1205) );
  INVX1 U479 ( .A(n670), .Y(n671) );
  AOI21XL U480 ( .A0(n710), .A1(n753), .B0(n712), .Y(n713) );
  INVXL U481 ( .A(n1268), .Y(n366) );
  INVXL U482 ( .A(n1273), .Y(n403) );
  NAND2XL U483 ( .A(n439), .B(n443), .Y(n405) );
  INVXL U484 ( .A(n1282), .Y(n631) );
  NAND2XL U485 ( .A(n557), .B(n669), .Y(n559) );
  AOI21XL U486 ( .A0(n670), .A1(n557), .B0(n556), .Y(n558) );
  INVXL U487 ( .A(n555), .Y(n590) );
  INVXL U488 ( .A(n1278), .Y(n560) );
  INVXL U489 ( .A(n439), .Y(n442) );
  INVXL U490 ( .A(n440), .Y(n441) );
  INVXL U491 ( .A(n1272), .Y(n443) );
  NAND2XL U492 ( .A(n1204), .B(n1203), .Y(n1196) );
  INVXL U493 ( .A(n1258), .Y(n1206) );
  INVXL U494 ( .A(n1299), .Y(n938) );
  INVXL U495 ( .A(n710), .Y(n711) );
  INVX1 U496 ( .A(n709), .Y(n753) );
  XNOR2XL U497 ( .A(n905), .B(A[11]), .Y(n239) );
  XNOR2XL U498 ( .A(n1156), .B(A[18]), .Y(n309) );
  XNOR2XL U499 ( .A(n1156), .B(A[10]), .Y(n511) );
  XNOR2XL U500 ( .A(n650), .B(A[21]), .Y(n523) );
  XNOR2X1 U501 ( .A(n922), .B(A[7]), .Y(n832) );
  XNOR2XL U502 ( .A(n919), .B(A[15]), .Y(n833) );
  XNOR2XL U503 ( .A(n1120), .B(A[5]), .Y(n863) );
  XNOR2X1 U504 ( .A(n1138), .B(A[3]), .Y(n861) );
  OAI22XL U505 ( .A0(n240), .A1(n871), .B0(n830), .B1(n1085), .Y(n867) );
  NOR2XL U506 ( .A(n1158), .B(n831), .Y(n866) );
  NAND2BXL U507 ( .AN(A[0]), .B(n1156), .Y(n831) );
  XNOR2X1 U508 ( .A(n908), .B(A[8]), .Y(n873) );
  XNOR2XL U509 ( .A(n1120), .B(A[4]), .Y(n875) );
  XNOR2XL U510 ( .A(n919), .B(n904), .Y(n874) );
  XNOR2XL U511 ( .A(n905), .B(A[16]), .Y(n871) );
  XNOR2XL U512 ( .A(n905), .B(A[15]), .Y(n906) );
  XNOR2XL U513 ( .A(n905), .B(n904), .Y(n951) );
  XNOR2X1 U514 ( .A(n1120), .B(A[3]), .Y(n912) );
  XNOR2X1 U515 ( .A(n1120), .B(A[2]), .Y(n953) );
  XNOR2XL U516 ( .A(n908), .B(A[6]), .Y(n959) );
  XNOR2XL U517 ( .A(n919), .B(A[13]), .Y(n920) );
  XNOR2XL U518 ( .A(n922), .B(A[5]), .Y(n923) );
  XNOR2XL U519 ( .A(n922), .B(A[4]), .Y(n963) );
  XNOR2XL U520 ( .A(n919), .B(A[12]), .Y(n967) );
  XNOR2XL U521 ( .A(n908), .B(A[15]), .Y(n642) );
  CMPR32X1 U522 ( .A(n577), .B(n576), .C(n575), .CO(n578), .S(n622) );
  OAI22XL U523 ( .A0(n962), .A1(n605), .B0(n685), .B1(n527), .Y(n577) );
  ADDFX2 U524 ( .A(n574), .B(n573), .CI(n572), .CO(n580), .S(n623) );
  OAI22XL U525 ( .A0(n976), .A1(n571), .B0(n9), .B1(n523), .Y(n572) );
  OAI22X1 U526 ( .A0(n970), .A1(n570), .B0(n968), .B1(n522), .Y(n573) );
  XNOR2X1 U527 ( .A(n924), .B(A[17]), .Y(n636) );
  ADDFX2 U528 ( .A(n615), .B(n614), .CI(n613), .CO(n624), .S(n662) );
  OAI22XL U529 ( .A0(n976), .A1(n612), .B0(n9), .B1(n571), .Y(n613) );
  OAI22X1 U530 ( .A0(n970), .A1(n611), .B0(n968), .B1(n570), .Y(n614) );
  XNOR2XL U531 ( .A(n1156), .B(A[16]), .Y(n302) );
  XNOR2XL U532 ( .A(n1156), .B(A[15]), .Y(n346) );
  XNOR2XL U533 ( .A(n1138), .B(n904), .Y(n420) );
  XNOR2XL U534 ( .A(n908), .B(A[20]), .Y(n422) );
  XNOR2XL U535 ( .A(n919), .B(A[6]), .Y(n167) );
  XNOR2XL U536 ( .A(n650), .B(A[4]), .Y(n163) );
  NAND2XL U537 ( .A(n1173), .B(n1267), .Y(n341) );
  NAND2XL U538 ( .A(n1175), .B(n1265), .Y(n299) );
  XNOR2X1 U539 ( .A(n595), .B(n594), .Y(PRODUCT[27]) );
  NAND2XL U540 ( .A(n593), .B(n1281), .Y(n594) );
  OAI21XL U541 ( .A0(n1086), .A1(n592), .B0(n591), .Y(n595) );
  NAND2XL U542 ( .A(n1186), .B(n1261), .Y(n1187) );
  NAND2XL U543 ( .A(n1087), .B(n1289), .Y(n1088) );
  OAI22XL U544 ( .A0(n970), .A1(n210), .B0(n968), .B1(n214), .Y(n215) );
  OAI22XL U545 ( .A0(n926), .A1(n207), .B0(n757), .B1(n211), .Y(n217) );
  OAI22XL U546 ( .A0(n970), .A1(n214), .B0(n968), .B1(n243), .Y(n257) );
  OAI22XL U547 ( .A0(n979), .A1(n211), .B0(n757), .B1(n242), .Y(n259) );
  OAI22XL U548 ( .A0(n976), .A1(n244), .B0(n9), .B1(n249), .Y(n263) );
  OAI22XL U549 ( .A0(n926), .A1(n242), .B0(n757), .B1(n245), .Y(n265) );
  OAI22XL U550 ( .A0(n970), .A1(n243), .B0(n968), .B1(n248), .Y(n264) );
  OAI22XL U551 ( .A0(n240), .A1(n238), .B0(n952), .B1(n1085), .Y(n981) );
  OAI22XL U552 ( .A0(n1135), .A1(n300), .B0(n1136), .B1(n236), .Y(n980) );
  INVXL U553 ( .A(n1120), .Y(n300) );
  OAI22XL U554 ( .A0(n976), .A1(n249), .B0(n9), .B1(n975), .Y(n1004) );
  OAI22X1 U555 ( .A0(n962), .A1(n250), .B0(n960), .B1(n961), .Y(n1006) );
  OAI22XL U556 ( .A0(n921), .A1(n248), .B0(n968), .B1(n969), .Y(n1005) );
  XNOR2XL U557 ( .A(n1120), .B(A[25]), .Y(n1133) );
  XNOR2XL U558 ( .A(n1156), .B(A[22]), .Y(n1132) );
  XNOR2XL U559 ( .A(n1156), .B(A[21]), .Y(n1119) );
  XNOR2XL U560 ( .A(n1127), .B(A[20]), .Y(n324) );
  XNOR2XL U561 ( .A(n1156), .B(A[19]), .Y(n325) );
  INVXL U562 ( .A(n329), .Y(n318) );
  OAI22XL U563 ( .A0(n962), .A1(n527), .B0(n685), .B1(n516), .Y(n543) );
  CMPR32X1 U564 ( .A(n540), .B(n539), .C(n538), .CO(n534), .S(n582) );
  OAI22XL U565 ( .A0(n1135), .A1(n537), .B0(n1136), .B1(n512), .Y(n538) );
  OAI22XL U566 ( .A0(n976), .A1(n523), .B0(n9), .B1(n510), .Y(n540) );
  NOR2XL U567 ( .A(n1158), .B(n511), .Y(n539) );
  CMPR32X1 U568 ( .A(n515), .B(n514), .C(n513), .CO(n499), .S(n533) );
  NOR2XL U569 ( .A(n384), .B(n459), .Y(n514) );
  OAI22X1 U570 ( .A0(n926), .A1(n482), .B0(n757), .B1(n458), .Y(n515) );
  ADDFX2 U571 ( .A(n826), .B(n825), .CI(n824), .CO(n807), .S(n843) );
  OAI22X1 U572 ( .A0(n7), .A1(n797), .B0(n8), .B1(n787), .Y(n825) );
  OAI22XL U573 ( .A0(n926), .A1(n827), .B0(n757), .B1(n786), .Y(n826) );
  OAI22XL U574 ( .A0(n966), .A1(n247), .B0(n964), .B1(n965), .Y(n1024) );
  OAI22XL U575 ( .A0(n962), .A1(n251), .B0(n960), .B1(n250), .Y(n268) );
  OAI22XL U576 ( .A0(n127), .A1(n728), .B0(n688), .B1(n1085), .Y(n727) );
  XNOR2XL U577 ( .A(n1120), .B(A[10]), .Y(n680) );
  OAI22XL U578 ( .A0(n976), .A1(n651), .B0(n9), .B1(n612), .Y(n652) );
  XNOR2XL U579 ( .A(n924), .B(A[15]), .Y(n719) );
  XNOR2XL U580 ( .A(n1120), .B(A[9]), .Y(n721) );
  XNOR2XL U581 ( .A(n924), .B(n904), .Y(n756) );
  XNOR2XL U582 ( .A(n1120), .B(A[8]), .Y(n759) );
  XNOR2XL U583 ( .A(n1120), .B(A[7]), .Y(n788) );
  XNOR2XL U584 ( .A(n924), .B(A[13]), .Y(n786) );
  OAI22XL U585 ( .A0(n127), .A1(n795), .B0(n766), .B1(n1085), .Y(n794) );
  OAI22XL U586 ( .A0(n976), .A1(n822), .B0(n9), .B1(n770), .Y(n799) );
  OAI22XL U587 ( .A0(n976), .A1(n732), .B0(n9), .B1(n691), .Y(n733) );
  OAI22XL U588 ( .A0(n976), .A1(n691), .B0(n9), .B1(n651), .Y(n692) );
  ADDFX2 U589 ( .A(n526), .B(n525), .CI(n524), .CO(n568), .S(n579) );
  OAI2BB1XL U590 ( .A0N(n1085), .A1N(n240), .B0(n490), .Y(n524) );
  OAI22X1 U591 ( .A0(n970), .A1(n522), .B0(n968), .B1(n488), .Y(n525) );
  ADDFX2 U592 ( .A(n583), .B(n582), .CI(n581), .CO(n584), .S(n625) );
  OAI22XL U593 ( .A0(n1135), .A1(n344), .B0(n1136), .B1(n317), .Y(n349) );
  OAI22XL U594 ( .A0(n962), .A1(n345), .B0(n685), .B1(n315), .Y(n351) );
  OAI2BB1XL U595 ( .A0N(n9), .A1N(n976), .B0(n371), .Y(n389) );
  NOR2XL U596 ( .A(n1158), .B(n369), .Y(n391) );
  INVXL U597 ( .A(n370), .Y(n371) );
  OAI22XL U598 ( .A0(n962), .A1(n415), .B0(n685), .B1(n380), .Y(n392) );
  OAI22XL U599 ( .A0(n7), .A1(n387), .B0(n8), .B1(n379), .Y(n393) );
  OAI22XL U600 ( .A0(n1100), .A1(n388), .B0(n1101), .B1(n381), .Y(n414) );
  OAI22XL U601 ( .A0(n1135), .A1(n383), .B0(n1136), .B1(n382), .Y(n413) );
  CMPR32X1 U602 ( .A(n493), .B(n492), .C(n491), .CO(n502), .S(n567) );
  INVXL U603 ( .A(n478), .Y(n491) );
  OAI22XL U604 ( .A0(n1135), .A1(n512), .B0(n1136), .B1(n475), .Y(n493) );
  OAI22XL U605 ( .A0(n962), .A1(n516), .B0(n685), .B1(n480), .Y(n496) );
  OR2XL U606 ( .A(n520), .B(n519), .Y(n494) );
  ADDFX2 U607 ( .A(n479), .B(n478), .CI(n477), .CO(n456), .S(n501) );
  NOR2X1 U608 ( .A(n1158), .B(n416), .Y(n479) );
  INVXL U609 ( .A(n417), .Y(n418) );
  XNOR2XL U610 ( .A(n905), .B(A[2]), .Y(n132) );
  OR2X2 U611 ( .A(n141), .B(n968), .Y(n92) );
  XOR2XL U612 ( .A(n919), .B(n94), .Y(n93) );
  INVXL U613 ( .A(A[1]), .Y(n94) );
  XNOR2XL U614 ( .A(n919), .B(A[2]), .Y(n141) );
  OAI22XL U615 ( .A0(n240), .A1(n139), .B0(n112), .B1(n1085), .Y(n125) );
  INVXL U616 ( .A(n650), .Y(n115) );
  XOR2XL U617 ( .A(n117), .B(n116), .Y(n82) );
  XNOR2XL U618 ( .A(n919), .B(A[3]), .Y(n121) );
  OAI22X1 U619 ( .A0(n240), .A1(n112), .B0(n106), .B1(n1085), .Y(n116) );
  NAND2BXL U620 ( .AN(A[0]), .B(n924), .Y(n104) );
  ADDFX2 U621 ( .A(n179), .B(n178), .CI(n177), .CO(n184), .S(n186) );
  OAI22X1 U622 ( .A0(n926), .A1(n109), .B0(n757), .B1(n173), .Y(n178) );
  OAI22XL U623 ( .A0(n970), .A1(n111), .B0(n968), .B1(n162), .Y(n179) );
  ADDFX2 U624 ( .A(n182), .B(n181), .CI(n180), .CO(n228), .S(n183) );
  OAI22XL U625 ( .A0(n921), .A1(n162), .B0(n968), .B1(n167), .Y(n182) );
  OAI22X1 U626 ( .A0(n976), .A1(n164), .B0(n9), .B1(n163), .Y(n181) );
  OAI22XL U627 ( .A0(n240), .A1(n171), .B0(n170), .B1(n1085), .Y(n175) );
  OAI22XL U628 ( .A0(n979), .A1(n173), .B0(n757), .B1(n172), .Y(n174) );
  NAND2XL U629 ( .A(n1213), .B(n1257), .Y(n1214) );
  INVXL U630 ( .A(n1247), .Y(n1248) );
  INVXL U631 ( .A(B[0]), .Y(n489) );
  OAI22XL U632 ( .A0(n1100), .A1(n348), .B0(n1101), .B1(n343), .Y(n357) );
  OAI22XL U633 ( .A0(n1135), .A1(n317), .B0(n1136), .B1(n313), .Y(n323) );
  XNOR2XL U634 ( .A(n1156), .B(A[17]), .Y(n301) );
  OAI22XL U635 ( .A0(n1135), .A1(n327), .B0(n1136), .B1(n1102), .Y(n1109) );
  OAI22XL U636 ( .A0(n1135), .A1(n1102), .B0(n1136), .B1(n1121), .Y(n1124) );
  OAI2BB1XL U637 ( .A0N(n1101), .A1N(n1100), .B0(n1099), .Y(n1115) );
  INVXL U638 ( .A(n1098), .Y(n1099) );
  XNOR3X2 U639 ( .A(n89), .B(n933), .C(n934), .Y(n942) );
  ADDFX2 U640 ( .A(n762), .B(n761), .CI(n760), .CO(n741), .S(n778) );
  OAI22XL U641 ( .A0(n926), .A1(n756), .B0(n757), .B1(n719), .Y(n762) );
  OAI22XL U642 ( .A0(n1135), .A1(n759), .B0(n954), .B1(n721), .Y(n760) );
  ADDFX2 U643 ( .A(n791), .B(n790), .CI(n789), .CO(n779), .S(n806) );
  OAI22XL U644 ( .A0(n1135), .A1(n788), .B0(n954), .B1(n759), .Y(n789) );
  OAI22X1 U645 ( .A0(n7), .A1(n787), .B0(n8), .B1(n758), .Y(n790) );
  OAI22XL U646 ( .A0(n926), .A1(n786), .B0(n757), .B1(n756), .Y(n791) );
  ADDFX2 U647 ( .A(n486), .B(n485), .CI(n484), .CO(n503), .S(n548) );
  INVX4 U648 ( .A(n102), .Y(n905) );
  INVX1 U649 ( .A(B[1]), .Y(n102) );
  NOR2BXL U650 ( .AN(A[0]), .B(n968), .Y(n129) );
  OAI22XL U651 ( .A0(n240), .A1(n126), .B0(n132), .B1(n1085), .Y(n130) );
  OAI22XL U652 ( .A0(n1161), .A1(n1128), .B0(n8), .B1(n1139), .Y(n1148) );
  NAND2X1 U653 ( .A(n72), .B(n96), .Y(n936) );
  NAND2X1 U654 ( .A(n88), .B(n87), .Y(n899) );
  NAND2X1 U655 ( .A(n934), .B(n935), .Y(n87) );
  OAI21XL U656 ( .A0(n934), .A1(n935), .B0(n933), .Y(n88) );
  XOR3X2 U657 ( .A(n944), .B(n942), .C(n943), .Y(n986) );
  OAI2BB1X1 U658 ( .A0N(n69), .A1N(n1010), .B0(n68), .Y(n990) );
  XOR3X2 U659 ( .A(n1012), .B(n1011), .C(n1010), .Y(n1018) );
  INVXL U660 ( .A(mult_x_1_n306), .Y(n1063) );
  INVXL U661 ( .A(n275), .Y(n1065) );
  AOI21XL U662 ( .A0(n289), .A1(n235), .B0(n234), .Y(n1066) );
  NAND2XL U663 ( .A(n130), .B(n129), .Y(n1216) );
  NAND2XL U664 ( .A(n1152), .B(n1151), .Y(mult_x_1_n121) );
  NOR2BXL U665 ( .AN(A[0]), .B(n1085), .Y(n1335) );
  XOR2XL U666 ( .A(n1073), .B(n1072), .Y(n1325) );
  NAND2XL U667 ( .A(n1076), .B(n1075), .Y(n1077) );
  NOR2XL U668 ( .A(n1093), .B(n1092), .Y(mult_x_1_n151) );
  NOR2XL U669 ( .A(n1111), .B(n1110), .Y(mult_x_1_n136) );
  NOR2XL U670 ( .A(n551), .B(n550), .Y(mult_x_1_n197) );
  NAND2XL U671 ( .A(n1168), .B(n1167), .Y(mult_x_1_n58) );
  NAND2XL U672 ( .A(n1166), .B(n1165), .Y(n1167) );
  NOR2XL U673 ( .A(n1150), .B(n1149), .Y(mult_x_1_n109) );
  NAND2XL U674 ( .A(n1150), .B(n1149), .Y(mult_x_1_n110) );
  NOR2XL U675 ( .A(n1152), .B(n1151), .Y(mult_x_1_n120) );
  NOR2XL U676 ( .A(n1126), .B(n1125), .Y(mult_x_1_n129) );
  NAND2XL U677 ( .A(n1126), .B(n1125), .Y(mult_x_1_n130) );
  NAND2XL U678 ( .A(n1111), .B(n1110), .Y(mult_x_1_n137) );
  NOR2XL U679 ( .A(n588), .B(n587), .Y(mult_x_1_n206) );
  NAND2XL U680 ( .A(n1014), .B(n1013), .Y(mult_x_1_n287) );
  XNOR2XL U681 ( .A(n1219), .B(n1218), .Y(n1333) );
  NAND2XL U682 ( .A(n1217), .B(n1216), .Y(n1219) );
  NAND2XL U683 ( .A(n1229), .B(n1228), .Y(n1231) );
  INVXL U684 ( .A(n1227), .Y(n1229) );
  NAND2XL U685 ( .A(n144), .B(n1224), .Y(n1226) );
  NAND2XL U686 ( .A(n1234), .B(n1233), .Y(n1236) );
  INVXL U687 ( .A(n1232), .Y(n1234) );
  XOR2XL U688 ( .A(n1202), .B(n1201), .Y(n1329) );
  NAND2XL U689 ( .A(n85), .B(n1200), .Y(n1202) );
  NAND2XL U690 ( .A(n1192), .B(n1191), .Y(n1193) );
  XNOR2XL U691 ( .A(n1172), .B(n1171), .Y(n1327) );
  NAND2XL U692 ( .A(n1170), .B(n1169), .Y(n1171) );
  OAI21XL U693 ( .A0(n1288), .A1(n1291), .B0(n1289), .Y(n710) );
  CLKINVX3 U694 ( .A(B[7]), .Y(n303) );
  AND2X1 U695 ( .A(n292), .B(n291), .Y(n66) );
  XNOR2X1 U696 ( .A(n474), .B(n473), .Y(PRODUCT[30]) );
  CMPR22X1 U697 ( .A(n645), .B(n644), .CO(n616), .S(n656) );
  CMPR22X1 U698 ( .A(n687), .B(n686), .CO(n655), .S(n696) );
  CMPR22X1 U699 ( .A(n765), .B(n764), .CO(n736), .S(n775) );
  CMPR22X1 U700 ( .A(n829), .B(n828), .CO(n802), .S(n840) );
  OAI22X1 U701 ( .A0(n926), .A1(n378), .B0(n757), .B1(n304), .Y(n353) );
  BUFX1 U702 ( .A(n119), .Y(n67) );
  CMPR22X1 U703 ( .A(n253), .B(n252), .CO(n267), .S(n260) );
  CMPR22X1 U704 ( .A(n166), .B(n165), .CO(n180), .S(n188) );
  OAI22X1 U705 ( .A0(n926), .A1(n303), .B0(n757), .B1(n104), .Y(n165) );
  CMPR22X1 U706 ( .A(n607), .B(n606), .CO(n575), .S(n617) );
  OAI22X1 U707 ( .A0(n643), .A1(n315), .B0(n960), .B1(n310), .Y(n329) );
  CMPR22X1 U708 ( .A(n143), .B(n142), .CO(n145), .S(n138) );
  OAI22X1 U709 ( .A0(n133), .A1(n970), .B0(n968), .B1(n93), .Y(n142) );
  XNOR2X1 U710 ( .A(n1089), .B(n1088), .Y(PRODUCT[22]) );
  XNOR2XL U711 ( .A(n1156), .B(A[1]), .Y(n862) );
  CMPR22X1 U712 ( .A(n529), .B(n528), .CO(n542), .S(n576) );
  OAI21XL U713 ( .A0(n116), .A1(n117), .B0(n79), .Y(n76) );
  AOI2BB1X1 U714 ( .A0N(n275), .A1N(n1068), .B0(n286), .Y(n287) );
  OAI22X1 U715 ( .A0(n307), .A1(n308), .B0(n1101), .B1(n194), .Y(n252) );
  OAI21X1 U716 ( .A0(n1073), .A1(n1069), .B0(n1070), .Y(n293) );
  INVX4 U717 ( .A(n169), .Y(n908) );
  NAND2X4 U718 ( .A(n75), .B(n237), .Y(n1135) );
  OAI21XL U719 ( .A0(n110), .A1(n9), .B0(n80), .Y(n79) );
  NAND3BX1 U720 ( .AN(n1190), .B(n1189), .C(n85), .Y(n84) );
  XOR2X1 U721 ( .A(n293), .B(n66), .Y(n1324) );
  INVX1 U722 ( .A(n289), .Y(n1073) );
  NAND3X1 U723 ( .A(n1172), .B(n1076), .C(n1170), .Y(n86) );
  XOR2X1 U724 ( .A(n650), .B(n91), .Y(n90) );
  OAI22X2 U725 ( .A0(n648), .A1(n964), .B0(n966), .B1(n98), .Y(n694) );
  XNOR2X1 U726 ( .A(B[6]), .B(B[5]), .Y(n105) );
  OAI22X1 U727 ( .A0(n962), .A1(n200), .B0(n960), .B1(n199), .Y(n204) );
  INVX1 U728 ( .A(n1308), .Y(n1062) );
  AOI21X1 U729 ( .A0(n295), .A1(n555), .B0(n294), .Y(n296) );
  CMPR22X1 U730 ( .A(n950), .B(n949), .CO(n958), .S(n999) );
  OAI22X1 U731 ( .A0(n966), .A1(n241), .B0(n964), .B1(n247), .Y(n254) );
  OAI22X1 U732 ( .A0(n966), .A1(n768), .B0(n964), .B1(n730), .Y(n773) );
  OAI22X1 U733 ( .A0(n966), .A1(n213), .B0(n964), .B1(n241), .Y(n258) );
  NAND2X2 U734 ( .A(n160), .B(n685), .Y(n643) );
  XOR2X1 U735 ( .A(n1250), .B(n509), .Y(PRODUCT[29]) );
  NAND2X2 U736 ( .A(n193), .B(n212), .Y(n307) );
  XNOR2X2 U737 ( .A(B[10]), .B(B[9]), .Y(n212) );
  XOR2XL U738 ( .A(B[2]), .B(B[3]), .Y(n108) );
  XNOR2X1 U739 ( .A(n650), .B(A[2]), .Y(n110) );
  BUFX3 U740 ( .A(n212), .Y(n964) );
  XNOR2X1 U741 ( .A(n650), .B(A[24]), .Y(n419) );
  XNOR2XL U742 ( .A(n905), .B(A[3]), .Y(n140) );
  OAI22X1 U743 ( .A0(n976), .A1(n419), .B0(n9), .B1(n370), .Y(n390) );
  OR2X2 U744 ( .A(n190), .B(n189), .Y(n1170) );
  OAI21XL U745 ( .A0(n1066), .A1(n288), .B0(n287), .Y(mult_x_1_n309) );
  NAND2X1 U746 ( .A(B[1]), .B(n489), .Y(n127) );
  BUFX3 U747 ( .A(n127), .Y(n240) );
  BUFX3 U748 ( .A(n489), .Y(n1085) );
  OAI22X1 U749 ( .A0(n240), .A1(n106), .B0(n171), .B1(n1085), .Y(n166) );
  BUFX3 U750 ( .A(n105), .Y(n757) );
  CLKINVX8 U751 ( .A(n303), .Y(n924) );
  XOR2X1 U752 ( .A(B[4]), .B(B[5]), .Y(n107) );
  XNOR2X1 U753 ( .A(B[4]), .B(B[3]), .Y(n113) );
  XNOR2XL U754 ( .A(B[2]), .B(B[1]), .Y(n134) );
  BUFX3 U755 ( .A(n134), .Y(n968) );
  XNOR2X1 U756 ( .A(n924), .B(A[0]), .Y(n109) );
  XNOR2X1 U757 ( .A(n924), .B(A[1]), .Y(n173) );
  XNOR2X1 U758 ( .A(n650), .B(A[3]), .Y(n164) );
  OAI22XL U759 ( .A0(n835), .A1(n110), .B0(n9), .B1(n164), .Y(n177) );
  OAI22XL U760 ( .A0(n976), .A1(n115), .B0(n9), .B1(n114), .Y(n124) );
  XNOR2X1 U761 ( .A(n650), .B(A[0]), .Y(n123) );
  OAI22XL U762 ( .A0(n835), .A1(n123), .B0(n9), .B1(n122), .Y(n149) );
  ADDHXL U763 ( .A(n125), .B(n124), .CO(n119), .S(n148) );
  OR2X2 U764 ( .A(n130), .B(n129), .Y(n1217) );
  OAI22X1 U765 ( .A0(n240), .A1(n132), .B0(n140), .B1(n1085), .Y(n143) );
  AOI21XL U766 ( .A0(n1225), .A1(n144), .B0(n147), .Y(n1235) );
  CMPR32X1 U767 ( .A(n150), .B(n149), .C(n148), .CO(n156), .S(n155) );
  CMPR32X1 U768 ( .A(n153), .B(n152), .C(n151), .CO(n154), .S(n146) );
  OAI21XL U769 ( .A0(n1235), .A1(n1232), .B0(n1233), .Y(n1189) );
  XNOR2X1 U770 ( .A(n924), .B(A[2]), .Y(n172) );
  XOR2X1 U771 ( .A(B[8]), .B(B[9]), .Y(n160) );
  INVX2 U772 ( .A(B[9]), .Y(n169) );
  XNOR2XL U773 ( .A(n908), .B(A[0]), .Y(n161) );
  XNOR2X1 U774 ( .A(n908), .B(A[1]), .Y(n200) );
  XNOR2X1 U775 ( .A(n650), .B(A[5]), .Y(n209) );
  XNOR2X1 U776 ( .A(n919), .B(A[7]), .Y(n210) );
  OAI22XL U777 ( .A0(n643), .A1(n169), .B0(n685), .B1(n168), .Y(n195) );
  CMPR32X1 U778 ( .A(n176), .B(n175), .C(n174), .CO(n218), .S(n185) );
  CMPR32X1 U779 ( .A(n188), .B(n187), .C(n186), .CO(n189), .S(n159) );
  NAND2XL U780 ( .A(n190), .B(n189), .Y(n1169) );
  INVXL U781 ( .A(n1169), .Y(n1074) );
  OAI22X1 U782 ( .A0(n976), .A1(n208), .B0(n9), .B1(n244), .Y(n262) );
  XNOR2XL U783 ( .A(n908), .B(A[2]), .Y(n199) );
  OAI22X1 U784 ( .A0(n962), .A1(n199), .B0(n960), .B1(n251), .Y(n261) );
  OAI22X1 U785 ( .A0(n240), .A1(n197), .B0(n239), .B1(n1085), .Y(n253) );
  XOR2X1 U786 ( .A(B[10]), .B(B[11]), .Y(n193) );
  INVX8 U787 ( .A(n308), .Y(n922) );
  CMPR32X1 U788 ( .A(n206), .B(n205), .C(n204), .CO(n271), .S(n222) );
  XNOR2X1 U789 ( .A(n924), .B(A[4]), .Y(n211) );
  OAI22X1 U790 ( .A0(n976), .A1(n209), .B0(n9), .B1(n208), .Y(n216) );
  XNOR2X1 U791 ( .A(n922), .B(A[0]), .Y(n213) );
  XNOR2X1 U792 ( .A(n922), .B(A[1]), .Y(n241) );
  ADDFHX1 U793 ( .A(n217), .B(n216), .CI(n215), .CO(n270), .S(n226) );
  CMPR32X1 U794 ( .A(n220), .B(n219), .C(n218), .CO(n225), .S(n227) );
  NOR2X1 U795 ( .A(n233), .B(n232), .Y(n290) );
  CMPR32X1 U796 ( .A(n226), .B(n225), .C(n224), .CO(n232), .S(n231) );
  NOR2XL U797 ( .A(n290), .B(n1069), .Y(n235) );
  NAND2XL U798 ( .A(n231), .B(n230), .Y(n1070) );
  NAND2XL U799 ( .A(n233), .B(n232), .Y(n291) );
  OAI21XL U800 ( .A0(n290), .A1(n1070), .B0(n291), .Y(n234) );
  BUFX3 U801 ( .A(n237), .Y(n1136) );
  BUFX3 U802 ( .A(n237), .Y(n954) );
  NOR2BX1 U803 ( .AN(A[0]), .B(n954), .Y(n256) );
  OAI22X1 U804 ( .A0(n240), .A1(n239), .B0(n238), .B1(n1085), .Y(n255) );
  XNOR2X1 U805 ( .A(n922), .B(A[2]), .Y(n247) );
  XNOR2X1 U806 ( .A(n924), .B(A[6]), .Y(n245) );
  XNOR2X1 U807 ( .A(n650), .B(A[8]), .Y(n249) );
  OAI22XL U808 ( .A0(n926), .A1(n245), .B0(n757), .B1(n978), .Y(n1026) );
  OAI22X1 U809 ( .A0(n1135), .A1(n246), .B0(n954), .B1(n955), .Y(n1025) );
  XNOR2X1 U810 ( .A(n922), .B(A[3]), .Y(n965) );
  XNOR2X1 U811 ( .A(n919), .B(A[11]), .Y(n969) );
  XNOR2X1 U812 ( .A(n650), .B(A[9]), .Y(n975) );
  CMPR32X1 U813 ( .A(n256), .B(n255), .C(n254), .CO(n1031), .S(n266) );
  CMPR32X1 U814 ( .A(n259), .B(n258), .C(n257), .CO(n274), .S(n269) );
  CMPR32X1 U815 ( .A(n262), .B(n261), .C(n260), .CO(n273), .S(n281) );
  CMPR32X1 U816 ( .A(n265), .B(n264), .C(n263), .CO(n1030), .S(n272) );
  CMPR32X1 U817 ( .A(n268), .B(n267), .C(n266), .CO(n1041), .S(n278) );
  CMPR32X1 U818 ( .A(n271), .B(n270), .C(n269), .CO(n277), .S(n279) );
  CMPR32X1 U819 ( .A(n274), .B(n273), .C(n272), .CO(n1047), .S(n276) );
  NOR2X1 U820 ( .A(n285), .B(n284), .Y(n275) );
  CMPR32X1 U821 ( .A(n281), .B(n280), .C(n279), .CO(n282), .S(n233) );
  NAND2XL U822 ( .A(n1065), .B(n6), .Y(n288) );
  INVXL U823 ( .A(n1068), .Y(n1067) );
  NAND2XL U824 ( .A(n285), .B(n284), .Y(n1064) );
  INVXL U825 ( .A(n1064), .Y(n286) );
  INVXL U826 ( .A(n290), .Y(n292) );
  NOR2X1 U827 ( .A(n1280), .B(n1278), .Y(n295) );
  OAI21XL U828 ( .A0(n1278), .A1(n1281), .B0(n1279), .Y(n294) );
  NOR2XL U829 ( .A(n1272), .B(n1270), .Y(n298) );
  NAND2XL U830 ( .A(n439), .B(n298), .Y(n1239) );
  OAI21XL U831 ( .A0(n1270), .A1(n1273), .B0(n1271), .Y(n297) );
  XNOR2X2 U832 ( .A(B[16]), .B(B[15]), .Y(n384) );
  BUFX3 U833 ( .A(n384), .Y(n1158) );
  BUFX8 U834 ( .A(B[16]), .Y(n1156) );
  XNOR2XL U835 ( .A(n924), .B(A[24]), .Y(n378) );
  XNOR2XL U836 ( .A(n924), .B(A[25]), .Y(n304) );
  INVXL U837 ( .A(n304), .Y(n305) );
  CLKINVX3 U838 ( .A(n306), .Y(n1127) );
  XNOR2XL U839 ( .A(n1127), .B(A[18]), .Y(n316) );
  OAI22XL U840 ( .A0(n1161), .A1(n316), .B0(n8), .B1(n312), .Y(n320) );
  BUFX3 U841 ( .A(n307), .Y(n1100) );
  OAI22XL U842 ( .A0(n1100), .A1(n343), .B0(n1101), .B1(n314), .Y(n319) );
  XNOR2XL U843 ( .A(n908), .B(A[25]), .Y(n310) );
  OAI22XL U844 ( .A0(n1161), .A1(n312), .B0(n8), .B1(n324), .Y(n333) );
  XNOR2X1 U845 ( .A(n1127), .B(A[17]), .Y(n347) );
  OAI22XL U846 ( .A0(n1161), .A1(n347), .B0(n8), .B1(n316), .Y(n350) );
  CMPR32X1 U847 ( .A(n320), .B(n319), .C(n318), .CO(n336), .S(n359) );
  CMPR32X1 U848 ( .A(n323), .B(n322), .C(n321), .CO(n363), .S(n358) );
  XNOR2X1 U849 ( .A(n922), .B(A[25]), .Y(n1098) );
  OAI22X1 U850 ( .A0(n1100), .A1(n326), .B0(n1101), .B1(n1098), .Y(n1116) );
  CMPR32X1 U851 ( .A(n330), .B(n329), .C(n328), .CO(n1108), .S(n335) );
  CMPR32X1 U852 ( .A(n333), .B(n332), .C(n331), .CO(n1107), .S(n334) );
  CMPR32X1 U853 ( .A(n336), .B(n335), .C(n334), .CO(n1094), .S(n362) );
  NAND2XL U854 ( .A(n1093), .B(n1092), .Y(mult_x_1_n152) );
  INVXL U855 ( .A(n337), .Y(n340) );
  INVXL U856 ( .A(n338), .Y(n339) );
  XNOR2X1 U857 ( .A(n342), .B(n341), .Y(PRODUCT[34]) );
  INVXL U858 ( .A(n353), .Y(n375) );
  CMPR32X1 U859 ( .A(n351), .B(n350), .C(n349), .CO(n360), .S(n397) );
  CMPR32X1 U860 ( .A(n354), .B(n353), .C(n352), .CO(n321), .S(n396) );
  ADDFHX1 U861 ( .A(n357), .B(n356), .CI(n355), .CO(n400), .S(n395) );
  CMPR32X1 U862 ( .A(n360), .B(n359), .C(n358), .CO(n361), .S(n398) );
  CMPR32X1 U863 ( .A(n363), .B(n362), .C(n361), .CO(n1093), .S(n364) );
  NOR2XL U864 ( .A(n365), .B(n364), .Y(mult_x_1_n160) );
  NAND2XL U865 ( .A(n365), .B(n364), .Y(mult_x_1_n161) );
  CMPR32X1 U866 ( .A(n374), .B(n373), .C(n372), .CO(n355), .S(n410) );
  XNOR2X1 U867 ( .A(n924), .B(A[23]), .Y(n386) );
  OAI22XL U868 ( .A0(n926), .A1(n386), .B0(n757), .B1(n378), .Y(n394) );
  XNOR2X1 U869 ( .A(n1120), .B(A[17]), .Y(n383) );
  XNOR2X1 U870 ( .A(n1120), .B(A[16]), .Y(n423) );
  XNOR2XL U871 ( .A(n1156), .B(A[13]), .Y(n385) );
  NOR2XL U872 ( .A(n384), .B(n385), .Y(n426) );
  XNOR2X1 U873 ( .A(n924), .B(A[22]), .Y(n421) );
  OAI22XL U874 ( .A0(n926), .A1(n421), .B0(n757), .B1(n386), .Y(n430) );
  INVX8 U875 ( .A(n306), .Y(n1138) );
  OAI22X1 U876 ( .A0(n7), .A1(n420), .B0(n8), .B1(n387), .Y(n429) );
  OAI22XL U877 ( .A0(n1100), .A1(n424), .B0(n1101), .B1(n388), .Y(n428) );
  CMPR32X1 U878 ( .A(n391), .B(n390), .C(n389), .CO(n411), .S(n450) );
  CMPR32X1 U879 ( .A(n394), .B(n393), .C(n392), .CO(n433), .S(n449) );
  CMPR32X1 U880 ( .A(n397), .B(n396), .C(n395), .CO(n399), .S(n434) );
  CMPR32X1 U881 ( .A(n400), .B(n399), .C(n398), .CO(n365), .S(n401) );
  NOR2XL U882 ( .A(n402), .B(n401), .Y(mult_x_1_n169) );
  NAND2XL U883 ( .A(n402), .B(n401), .Y(mult_x_1_n170) );
  AOI21XL U884 ( .A0(n440), .A1(n443), .B0(n403), .Y(n404) );
  INVXL U885 ( .A(n1270), .Y(n406) );
  CMPR32X1 U886 ( .A(n411), .B(n410), .C(n409), .CO(n436), .S(n448) );
  CMPR32X1 U887 ( .A(n414), .B(n413), .C(n412), .CO(n432), .S(n454) );
  XNOR2XL U888 ( .A(n1156), .B(A[12]), .Y(n416) );
  XNOR2X1 U889 ( .A(n650), .B(A[23]), .Y(n476) );
  OAI22X1 U890 ( .A0(n976), .A1(n476), .B0(n9), .B1(n419), .Y(n463) );
  XNOR2X1 U891 ( .A(n1138), .B(A[13]), .Y(n460) );
  OAI22X2 U892 ( .A0(n7), .A1(n460), .B0(n8), .B1(n420), .Y(n462) );
  OAI22XL U893 ( .A0(n926), .A1(n458), .B0(n757), .B1(n421), .Y(n461) );
  XNOR2XL U894 ( .A(n908), .B(A[19]), .Y(n480) );
  OAI22XL U895 ( .A0(n962), .A1(n480), .B0(n960), .B1(n422), .Y(n466) );
  XNOR2X1 U896 ( .A(n1120), .B(A[15]), .Y(n475) );
  OAI22X1 U897 ( .A0(n1135), .A1(n475), .B0(n1136), .B1(n423), .Y(n465) );
  OAI22XL U898 ( .A0(n1100), .A1(n481), .B0(n1101), .B1(n424), .Y(n464) );
  ADDFHX1 U899 ( .A(n430), .B(n429), .CI(n428), .CO(n451), .S(n467) );
  ADDFHX1 U900 ( .A(n433), .B(n432), .CI(n431), .CO(n435), .S(n446) );
  CMPR32X1 U901 ( .A(n436), .B(n435), .C(n434), .CO(n402), .S(n437) );
  NOR2XL U902 ( .A(n438), .B(n437), .Y(mult_x_1_n176) );
  NAND2XL U903 ( .A(n438), .B(n437), .Y(mult_x_1_n177) );
  OAI21XL U904 ( .A0(n1250), .A1(n442), .B0(n441), .Y(n445) );
  ADDFHX1 U905 ( .A(n448), .B(n447), .CI(n446), .CO(n438), .S(n471) );
  CMPR32X1 U906 ( .A(n451), .B(n450), .C(n449), .CO(n431), .S(n505) );
  CMPR32X1 U907 ( .A(n454), .B(n453), .C(n452), .CO(n447), .S(n504) );
  XNOR2X1 U908 ( .A(n924), .B(A[20]), .Y(n482) );
  XNOR2X1 U909 ( .A(n1156), .B(A[11]), .Y(n459) );
  XNOR2X1 U910 ( .A(n1138), .B(A[12]), .Y(n483) );
  OAI22XL U911 ( .A0(n7), .A1(n483), .B0(n8), .B1(n460), .Y(n513) );
  CMPR32X1 U912 ( .A(n466), .B(n465), .C(n464), .CO(n469), .S(n497) );
  CMPR32X1 U913 ( .A(n469), .B(n468), .C(n467), .CO(n452), .S(n484) );
  NOR2XL U914 ( .A(n471), .B(n470), .Y(mult_x_1_n183) );
  NAND2XL U915 ( .A(n471), .B(n470), .Y(mult_x_1_n184) );
  OAI21X2 U916 ( .A0(n1250), .A1(n1276), .B0(n1277), .Y(n474) );
  INVXL U917 ( .A(n1274), .Y(n472) );
  XNOR2X1 U918 ( .A(n650), .B(A[22]), .Y(n510) );
  OAI22XL U919 ( .A0(n976), .A1(n510), .B0(n9), .B1(n476), .Y(n492) );
  OAI22XL U920 ( .A0(n1100), .A1(n487), .B0(n1101), .B1(n481), .Y(n495) );
  XNOR2X1 U921 ( .A(n924), .B(A[19]), .Y(n535) );
  OAI22X1 U922 ( .A0(n1100), .A1(n521), .B0(n1101), .B1(n487), .Y(n526) );
  XNOR2X1 U923 ( .A(n919), .B(A[23]), .Y(n522) );
  CMPR32X1 U924 ( .A(n496), .B(n495), .C(n494), .CO(n500), .S(n566) );
  CMPR32X1 U925 ( .A(n502), .B(n501), .C(n500), .CO(n549), .S(n544) );
  ADDFHX1 U926 ( .A(n505), .B(n504), .CI(n503), .CO(n470), .S(n506) );
  NOR2XL U927 ( .A(n507), .B(n506), .Y(mult_x_1_n194) );
  NAND2XL U928 ( .A(n507), .B(n506), .Y(mult_x_1_n195) );
  NAND2XL U929 ( .A(n508), .B(n1277), .Y(n509) );
  XNOR2X1 U930 ( .A(n1120), .B(A[13]), .Y(n537) );
  OAI22X1 U931 ( .A0(n240), .A1(n530), .B0(n517), .B1(n1085), .Y(n529) );
  XNOR2X1 U932 ( .A(n1156), .B(A[9]), .Y(n518) );
  NOR2XL U933 ( .A(n384), .B(n518), .Y(n528) );
  XNOR2X1 U934 ( .A(n922), .B(n904), .Y(n569) );
  XNOR2X1 U935 ( .A(n650), .B(A[20]), .Y(n571) );
  XNOR2XL U936 ( .A(n908), .B(A[16]), .Y(n605) );
  OAI22X1 U937 ( .A0(n127), .A1(n608), .B0(n530), .B1(n1085), .Y(n607) );
  XNOR2XL U938 ( .A(n1156), .B(A[8]), .Y(n531) );
  NOR2XL U939 ( .A(n384), .B(n531), .Y(n606) );
  XNOR2X1 U940 ( .A(n924), .B(A[18]), .Y(n599) );
  OAI22X1 U941 ( .A0(n926), .A1(n599), .B0(n757), .B1(n535), .Y(n604) );
  XNOR2X2 U942 ( .A(n1138), .B(A[10]), .Y(n600) );
  OAI22X2 U943 ( .A0(n7), .A1(n600), .B0(n8), .B1(n536), .Y(n603) );
  XNOR2X1 U944 ( .A(n1120), .B(A[12]), .Y(n601) );
  OAI22X1 U945 ( .A0(n1135), .A1(n601), .B0(n954), .B1(n537), .Y(n602) );
  CMPR32X1 U946 ( .A(n543), .B(n542), .C(n541), .CO(n532), .S(n581) );
  CMPR32X1 U947 ( .A(n546), .B(n545), .C(n544), .CO(n547), .S(n563) );
  INVXL U948 ( .A(n552), .Y(n589) );
  NOR2XL U949 ( .A(n589), .B(n1280), .Y(n557) );
  OAI21XL U950 ( .A0(n590), .A1(n1280), .B0(n1281), .Y(n556) );
  OAI22X1 U951 ( .A0(n1100), .A1(n610), .B0(n1101), .B1(n569), .Y(n615) );
  XNOR2X1 U952 ( .A(n650), .B(A[19]), .Y(n612) );
  NAND2XL U953 ( .A(n588), .B(n587), .Y(mult_x_1_n207) );
  AOI21XL U954 ( .A0(n670), .A1(n552), .B0(n555), .Y(n591) );
  ADDFHX1 U955 ( .A(n598), .B(n597), .CI(n596), .CO(n587), .S(n629) );
  OAI22X1 U956 ( .A0(n926), .A1(n636), .B0(n757), .B1(n599), .Y(n641) );
  OAI22X2 U957 ( .A0(n7), .A1(n637), .B0(n8), .B1(n600), .Y(n640) );
  OAI22XL U958 ( .A0(n643), .A1(n642), .B0(n960), .B1(n605), .Y(n618) );
  OAI22X1 U959 ( .A0(n240), .A1(n646), .B0(n608), .B1(n1085), .Y(n645) );
  XNOR2XL U960 ( .A(n1156), .B(A[7]), .Y(n609) );
  NOR2XL U961 ( .A(n384), .B(n609), .Y(n644) );
  XNOR2X1 U962 ( .A(n922), .B(A[12]), .Y(n648) );
  OAI22X2 U963 ( .A0(n970), .A1(n649), .B0(n968), .B1(n611), .Y(n653) );
  XNOR2X1 U964 ( .A(n650), .B(A[18]), .Y(n651) );
  CMPR32X1 U965 ( .A(n618), .B(n617), .C(n616), .CO(n619), .S(n661) );
  CMPR32X1 U966 ( .A(n621), .B(n620), .C(n619), .CO(n635), .S(n665) );
  NOR2XL U967 ( .A(n629), .B(n628), .Y(mult_x_1_n215) );
  NAND2XL U968 ( .A(n629), .B(n628), .Y(mult_x_1_n216) );
  ADDFHX1 U969 ( .A(n635), .B(n634), .CI(n633), .CO(n628), .S(n668) );
  XNOR2X1 U970 ( .A(n924), .B(A[16]), .Y(n678) );
  OAI22X1 U971 ( .A0(n926), .A1(n678), .B0(n757), .B1(n636), .Y(n683) );
  XNOR2X1 U972 ( .A(n1138), .B(A[8]), .Y(n679) );
  OAI22X2 U973 ( .A0(n7), .A1(n679), .B0(n8), .B1(n637), .Y(n682) );
  OAI22X1 U974 ( .A0(n1135), .A1(n680), .B0(n954), .B1(n638), .Y(n681) );
  XNOR2X1 U975 ( .A(n908), .B(n904), .Y(n684) );
  OAI22XL U976 ( .A0(n643), .A1(n684), .B0(n960), .B1(n642), .Y(n657) );
  OAI22X1 U977 ( .A0(n127), .A1(n688), .B0(n646), .B1(n1085), .Y(n687) );
  XNOR2XL U978 ( .A(n1156), .B(A[6]), .Y(n647) );
  NOR2XL U979 ( .A(n384), .B(n647), .Y(n686) );
  OAI22X2 U980 ( .A0(n970), .A1(n690), .B0(n968), .B1(n649), .Y(n693) );
  XNOR2X1 U981 ( .A(n650), .B(A[17]), .Y(n691) );
  CMPR32X1 U982 ( .A(n657), .B(n656), .C(n655), .CO(n658), .S(n701) );
  CMPR32X1 U983 ( .A(n660), .B(n659), .C(n658), .CO(n677), .S(n705) );
  CMPR32X1 U984 ( .A(n666), .B(n665), .C(n664), .CO(n634), .S(n675) );
  NOR2XL U985 ( .A(n668), .B(n667), .Y(mult_x_1_n226) );
  NAND2XL U986 ( .A(n668), .B(n667), .Y(mult_x_1_n227) );
  OAI21XL U987 ( .A0(n1086), .A1(n553), .B0(n671), .Y(n674) );
  XNOR2X1 U988 ( .A(n674), .B(n673), .Y(PRODUCT[25]) );
  ADDFHX1 U989 ( .A(n677), .B(n676), .CI(n675), .CO(n667), .S(n708) );
  OAI22X1 U990 ( .A0(n926), .A1(n719), .B0(n757), .B1(n678), .Y(n724) );
  OAI22X1 U991 ( .A0(n1135), .A1(n721), .B0(n954), .B1(n680), .Y(n722) );
  OAI22XL U992 ( .A0(n962), .A1(n725), .B0(n685), .B1(n684), .Y(n697) );
  XNOR2XL U993 ( .A(n1156), .B(A[5]), .Y(n689) );
  NOR2XL U994 ( .A(n384), .B(n689), .Y(n726) );
  XNOR2X1 U995 ( .A(n922), .B(A[10]), .Y(n730) );
  OAI22X2 U996 ( .A0(n970), .A1(n731), .B0(n968), .B1(n690), .Y(n734) );
  XNOR2X1 U997 ( .A(n650), .B(A[16]), .Y(n732) );
  CMPR32X1 U998 ( .A(n697), .B(n696), .C(n695), .CO(n698), .S(n742) );
  CMPR32X1 U999 ( .A(n700), .B(n699), .C(n698), .CO(n718), .S(n746) );
  CMPR32X1 U1000 ( .A(n706), .B(n705), .C(n704), .CO(n676), .S(n716) );
  NOR2XL U1001 ( .A(n708), .B(n707), .Y(mult_x_1_n233) );
  NAND2XL U1002 ( .A(n750), .B(n753), .Y(n714) );
  INVXL U1003 ( .A(n752), .Y(n712) );
  INVXL U1004 ( .A(n1286), .Y(n715) );
  ADDFHX1 U1005 ( .A(n718), .B(n717), .CI(n716), .CO(n707), .S(n749) );
  XNOR2XL U1006 ( .A(n908), .B(A[12]), .Y(n763) );
  OAI22XL U1007 ( .A0(n962), .A1(n763), .B0(n960), .B1(n725), .Y(n738) );
  ADDHXL U1008 ( .A(n727), .B(n726), .CO(n695), .S(n737) );
  OAI22X1 U1009 ( .A0(n127), .A1(n766), .B0(n728), .B1(n1085), .Y(n765) );
  XNOR2XL U1010 ( .A(n1156), .B(A[4]), .Y(n729) );
  NOR2XL U1011 ( .A(n384), .B(n729), .Y(n764) );
  XNOR2X1 U1012 ( .A(n922), .B(A[9]), .Y(n768) );
  XNOR2X1 U1013 ( .A(n650), .B(A[15]), .Y(n770) );
  CMPR32X1 U1014 ( .A(n738), .B(n736), .C(n737), .CO(n739), .S(n780) );
  CMPR32X1 U1015 ( .A(n747), .B(n746), .C(n745), .CO(n717), .S(n1079) );
  NOR2XL U1016 ( .A(n749), .B(n748), .Y(mult_x_1_n244) );
  NAND2XL U1017 ( .A(n749), .B(n748), .Y(mult_x_1_n245) );
  INVXL U1018 ( .A(n750), .Y(n751) );
  OAI21XL U1019 ( .A0(n1086), .A1(n751), .B0(n711), .Y(n755) );
  NAND2X1 U1020 ( .A(n753), .B(n752), .Y(n754) );
  XNOR2X1 U1021 ( .A(n755), .B(n754), .Y(PRODUCT[23]) );
  XNOR2XL U1022 ( .A(n908), .B(A[11]), .Y(n792) );
  OAI22XL U1023 ( .A0(n962), .A1(n792), .B0(n960), .B1(n763), .Y(n776) );
  XNOR2XL U1024 ( .A(n1156), .B(A[3]), .Y(n767) );
  NOR2XL U1025 ( .A(n384), .B(n767), .Y(n793) );
  XNOR2XL U1026 ( .A(n919), .B(A[16]), .Y(n798) );
  OAI22X2 U1027 ( .A0(n970), .A1(n798), .B0(n968), .B1(n769), .Y(n800) );
  CMPR32X1 U1028 ( .A(n776), .B(n775), .C(n774), .CO(n777), .S(n808) );
  XNOR2X1 U1029 ( .A(n924), .B(A[12]), .Y(n827) );
  XNOR2X1 U1030 ( .A(n1138), .B(A[4]), .Y(n797) );
  OAI22XL U1031 ( .A0(n1135), .A1(n823), .B0(n954), .B1(n788), .Y(n824) );
  XNOR2X1 U1032 ( .A(n908), .B(A[10]), .Y(n821) );
  OAI22XL U1033 ( .A0(n962), .A1(n821), .B0(n960), .B1(n792), .Y(n804) );
  ADDHXL U1034 ( .A(n794), .B(n793), .CO(n774), .S(n803) );
  OAI22X1 U1035 ( .A0(n240), .A1(n830), .B0(n795), .B1(n1085), .Y(n829) );
  XNOR2XL U1036 ( .A(n1156), .B(A[2]), .Y(n796) );
  NOR2XL U1037 ( .A(n384), .B(n796), .Y(n828) );
  OAI22X1 U1038 ( .A0(n970), .A1(n833), .B0(n968), .B1(n798), .Y(n868) );
  CMPR32X1 U1039 ( .A(n804), .B(n802), .C(n803), .CO(n805), .S(n845) );
  ADDFHX1 U1040 ( .A(n810), .B(n809), .CI(n808), .CO(n813), .S(n848) );
  NOR2XL U1041 ( .A(n815), .B(n814), .Y(mult_x_1_n262) );
  NAND2XL U1042 ( .A(n816), .B(n1291), .Y(n817) );
  ADDFHX1 U1043 ( .A(n820), .B(n819), .CI(n818), .CO(n814), .S(n852) );
  XNOR2X1 U1044 ( .A(n908), .B(A[9]), .Y(n865) );
  OAI22X1 U1045 ( .A0(n962), .A1(n865), .B0(n960), .B1(n821), .Y(n838) );
  OAI22X1 U1046 ( .A0(n976), .A1(n834), .B0(n9), .B1(n822), .Y(n837) );
  OAI22XL U1047 ( .A0(n1135), .A1(n863), .B0(n954), .B1(n823), .Y(n836) );
  XNOR2XL U1048 ( .A(n924), .B(A[11]), .Y(n864) );
  OAI22XL U1049 ( .A0(n979), .A1(n864), .B0(n757), .B1(n827), .Y(n841) );
  XNOR2X1 U1050 ( .A(n922), .B(A[6]), .Y(n879) );
  OAI22X1 U1051 ( .A0(n970), .A1(n874), .B0(n968), .B1(n833), .Y(n877) );
  CMPR32X1 U1052 ( .A(n838), .B(n837), .C(n836), .CO(n844), .S(n888) );
  CMPR32X1 U1053 ( .A(n841), .B(n840), .C(n839), .CO(n842), .S(n887) );
  NOR2XL U1054 ( .A(n852), .B(n851), .Y(mult_x_1_n265) );
  NAND2XL U1055 ( .A(n852), .B(n851), .Y(mult_x_1_n266) );
  INVXL U1056 ( .A(n1292), .Y(n856) );
  ADDFHX1 U1057 ( .A(n860), .B(n859), .CI(n858), .CO(n851), .S(n894) );
  NOR2XL U1058 ( .A(n384), .B(n862), .Y(n882) );
  OAI22XL U1059 ( .A0(n1135), .A1(n875), .B0(n954), .B1(n863), .Y(n881) );
  XNOR2XL U1060 ( .A(n924), .B(A[10]), .Y(n880) );
  OAI22XL U1061 ( .A0(n926), .A1(n880), .B0(n757), .B1(n864), .Y(n886) );
  OAI22XL U1062 ( .A0(n962), .A1(n873), .B0(n960), .B1(n865), .Y(n885) );
  ADDHXL U1063 ( .A(n867), .B(n866), .CO(n839), .S(n884) );
  XNOR2X1 U1064 ( .A(n1138), .B(A[1]), .Y(n910) );
  XNOR2X1 U1065 ( .A(n908), .B(A[7]), .Y(n909) );
  OAI22X2 U1066 ( .A0(n970), .A1(n920), .B0(n968), .B1(n874), .Y(n928) );
  XNOR2X1 U1067 ( .A(n650), .B(A[11]), .Y(n948) );
  XNOR2XL U1068 ( .A(n924), .B(A[9]), .Y(n925) );
  OAI22XL U1069 ( .A0(n926), .A1(n925), .B0(n757), .B1(n880), .Y(n930) );
  CMPR32X1 U1070 ( .A(n883), .B(n882), .C(n881), .CO(n903), .S(n946) );
  CMPR32X1 U1071 ( .A(n886), .B(n885), .C(n884), .CO(n902), .S(n945) );
  NOR2XL U1072 ( .A(n894), .B(n893), .Y(mult_x_1_n273) );
  NAND2XL U1073 ( .A(n894), .B(n893), .Y(mult_x_1_n274) );
  ADDFHX1 U1074 ( .A(n900), .B(n899), .CI(n898), .CO(n893), .S(n937) );
  CMPR32X1 U1075 ( .A(n903), .B(n902), .C(n901), .CO(n900), .S(n944) );
  OAI22X1 U1076 ( .A0(n240), .A1(n951), .B0(n906), .B1(n1085), .Y(n950) );
  XNOR2X1 U1077 ( .A(n1138), .B(A[0]), .Y(n911) );
  OAI22XL U1078 ( .A0(n1135), .A1(n953), .B0(n954), .B1(n912), .Y(n971) );
  OAI22XL U1079 ( .A0(n921), .A1(n967), .B0(n968), .B1(n920), .Y(n997) );
  OAI22X1 U1080 ( .A0(n966), .A1(n963), .B0(n964), .B1(n923), .Y(n996) );
  OAI22XL U1081 ( .A0(n926), .A1(n977), .B0(n757), .B1(n925), .Y(n995) );
  NOR2XL U1082 ( .A(n937), .B(n936), .Y(mult_x_1_n276) );
  NAND2XL U1083 ( .A(n937), .B(n936), .Y(mult_x_1_n277) );
  INVXL U1084 ( .A(n1296), .Y(n939) );
  NAND2X1 U1085 ( .A(n939), .B(n1297), .Y(n940) );
  XNOR2XL U1086 ( .A(n650), .B(A[10]), .Y(n974) );
  ADDFHX1 U1087 ( .A(n958), .B(n957), .CI(n956), .CO(n984), .S(n1011) );
  OAI22X1 U1088 ( .A0(n966), .A1(n965), .B0(n964), .B1(n963), .Y(n1008) );
  OAI22XL U1089 ( .A0(n976), .A1(n975), .B0(n9), .B1(n974), .Y(n1029) );
  OAI22XL U1090 ( .A0(n979), .A1(n978), .B0(n757), .B1(n977), .Y(n1028) );
  ADDHXL U1091 ( .A(n981), .B(n980), .CO(n1027), .S(n1032) );
  CMPR32X1 U1092 ( .A(n984), .B(n983), .C(n982), .CO(n943), .S(n989) );
  NOR2XL U1093 ( .A(n986), .B(n985), .Y(mult_x_1_n281) );
  NAND2XL U1094 ( .A(n986), .B(n985), .Y(mult_x_1_n282) );
  CMPR32X1 U1095 ( .A(n994), .B(n993), .C(n992), .CO(n982), .S(n1020) );
  CMPR32X1 U1096 ( .A(n1000), .B(n999), .C(n998), .CO(n1012), .S(n1034) );
  CMPR32X1 U1097 ( .A(n1003), .B(n1002), .C(n1001), .CO(n998), .S(n1040) );
  CMPR32X1 U1098 ( .A(n1006), .B(n1005), .C(n1004), .CO(n1039), .S(n1042) );
  NOR2XL U1099 ( .A(n1014), .B(n1013), .Y(mult_x_1_n286) );
  OAI21XL U1100 ( .A0(n1062), .A1(n1302), .B0(n1307), .Y(n1017) );
  INVXL U1101 ( .A(n1300), .Y(n1015) );
  NAND2XL U1102 ( .A(n1015), .B(n1301), .Y(n1016) );
  CMPR32X1 U1103 ( .A(n1023), .B(n1022), .C(n1021), .CO(n1010), .S(n1052) );
  CMPR32X1 U1104 ( .A(n1029), .B(n1028), .C(n1027), .CO(n1021), .S(n1045) );
  ADDFHX1 U1105 ( .A(n1032), .B(n1031), .CI(n1030), .CO(n1044), .S(n1049) );
  CMPR32X1 U1106 ( .A(n1035), .B(n1034), .C(n1033), .CO(n1019), .S(n1050) );
  NOR2XL U1107 ( .A(n1037), .B(n1036), .Y(mult_x_1_n292) );
  NAND2XL U1108 ( .A(n1037), .B(n1036), .Y(mult_x_1_n293) );
  CMPR32X1 U1109 ( .A(n1040), .B(n1039), .C(n1038), .CO(n1033), .S(n1055) );
  CMPR32X1 U1110 ( .A(n1043), .B(n1042), .C(n1041), .CO(n1054), .S(n1048) );
  ADDFHX1 U1111 ( .A(n1049), .B(n1048), .CI(n1047), .CO(n1056), .S(n285) );
  CMPR32X1 U1112 ( .A(n1052), .B(n1051), .C(n1050), .CO(n1036), .S(n1059) );
  OR2X2 U1113 ( .A(n1059), .B(n1058), .Y(n1091) );
  NAND2XL U1114 ( .A(n1091), .B(n1063), .Y(mult_x_1_n295) );
  INVXL U1115 ( .A(mult_x_1_n307), .Y(n1061) );
  NAND2XL U1116 ( .A(n1059), .B(n1058), .Y(n1090) );
  INVXL U1117 ( .A(n1090), .Y(n1060) );
  AOI21XL U1118 ( .A0(n1091), .A1(n1061), .B0(n1060), .Y(mult_x_1_n296) );
  NAND2XL U1119 ( .A(n1063), .B(mult_x_1_n307), .Y(mult_x_1_n84) );
  XOR2X1 U1120 ( .A(n1309), .B(n1305), .Y(PRODUCT[13]) );
  NAND2XL U1121 ( .A(n1065), .B(n1064), .Y(mult_x_1_n85) );
  XNOR2X1 U1122 ( .A(n1254), .B(n1306), .Y(PRODUCT[12]) );
  INVXL U1123 ( .A(n1066), .Y(mult_x_1_n321) );
  AOI21XL U1124 ( .A0(mult_x_1_n321), .A1(n6), .B0(n1067), .Y(mult_x_1_n316)
         );
  NAND2XL U1125 ( .A(n6), .B(n1068), .Y(mult_x_1_n86) );
  INVXL U1126 ( .A(n1069), .Y(n1071) );
  NAND2XL U1127 ( .A(n1071), .B(n1070), .Y(n1072) );
  AOI21XL U1128 ( .A0(n1172), .A1(n1170), .B0(n1074), .Y(n1078) );
  ADDFHX1 U1129 ( .A(n1081), .B(n1080), .CI(n1079), .CO(n748), .S(
        mult_x_1_n586) );
  INVXL U1130 ( .A(n1288), .Y(n1087) );
  NAND2XL U1131 ( .A(n1091), .B(n1090), .Y(mult_x_1_n83) );
  CMPR32X1 U1132 ( .A(n1096), .B(n1095), .C(n1094), .CO(n1111), .S(n1092) );
  XNOR2X1 U1133 ( .A(n1120), .B(A[24]), .Y(n1121) );
  OAI22XL U1134 ( .A0(n1161), .A1(n1103), .B0(n8), .B1(n1118), .Y(n1123) );
  CMPR32X1 U1135 ( .A(n1106), .B(n1105), .C(n1104), .CO(n1122), .S(n1096) );
  CMPR32X1 U1136 ( .A(n1109), .B(n1108), .C(n1107), .CO(n1112), .S(n1095) );
  CMPR32X1 U1137 ( .A(n1114), .B(n1113), .C(n1112), .CO(n1126), .S(n1110) );
  CMPR32X1 U1138 ( .A(n1117), .B(n1116), .C(n1115), .CO(n1145), .S(n1114) );
  OAI22XL U1139 ( .A0(n1161), .A1(n1118), .B0(n8), .B1(n1128), .Y(n1131) );
  OAI22X1 U1140 ( .A0(n1135), .A1(n1121), .B0(n1136), .B1(n1133), .Y(n1142) );
  CMPR32X1 U1141 ( .A(n1124), .B(n1123), .C(n1122), .CO(n1143), .S(n1113) );
  CMPR32X1 U1142 ( .A(n1131), .B(n1130), .C(n1129), .CO(n1147), .S(n1144) );
  CMPR32X1 U1143 ( .A(n1142), .B(n1141), .C(n1140), .CO(n1153), .S(n1146) );
  CMPR32X1 U1144 ( .A(n1145), .B(n1144), .C(n1143), .CO(n1152), .S(n1125) );
  CMPR32X1 U1145 ( .A(n1148), .B(n1147), .C(n1146), .CO(n1150), .S(n1151) );
  CMPR32X1 U1146 ( .A(n1155), .B(n1154), .C(n1153), .CO(n1166), .S(n1149) );
  XOR3X2 U1147 ( .A(n1164), .B(n1163), .C(n1162), .Y(n1165) );
  OAI21XL U1148 ( .A0(n1178), .A1(n1269), .B0(n1177), .Y(n1243) );
  AOI21XL U1149 ( .A0(n1210), .A1(n1183), .B0(n1182), .Y(n1184) );
  OAI21XL U1150 ( .A0(n1250), .A1(n1185), .B0(n1184), .Y(n1188) );
  OAI21XL U1151 ( .A0(n1201), .A1(n1199), .B0(n1200), .Y(n1194) );
  INVXL U1152 ( .A(n1190), .Y(n1192) );
  OAI21XL U1153 ( .A0(n1260), .A1(n1263), .B0(n1261), .Y(n1207) );
  AOI21XL U1154 ( .A0(n1210), .A1(n1203), .B0(n1207), .Y(n1195) );
  OAI21XL U1155 ( .A0(n1250), .A1(n1196), .B0(n1195), .Y(n1198) );
  AOI21XL U1156 ( .A0(n1210), .A1(n1209), .B0(n1208), .Y(n1211) );
  OAI21XL U1157 ( .A0(n1250), .A1(n1212), .B0(n1211), .Y(n1215) );
  XNOR2XL U1158 ( .A(n1226), .B(n1225), .Y(n1331) );
  XOR2XL U1159 ( .A(n1231), .B(n1230), .Y(n1332) );
  XOR2XL U1160 ( .A(n1236), .B(n1235), .Y(n1330) );
  OAI21XL U1161 ( .A0(n1240), .A1(n1256), .B0(n1257), .Y(n1241) );
  OAI21XL U1162 ( .A0(n1246), .A1(n1245), .B0(n1244), .Y(n1247) );
  OAI21XL U1163 ( .A0(n1250), .A1(n1249), .B0(n1248), .Y(n1251) );
  XNOR2XL U1164 ( .A(n1251), .B(n1255), .Y(PRODUCT[40]) );
endmodule


module FFT2048_DW02_mult_2_stage_J1_9 ( A, B, TC, CLK, PRODUCT );
  input [25:0] A;
  input [16:0] B;
  output [42:0] PRODUCT;
  input TC, CLK;
  wire   n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, mult_x_1_n665, mult_x_1_n650, mult_x_1_n649,
         mult_x_1_n634, mult_x_1_n633, mult_x_1_n618, mult_x_1_n617,
         mult_x_1_n602, mult_x_1_n601, mult_x_1_n586, mult_x_1_n569,
         mult_x_1_n554, mult_x_1_n553, mult_x_1_n538, mult_x_1_n537,
         mult_x_1_n522, mult_x_1_n521, mult_x_1_n508, mult_x_1_n507,
         mult_x_1_n321, mult_x_1_n316, mult_x_1_n309, mult_x_1_n307,
         mult_x_1_n306, mult_x_1_n296, mult_x_1_n295, mult_x_1_n293,
         mult_x_1_n292, mult_x_1_n287, mult_x_1_n286, mult_x_1_n282,
         mult_x_1_n281, mult_x_1_n245, mult_x_1_n244, mult_x_1_n195,
         mult_x_1_n194, mult_x_1_n184, mult_x_1_n183, mult_x_1_n177,
         mult_x_1_n176, mult_x_1_n170, mult_x_1_n169, mult_x_1_n161,
         mult_x_1_n160, mult_x_1_n152, mult_x_1_n151, mult_x_1_n137,
         mult_x_1_n136, mult_x_1_n130, mult_x_1_n129, mult_x_1_n121,
         mult_x_1_n120, mult_x_1_n110, mult_x_1_n109, mult_x_1_n86,
         mult_x_1_n85, mult_x_1_n84, mult_x_1_n83, mult_x_1_n58, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377;

  DFFHQXL mult_x_1_clk_r_REG12_S1 ( .D(mult_x_1_n183), .CK(CLK), .Q(n1338) );
  DFFHQXL mult_x_1_clk_r_REG16_S1 ( .D(mult_x_1_n169), .CK(CLK), .Q(n1334) );
  DFFHQXL mult_x_1_clk_r_REG18_S1 ( .D(mult_x_1_n160), .CK(CLK), .Q(n1332) );
  DFFHQXL mult_x_1_clk_r_REG20_S1 ( .D(mult_x_1_n151), .CK(CLK), .Q(n1330) );
  DFFHQX4 mult_x_1_clk_r_REG42_S1 ( .D(mult_x_1_n665), .CK(CLK), .Q(n1377) );
  DFFHQX4 mult_x_1_clk_r_REG41_S1 ( .D(mult_x_1_n650), .CK(CLK), .Q(n1376) );
  DFFHQX4 mult_x_1_clk_r_REG40_S1 ( .D(mult_x_1_n649), .CK(CLK), .Q(n1375) );
  DFFHQX4 mult_x_1_clk_r_REG39_S1 ( .D(mult_x_1_n634), .CK(CLK), .Q(n1374) );
  DFFHQX4 mult_x_1_clk_r_REG38_S1 ( .D(mult_x_1_n633), .CK(CLK), .Q(n1373) );
  DFFHQX4 mult_x_1_clk_r_REG37_S1 ( .D(mult_x_1_n618), .CK(CLK), .Q(n1372) );
  DFFHQX4 mult_x_1_clk_r_REG36_S1 ( .D(mult_x_1_n617), .CK(CLK), .Q(n1371) );
  DFFHQX4 mult_x_1_clk_r_REG35_S1 ( .D(mult_x_1_n602), .CK(CLK), .Q(n1370) );
  DFFHQX4 mult_x_1_clk_r_REG34_S1 ( .D(mult_x_1_n601), .CK(CLK), .Q(n1369) );
  DFFHQX4 mult_x_1_clk_r_REG30_S1 ( .D(mult_x_1_n569), .CK(CLK), .Q(n1367) );
  DFFHQX4 mult_x_1_clk_r_REG1_S1 ( .D(mult_x_1_n554), .CK(CLK), .Q(n1366) );
  DFFHQX4 mult_x_1_clk_r_REG3_S1 ( .D(mult_x_1_n538), .CK(CLK), .Q(n1364) );
  DFFHQX4 mult_x_1_clk_r_REG56_S1 ( .D(mult_x_1_n309), .CK(CLK), .Q(n1356) );
  DFFHQX4 mult_x_1_clk_r_REG50_S1 ( .D(mult_x_1_n296), .CK(CLK), .Q(n1355) );
  DFFHQX4 mult_x_1_clk_r_REG48_S1 ( .D(mult_x_1_n292), .CK(CLK), .Q(n1348) );
  DFFHQX1 mult_x_1_clk_r_REG54_S1 ( .D(mult_x_1_n306), .CK(CLK), .Q(n1318) );
  DFFHQX4 mult_x_1_clk_r_REG32_S1 ( .D(mult_x_1_n244), .CK(CLK), .Q(n1342) );
  DFFHQXL mult_x_1_clk_r_REG9_S1 ( .D(mult_x_1_n195), .CK(CLK), .Q(n1341) );
  DFFHQXL clk_r_REG63_S1 ( .D(n1393), .CK(CLK), .Q(PRODUCT[8]) );
  DFFHQXL mult_x_1_clk_r_REG49_S1 ( .D(mult_x_1_n83), .CK(CLK), .Q(n1351) );
  DFFHQXL mult_x_1_clk_r_REG21_S1 ( .D(mult_x_1_n137), .CK(CLK), .Q(n1329) );
  DFFHQXL mult_x_1_clk_r_REG17_S1 ( .D(mult_x_1_n161), .CK(CLK), .Q(n1333) );
  DFFHQXL mult_x_1_clk_r_REG19_S1 ( .D(mult_x_1_n152), .CK(CLK), .Q(n1331) );
  DFFHQXL mult_x_1_clk_r_REG60_S1 ( .D(mult_x_1_n321), .CK(CLK), .Q(n1320) );
  DFFHQXL clk_r_REG59_S1 ( .D(n1390), .CK(CLK), .Q(PRODUCT[11]) );
  DFFHQXL clk_r_REG61_S1 ( .D(n1391), .CK(CLK), .Q(PRODUCT[10]) );
  DFFHQXL mult_x_1_clk_r_REG31_S1 ( .D(mult_x_1_n245), .CK(CLK), .Q(n1343) );
  DFFHQXL clk_r_REG62_S1 ( .D(n1392), .CK(CLK), .Q(PRODUCT[9]) );
  DFFHQXL clk_r_REG71_S1 ( .D(n1401), .CK(CLK), .Q(PRODUCT[0]) );
  DFFHQXL mult_x_1_clk_r_REG28_S1 ( .D(mult_x_1_n109), .CK(CLK), .Q(n1322) );
  DFFHQXL mult_x_1_clk_r_REG22_S1 ( .D(mult_x_1_n136), .CK(CLK), .Q(n1328) );
  DFFHQXL clk_r_REG64_S1 ( .D(n1394), .CK(CLK), .Q(PRODUCT[7]) );
  DFFHQXL clk_r_REG65_S1 ( .D(n1395), .CK(CLK), .Q(PRODUCT[6]) );
  DFFHQXL clk_r_REG66_S1 ( .D(n1396), .CK(CLK), .Q(PRODUCT[5]) );
  DFFHQXL clk_r_REG67_S1 ( .D(n1397), .CK(CLK), .Q(PRODUCT[4]) );
  DFFHQXL clk_r_REG68_S1 ( .D(n1398), .CK(CLK), .Q(PRODUCT[3]) );
  DFFHQXL clk_r_REG69_S1 ( .D(n1399), .CK(CLK), .Q(PRODUCT[2]) );
  DFFHQXL clk_r_REG70_S1 ( .D(n1400), .CK(CLK), .Q(PRODUCT[1]) );
  DFFHQX2 mult_x_1_clk_r_REG5_S1 ( .D(mult_x_1_n522), .CK(CLK), .Q(n1362) );
  DFFHQX1 mult_x_1_clk_r_REG4_S1 ( .D(mult_x_1_n521), .CK(CLK), .Q(n1361) );
  DFFHQX1 mult_x_1_clk_r_REG58_S1 ( .D(mult_x_1_n316), .CK(CLK), .Q(n1357) );
  DFFHQXL mult_x_1_clk_r_REG57_S1 ( .D(mult_x_1_n86), .CK(CLK), .Q(n1354) );
  DFFHQX1 mult_x_1_clk_r_REG55_S1 ( .D(mult_x_1_n85), .CK(CLK), .Q(n1353) );
  DFFHQXL mult_x_1_clk_r_REG10_S1 ( .D(mult_x_1_n194), .CK(CLK), .Q(n1340) );
  DFFHQXL mult_x_1_clk_r_REG11_S1 ( .D(mult_x_1_n184), .CK(CLK), .Q(n1339) );
  DFFHQXL mult_x_1_clk_r_REG13_S1 ( .D(mult_x_1_n177), .CK(CLK), .Q(n1337) );
  DFFHQXL mult_x_1_clk_r_REG14_S1 ( .D(mult_x_1_n176), .CK(CLK), .Q(n1336) );
  DFFHQXL mult_x_1_clk_r_REG15_S1 ( .D(mult_x_1_n170), .CK(CLK), .Q(n1335) );
  DFFHQXL mult_x_1_clk_r_REG23_S1 ( .D(mult_x_1_n130), .CK(CLK), .Q(n1327) );
  DFFHQXL mult_x_1_clk_r_REG24_S1 ( .D(mult_x_1_n129), .CK(CLK), .Q(n1326) );
  DFFHQXL mult_x_1_clk_r_REG25_S1 ( .D(mult_x_1_n121), .CK(CLK), .Q(n1325) );
  DFFHQXL mult_x_1_clk_r_REG26_S1 ( .D(mult_x_1_n120), .CK(CLK), .Q(n1324) );
  DFFHQXL mult_x_1_clk_r_REG27_S1 ( .D(mult_x_1_n110), .CK(CLK), .Q(n1323) );
  DFFHQXL mult_x_1_clk_r_REG29_S1 ( .D(mult_x_1_n58), .CK(CLK), .Q(n1321) );
  DFFHQXL mult_x_1_clk_r_REG53_S1 ( .D(mult_x_1_n307), .CK(CLK), .Q(n1319) );
  DFFHQX1 mult_x_1_clk_r_REG52_S1 ( .D(mult_x_1_n84), .CK(CLK), .Q(n1352) );
  DFFHQX4 mult_x_1_clk_r_REG51_S1 ( .D(mult_x_1_n295), .CK(CLK), .Q(n1350) );
  DFFHQX2 mult_x_1_clk_r_REG44_S1 ( .D(mult_x_1_n281), .CK(CLK), .Q(n1344) );
  DFFHQX1 mult_x_1_clk_r_REG7_S1 ( .D(mult_x_1_n508), .CK(CLK), .Q(n1360) );
  DFFHQX1 mult_x_1_clk_r_REG47_S1 ( .D(mult_x_1_n293), .CK(CLK), .Q(n1349) );
  DFFHQX2 mult_x_1_clk_r_REG33_S1 ( .D(mult_x_1_n586), .CK(CLK), .Q(n1368) );
  DFFHQX1 mult_x_1_clk_r_REG46_S1 ( .D(mult_x_1_n286), .CK(CLK), .Q(n1346) );
  DFFHQX1 mult_x_1_clk_r_REG6_S1 ( .D(mult_x_1_n507), .CK(CLK), .Q(n1359) );
  DFFHQX1 mult_x_1_clk_r_REG43_S1 ( .D(mult_x_1_n282), .CK(CLK), .Q(n1345) );
  DFFHQX1 mult_x_1_clk_r_REG8_S1 ( .D(n62), .CK(CLK), .Q(n1358) );
  DFFHQX2 mult_x_1_clk_r_REG45_S1 ( .D(mult_x_1_n287), .CK(CLK), .Q(n1347) );
  DFFHQX2 mult_x_1_clk_r_REG2_S1 ( .D(mult_x_1_n537), .CK(CLK), .Q(n1363) );
  DFFHQX2 mult_x_1_clk_r_REG0_S1 ( .D(mult_x_1_n553), .CK(CLK), .Q(n1365) );
  OAI21XL U1 ( .A0(n118), .A1(n117), .B0(n116), .Y(n535) );
  ADDFHX1 U2 ( .A(n1143), .B(n1142), .CI(n1141), .CO(n1148), .S(n1150) );
  ADDFX2 U3 ( .A(n1004), .B(n1003), .CI(n1002), .CO(n982), .S(n1005) );
  ADDFHX1 U4 ( .A(n1146), .B(n1145), .CI(n1144), .CO(n1136), .S(n1147) );
  ADDFHX2 U5 ( .A(n980), .B(n979), .CI(n978), .CO(n958), .S(n981) );
  ADDFHX2 U6 ( .A(n726), .B(n725), .CI(n724), .CO(n1142), .S(n759) );
  CMPR32X1 U7 ( .A(n1107), .B(n1106), .C(n1105), .CO(n1110), .S(n1132) );
  ADDFHX1 U8 ( .A(n1125), .B(n1124), .CI(n1123), .CO(n1146), .S(n1141) );
  CMPR32X1 U9 ( .A(n499), .B(n498), .C(n497), .CO(n483), .S(n513) );
  CMPR32X1 U10 ( .A(n1059), .B(n1058), .C(n1057), .CO(n1068), .S(n1106) );
  ADDFX2 U11 ( .A(n424), .B(n423), .CI(n422), .CO(n445), .S(n481) );
  ADDFHX1 U12 ( .A(n623), .B(n622), .CI(n621), .CO(n614), .S(n639) );
  ADDFHX1 U13 ( .A(n1034), .B(n1033), .CI(n1032), .CO(n640), .S(n1064) );
  CMPR32X1 U14 ( .A(n819), .B(n818), .C(n817), .CO(n790), .S(n856) );
  ADDFHX1 U15 ( .A(n1084), .B(n1083), .CI(n1082), .CO(n1065), .S(n1103) );
  ADDFX2 U16 ( .A(n464), .B(n463), .CI(n462), .CO(n482), .S(n497) );
  CMPR32X1 U17 ( .A(n768), .B(n70), .C(n766), .CO(n784), .S(n818) );
  ADDFHX1 U18 ( .A(n886), .B(n885), .CI(n884), .CO(n888), .S(n285) );
  ADDFHX1 U19 ( .A(n410), .B(n409), .CI(n408), .CO(n388), .S(n443) );
  ADDFX2 U20 ( .A(n508), .B(n507), .CI(n506), .CO(n487), .S(n529) );
  CMPR32X1 U21 ( .A(n271), .B(n270), .C(n269), .CO(n885), .S(n281) );
  ADDFHX1 U22 ( .A(n843), .B(n842), .CI(n841), .CO(n838), .S(n1162) );
  NOR2X1 U23 ( .A(n212), .B(n213), .Y(n1255) );
  CLKBUFX8 U24 ( .A(n671), .Y(n1219) );
  CLKBUFX8 U25 ( .A(n266), .Y(n8) );
  CLKBUFX8 U26 ( .A(n417), .Y(n1046) );
  BUFX4 U27 ( .A(B[16]), .Y(n1044) );
  CLKINVX3 U28 ( .A(B[11]), .Y(n268) );
  XOR2X1 U29 ( .A(B[12]), .B(B[13]), .Y(n320) );
  BUFX4 U30 ( .A(n690), .Y(n1053) );
  XNOR2X1 U31 ( .A(B[12]), .B(B[11]), .Y(n567) );
  CLKINVX3 U32 ( .A(n402), .Y(n777) );
  BUFX4 U33 ( .A(n215), .Y(n1086) );
  BUFX4 U34 ( .A(n728), .Y(n1056) );
  BUFX4 U35 ( .A(n718), .Y(n1077) );
  BUFX3 U36 ( .A(n160), .Y(n6) );
  NAND2X1 U37 ( .A(n163), .B(n187), .Y(n690) );
  NAND2X1 U38 ( .A(n158), .B(n160), .Y(n718) );
  CLKINVX3 U39 ( .A(B[7]), .Y(n355) );
  XOR2X1 U40 ( .A(n52), .B(n503), .Y(PRODUCT[30]) );
  XNOR2X1 U41 ( .A(n546), .B(n545), .Y(PRODUCT[27]) );
  NOR2X1 U42 ( .A(n1370), .B(n1371), .Y(n315) );
  NAND2X1 U43 ( .A(n1377), .B(n1376), .Y(n661) );
  AND2X1 U44 ( .A(n438), .B(n309), .Y(n155) );
  XNOR2XL U45 ( .A(n746), .B(n1035), .Y(n807) );
  XNOR2XL U46 ( .A(n1281), .B(n1280), .Y(PRODUCT[39]) );
  XNOR2XL U47 ( .A(n774), .B(n1043), .Y(n174) );
  XNOR2XL U48 ( .A(n585), .B(n772), .Y(n278) );
  XNOR2XL U49 ( .A(n1036), .B(n1043), .Y(n833) );
  XNOR2XL U50 ( .A(n908), .B(n596), .Y(n929) );
  XNOR2XL U51 ( .A(n908), .B(n915), .Y(n605) );
  XNOR2XL U52 ( .A(n585), .B(n776), .Y(n744) );
  XNOR2XL U53 ( .A(n746), .B(A[14]), .Y(n731) );
  XNOR2XL U54 ( .A(n916), .B(n1201), .Y(n413) );
  XOR2XL U55 ( .A(n108), .B(n38), .Y(n171) );
  NAND2X2 U56 ( .A(n671), .B(n46), .Y(n673) );
  ADDFX2 U57 ( .A(n233), .B(n232), .CI(n231), .CO(n238), .S(n240) );
  BUFX3 U58 ( .A(n168), .Y(n9) );
  XNOR2XL U59 ( .A(n1185), .B(n1026), .Y(n946) );
  XNOR2XL U60 ( .A(n669), .B(n668), .Y(n1052) );
  XNOR2XL U61 ( .A(n746), .B(n732), .Y(n179) );
  ADDFX2 U62 ( .A(n877), .B(n876), .CI(n875), .CO(n853), .S(n1165) );
  ADDFX2 U63 ( .A(n965), .B(n964), .CI(n963), .CO(n1001), .S(n994) );
  ADDFX2 U64 ( .A(n825), .B(n824), .CI(n823), .CO(n817), .S(n861) );
  XOR2XL U65 ( .A(n19), .B(n616), .Y(n644) );
  AOI21XL U66 ( .A0(n874), .A1(n873), .B0(n872), .Y(n1172) );
  XOR2XL U67 ( .A(n1268), .B(n1267), .Y(n1395) );
  XNOR2XL U68 ( .A(n904), .B(n903), .Y(n1393) );
  CLKINVX2 U69 ( .A(n1348), .Y(n13) );
  NAND2XL U70 ( .A(n32), .B(n31), .Y(mult_x_1_n507) );
  NOR2XL U71 ( .A(n754), .B(n753), .Y(mult_x_1_n281) );
  XOR2X1 U72 ( .A(n61), .B(n1135), .Y(mult_x_1_n634) );
  OAI2BB1X1 U73 ( .A0N(n33), .A1N(n7), .B0(n957), .Y(n32) );
  NAND2X1 U74 ( .A(n285), .B(n284), .Y(n870) );
  INVX1 U75 ( .A(n1193), .Y(n1169) );
  NAND2X1 U76 ( .A(n958), .B(n959), .Y(n31) );
  NAND2X1 U77 ( .A(n244), .B(n243), .Y(n901) );
  OR2X2 U78 ( .A(n889), .B(n888), .Y(n887) );
  OAI21XL U79 ( .A0(n17), .A1(n16), .B0(n15), .Y(n857) );
  XOR2X1 U80 ( .A(n14), .B(n838), .Y(n859) );
  OAI21XL U81 ( .A0(n839), .A1(n840), .B0(n838), .Y(n15) );
  ADDFHX1 U82 ( .A(n1152), .B(n1151), .CI(n1150), .CO(mult_x_1_n665), .S(n754)
         );
  OAI2BB1XL U83 ( .A0N(n496), .A1N(n26), .B0(n24), .Y(n499) );
  OAI2BB1X1 U84 ( .A0N(n617), .A1N(n616), .B0(n18), .Y(n1013) );
  XOR2X1 U85 ( .A(n839), .B(n840), .Y(n14) );
  INVX1 U86 ( .A(n840), .Y(n17) );
  OAI21XL U87 ( .A0(n616), .A1(n617), .B0(n615), .Y(n18) );
  NAND2BXL U88 ( .AN(n496), .B(n29), .Y(n25) );
  INVXL U89 ( .A(n496), .Y(n27) );
  ADDFHX1 U90 ( .A(n584), .B(n583), .CI(n582), .CO(n1010), .S(n613) );
  NAND2XL U91 ( .A(n152), .B(n154), .Y(n351) );
  AOI2BB1X1 U92 ( .A0N(n457), .A1N(n5), .B0(n30), .Y(n29) );
  OAI2BB1XL U93 ( .A0N(n5), .A1N(n1205), .B0(n1204), .Y(n1212) );
  OAI22X1 U94 ( .A0(n1187), .A1(n797), .B0(n5), .B1(n796), .Y(n827) );
  OAI2BB1XL U95 ( .A0N(n1086), .A1N(n1088), .B0(n324), .Y(n330) );
  BUFX8 U96 ( .A(n625), .Y(n1088) );
  OAI22XL U97 ( .A0(n728), .A1(n165), .B0(n9), .B1(n219), .Y(n231) );
  NOR2BX1 U98 ( .AN(n1154), .B(n1086), .Y(n230) );
  XNOR2XL U99 ( .A(n774), .B(n1154), .Y(n186) );
  XOR2X1 U100 ( .A(n664), .B(n663), .Y(PRODUCT[19]) );
  XNOR2X1 U101 ( .A(n822), .B(n1351), .Y(PRODUCT[15]) );
  NAND2X1 U102 ( .A(n11), .B(n537), .Y(n538) );
  NAND2X1 U103 ( .A(n441), .B(n1337), .Y(n442) );
  NAND2X1 U104 ( .A(n474), .B(n1339), .Y(n475) );
  XOR2X1 U105 ( .A(n868), .B(n1352), .Y(PRODUCT[14]) );
  BUFX2 U106 ( .A(A[16]), .Y(n668) );
  XOR2X1 U107 ( .A(n957), .B(n23), .Y(mult_x_1_n508) );
  NAND2X1 U108 ( .A(n132), .B(n131), .Y(n785) );
  INVX1 U109 ( .A(n901), .Y(n896) );
  NAND2X1 U110 ( .A(n262), .B(n261), .Y(n891) );
  NOR2X1 U111 ( .A(n863), .B(n862), .Y(mult_x_1_n306) );
  NAND2X1 U112 ( .A(n863), .B(n862), .Y(mult_x_1_n307) );
  NAND2X1 U113 ( .A(n213), .B(n212), .Y(n1256) );
  NAND2X1 U114 ( .A(n889), .B(n888), .Y(n1193) );
  ADDFHX2 U115 ( .A(n1134), .B(n1133), .CI(n1132), .CO(n1112), .S(n1135) );
  ADDFHX1 U116 ( .A(n861), .B(n860), .CI(n859), .CO(n864), .S(n863) );
  INVX1 U117 ( .A(n959), .Y(n7) );
  ADDFHX1 U118 ( .A(n1013), .B(n1012), .CI(n1011), .CO(n1018), .S(n1021) );
  ADDFHX1 U119 ( .A(n614), .B(n613), .CI(n612), .CO(n1022), .S(n645) );
  INVXL U120 ( .A(n245), .Y(n90) );
  XOR2X2 U121 ( .A(n252), .B(n97), .Y(n36) );
  ADDFHX1 U122 ( .A(n701), .B(n700), .CI(n699), .CO(n1143), .S(n751) );
  INVXL U123 ( .A(n1064), .Y(n88) );
  XOR2X1 U124 ( .A(n615), .B(n617), .Y(n19) );
  NAND2XL U125 ( .A(n495), .B(n25), .Y(n24) );
  XOR2X1 U126 ( .A(n28), .B(n27), .Y(n525) );
  ADDFHX1 U127 ( .A(n989), .B(n988), .CI(n987), .CO(n977), .S(n997) );
  OAI22X1 U128 ( .A0(n1088), .A1(n216), .B0(n1086), .B1(n254), .Y(n256) );
  INVX4 U129 ( .A(n1088), .Y(n99) );
  XNOR2X1 U130 ( .A(n1246), .B(n1245), .Y(PRODUCT[36]) );
  XNOR2X1 U131 ( .A(n1253), .B(n1252), .Y(PRODUCT[37]) );
  XNOR2X1 U132 ( .A(n1263), .B(n1262), .Y(PRODUCT[38]) );
  INVXL U133 ( .A(n251), .Y(n37) );
  OAI22XL U134 ( .A0(n1056), .A1(n1054), .B0(n9), .B1(n631), .Y(n1057) );
  NAND2XL U135 ( .A(n151), .B(n1303), .Y(n400) );
  NOR2BX1 U136 ( .AN(n1154), .B(n8), .Y(n274) );
  OAI22XL U137 ( .A0(n1053), .A1(n249), .B0(n1051), .B1(n280), .Y(n275) );
  OR2XL U138 ( .A(n183), .B(n182), .Y(n1310) );
  XOR2X1 U139 ( .A(n560), .B(n56), .Y(PRODUCT[25]) );
  CLKBUFX8 U140 ( .A(n567), .Y(n5) );
  XOR2X1 U141 ( .A(n1159), .B(n1158), .Y(PRODUCT[21]) );
  OAI2BB1XL U142 ( .A0N(n144), .A1N(n561), .B0(n649), .Y(n156) );
  NOR2X1 U143 ( .A(n1296), .B(n1242), .Y(n1270) );
  XNOR2X1 U144 ( .A(n788), .B(n787), .Y(PRODUCT[16]) );
  INVX1 U145 ( .A(n536), .Y(n11) );
  BUFX2 U146 ( .A(A[18]), .Y(n719) );
  BUFX2 U147 ( .A(A[3]), .Y(n1043) );
  INVX1 U148 ( .A(n1332), .Y(n1235) );
  INVX1 U149 ( .A(n895), .Y(n904) );
  XNOR2X1 U150 ( .A(n1259), .B(n1258), .Y(n1394) );
  NAND2XL U151 ( .A(n869), .B(mult_x_1_n307), .Y(mult_x_1_n84) );
  INVXL U152 ( .A(mult_x_1_n307), .Y(n867) );
  NAND2X1 U153 ( .A(n865), .B(n864), .Y(n1155) );
  NAND2XL U154 ( .A(n898), .B(n897), .Y(n899) );
  NAND2XL U155 ( .A(n125), .B(n124), .Y(mult_x_1_n633) );
  ADDFHX1 U156 ( .A(n1007), .B(n1006), .CI(n1005), .CO(mult_x_1_n537), .S(
        mult_x_1_n538) );
  NAND2XL U157 ( .A(n133), .B(n789), .Y(n132) );
  NAND2XL U158 ( .A(n1136), .B(n1137), .Y(n124) );
  INVXL U159 ( .A(n906), .Y(n117) );
  NOR2X1 U160 ( .A(n1255), .B(n1264), .Y(n214) );
  NAND2BX2 U161 ( .AN(n246), .B(n90), .Y(n898) );
  INVX1 U162 ( .A(n22), .Y(n23) );
  ADDFHX1 U163 ( .A(n1019), .B(n1018), .CI(n1017), .CO(mult_x_1_n553), .S(
        mult_x_1_n554) );
  NAND2XL U164 ( .A(n790), .B(n791), .Y(n131) );
  INVXL U165 ( .A(n243), .Y(n94) );
  ADDFHX2 U166 ( .A(n515), .B(n514), .CI(n513), .CO(n531), .S(n906) );
  INVX1 U167 ( .A(n958), .Y(n33) );
  INVXL U168 ( .A(n982), .Y(n122) );
  INVXL U169 ( .A(n758), .Y(n103) );
  NAND2X1 U170 ( .A(n211), .B(n210), .Y(n1265) );
  XOR2X1 U171 ( .A(n250), .B(n35), .Y(n258) );
  INVXL U172 ( .A(n907), .Y(n118) );
  ADDFHX1 U173 ( .A(n1165), .B(n1164), .CI(n1163), .CO(n1166), .S(n889) );
  OAI2BB1XL U174 ( .A0N(n86), .A1N(n1063), .B0(n85), .Y(n1074) );
  OAI2BB1XL U175 ( .A0N(n111), .A1N(n387), .B0(n110), .Y(n433) );
  NAND2XL U176 ( .A(n88), .B(n87), .Y(n86) );
  ADDFHX1 U177 ( .A(n611), .B(n68), .CI(n609), .CO(n612), .S(n641) );
  INVXL U178 ( .A(n759), .Y(n104) );
  INVXL U179 ( .A(n791), .Y(n134) );
  OR2XL U180 ( .A(n1224), .B(n1223), .Y(n1226) );
  XOR2X1 U181 ( .A(n37), .B(n36), .Y(n35) );
  ADDFHX1 U182 ( .A(n173), .B(n171), .CI(n172), .CO(n212), .S(n211) );
  INVXL U183 ( .A(n63), .Y(n64) );
  NAND2XL U184 ( .A(n140), .B(n139), .Y(n484) );
  XOR2X1 U185 ( .A(n100), .B(n486), .Y(n515) );
  OR2XL U186 ( .A(n388), .B(n389), .Y(n111) );
  INVX1 U187 ( .A(n839), .Y(n16) );
  ADDFHX2 U188 ( .A(n640), .B(n639), .CI(n638), .CO(n1025), .S(n1070) );
  NOR2BX1 U189 ( .AN(n252), .B(n97), .Y(n271) );
  ADDFHX2 U190 ( .A(n974), .B(n973), .CI(n972), .CO(n980), .S(n1003) );
  ADDFHX1 U191 ( .A(n1119), .B(n1118), .CI(n1117), .CO(n1104), .S(n1127) );
  NAND2BXL U192 ( .AN(n837), .B(n43), .Y(n42) );
  ADDFHX1 U193 ( .A(n277), .B(n276), .CI(n275), .CO(n879), .S(n283) );
  ADDFHX1 U194 ( .A(n494), .B(n493), .CI(n492), .CO(n486), .S(n526) );
  INVXL U195 ( .A(n29), .Y(n26) );
  ADDFHX1 U196 ( .A(n742), .B(n741), .CI(n740), .CO(n734), .S(n793) );
  OAI2BB1XL U197 ( .A0N(n6), .A1N(n1077), .B0(n357), .Y(n384) );
  NAND2BXL U198 ( .AN(n175), .B(n40), .Y(n39) );
  INVXL U199 ( .A(n45), .Y(n43) );
  NAND2XL U200 ( .A(n45), .B(n837), .Y(n41) );
  OR2X2 U201 ( .A(n200), .B(n199), .Y(n198) );
  OAI2BB1XL U202 ( .A0N(n1051), .A1N(n1053), .B0(n452), .Y(n506) );
  XNOR2X2 U203 ( .A(n476), .B(n475), .Y(PRODUCT[31]) );
  INVXL U204 ( .A(n1056), .Y(n40) );
  NAND2BXL U205 ( .AN(n109), .B(n107), .Y(n106) );
  AND2XL U206 ( .A(n1285), .B(n1284), .Y(n1400) );
  NAND2BXL U207 ( .AN(n349), .B(n153), .Y(n152) );
  XNOR2XL U208 ( .A(n1044), .B(A[19]), .Y(n319) );
  XNOR2XL U209 ( .A(n1044), .B(n668), .Y(n354) );
  XNOR2XL U210 ( .A(n1044), .B(A[24]), .Y(n1215) );
  XNOR2XL U211 ( .A(n1210), .B(A[24]), .Y(n1211) );
  XNOR2XL U212 ( .A(n1210), .B(A[25]), .Y(n1216) );
  INVXL U213 ( .A(n1307), .Y(n153) );
  XNOR2XL U214 ( .A(n1044), .B(n1208), .Y(n1209) );
  OR2XL U215 ( .A(n1283), .B(n1282), .Y(n1285) );
  OAI22X1 U216 ( .A0(n180), .A1(n627), .B0(n572), .B1(n1153), .Y(n626) );
  BUFX3 U217 ( .A(n180), .Y(n808) );
  NAND2X1 U218 ( .A(B[1]), .B(n1040), .Y(n180) );
  AND2XL U219 ( .A(n559), .B(n558), .Y(n56) );
  INVXL U220 ( .A(n537), .Y(n53) );
  INVXL U221 ( .A(n1026), .Y(n21) );
  NAND2X1 U222 ( .A(n12), .B(n13), .Y(n49) );
  INVXL U223 ( .A(n314), .Y(n149) );
  NOR2X1 U224 ( .A(n551), .B(n547), .Y(n302) );
  INVXL U225 ( .A(n303), .Y(n145) );
  INVX1 U226 ( .A(B[0]), .Y(n1040) );
  INVXL U227 ( .A(n1346), .Y(n755) );
  INVXL U228 ( .A(n1154), .Y(n10) );
  BUFX2 U229 ( .A(A[1]), .Y(n732) );
  BUFX2 U230 ( .A(A[7]), .Y(n1030) );
  BUFX2 U231 ( .A(A[8]), .Y(n776) );
  BUFX2 U232 ( .A(A[4]), .Y(n772) );
  BUFX2 U233 ( .A(A[5]), .Y(n1028) );
  BUFX2 U234 ( .A(A[9]), .Y(n920) );
  BUFX2 U235 ( .A(A[21]), .Y(n1183) );
  BUFX2 U236 ( .A(A[20]), .Y(n596) );
  BUFX2 U237 ( .A(A[17]), .Y(n915) );
  BUFX2 U238 ( .A(A[11]), .Y(n1035) );
  BUFX2 U239 ( .A(A[12]), .Y(n745) );
  BUFX2 U240 ( .A(A[22]), .Y(n1201) );
  BUFX2 U241 ( .A(A[13]), .Y(n1026) );
  BUFX2 U242 ( .A(A[23]), .Y(n1208) );
  INVX1 U243 ( .A(n1355), .Y(n12) );
  OAI22X1 U244 ( .A0(n1218), .A1(n587), .B0(n1219), .B1(n945), .Y(n985) );
  AOI21X2 U245 ( .A0(n130), .A1(n653), .B0(n128), .Y(n127) );
  NAND2BX1 U246 ( .AN(n1296), .B(n78), .Y(n151) );
  NOR2BX1 U247 ( .AN(n1154), .B(n1219), .Y(n771) );
  AOI21X1 U248 ( .A0(n867), .A1(n1156), .B0(n866), .Y(mult_x_1_n296) );
  NOR2X1 U249 ( .A(n96), .B(n95), .Y(n895) );
  OAI22X1 U250 ( .A0(n1049), .A1(n695), .B0(n8), .B1(n686), .Y(n713) );
  NAND3X1 U251 ( .A(n48), .B(n51), .C(n1356), .Y(n50) );
  NOR2X1 U252 ( .A(n1367), .B(n1366), .Y(n547) );
  NOR2X1 U253 ( .A(n1365), .B(n1364), .Y(n551) );
  CLKINVX3 U254 ( .A(n78), .Y(n1307) );
  NAND3X2 U255 ( .A(n141), .B(n142), .C(n54), .Y(n78) );
  OAI22X1 U256 ( .A0(n574), .A1(n1049), .B0(n8), .B1(n20), .Y(n594) );
  OAI22X1 U257 ( .A0(n925), .A1(n8), .B0(n1049), .B1(n20), .Y(n965) );
  XOR2X1 U258 ( .A(n799), .B(n21), .Y(n20) );
  XOR2X1 U259 ( .A(n958), .B(n7), .Y(n22) );
  XOR2X1 U260 ( .A(n495), .B(n29), .Y(n28) );
  NOR2X1 U261 ( .A(n504), .B(n1205), .Y(n30) );
  NAND2X1 U262 ( .A(n898), .B(n902), .Y(n93) );
  OAI2BB2X1 U263 ( .B0(n36), .B1(n37), .A0N(n34), .A1N(n250), .Y(n282) );
  NAND2BXL U264 ( .AN(n251), .B(n36), .Y(n34) );
  OAI2BB1X1 U265 ( .A0N(n38), .A1N(n106), .B0(n105), .Y(n241) );
  OAI21XL U266 ( .A0(n165), .A1(n9), .B0(n39), .Y(n38) );
  NOR2X1 U267 ( .A(n211), .B(n210), .Y(n1264) );
  OAI2BB1X1 U268 ( .A0N(n836), .A1N(n42), .B0(n41), .Y(n842) );
  XNOR2X1 U269 ( .A(n836), .B(n44), .Y(n875) );
  XNOR2X1 U270 ( .A(n837), .B(n45), .Y(n44) );
  NOR2X1 U271 ( .A(n5), .B(n10), .Y(n45) );
  XNOR2X2 U272 ( .A(B[14]), .B(n47), .Y(n46) );
  INVX1 U273 ( .A(B[15]), .Y(n47) );
  XNOR2X4 U274 ( .A(B[14]), .B(B[13]), .Y(n671) );
  INVX1 U275 ( .A(n1350), .Y(n48) );
  CLKINVX3 U276 ( .A(n119), .Y(n296) );
  NAND3X2 U277 ( .A(n50), .B(n1349), .C(n49), .Y(n119) );
  CLKINVX2 U278 ( .A(n1348), .Y(n51) );
  CLKINVX2 U279 ( .A(B[3]), .Y(n189) );
  AOI21X1 U280 ( .A0(n78), .A1(n11), .B0(n53), .Y(n52) );
  OAI21X1 U281 ( .A0(n315), .A1(n314), .B0(n316), .Y(n563) );
  NAND2X2 U282 ( .A(n1372), .B(n1373), .Y(n314) );
  XOR2X1 U283 ( .A(B[10]), .B(B[11]), .Y(n120) );
  OAI22X1 U284 ( .A0(n1088), .A1(n737), .B0(n1086), .B1(n683), .Y(n742) );
  OAI22X1 U285 ( .A0(n1088), .A1(n683), .B0(n1086), .B1(n682), .Y(n693) );
  XNOR2X1 U286 ( .A(n1036), .B(n1035), .Y(n1085) );
  XNOR2X1 U287 ( .A(n1036), .B(n920), .Y(n714) );
  XNOR2X1 U288 ( .A(n1036), .B(n776), .Y(n682) );
  ADDFX2 U289 ( .A(n941), .B(n940), .CI(n939), .CO(n959), .S(n979) );
  XNOR2X1 U290 ( .A(n923), .B(n922), .Y(n951) );
  NOR2X1 U291 ( .A(n1046), .B(n921), .Y(n935) );
  XNOR2X1 U292 ( .A(n1210), .B(A[14]), .Y(n454) );
  XNOR2X1 U293 ( .A(n1210), .B(n745), .Y(n512) );
  OAI22X1 U294 ( .A0(n1077), .A1(n511), .B0(n6), .B1(n489), .Y(n914) );
  XNOR2X1 U295 ( .A(n585), .B(n1183), .Y(n489) );
  OAI22X1 U296 ( .A0(n1049), .A1(n925), .B0(n8), .B1(n924), .Y(n968) );
  OAI22X1 U297 ( .A0(n1218), .A1(n512), .B0(n1219), .B1(n491), .Y(n912) );
  XNOR2X1 U298 ( .A(n1210), .B(n1026), .Y(n491) );
  OAI22X2 U299 ( .A0(n1218), .A1(n944), .B0(n1219), .B1(n512), .Y(n922) );
  BUFX1 U300 ( .A(A[2]), .Y(n798) );
  NAND2X1 U301 ( .A(n147), .B(n556), .Y(n141) );
  NAND3X1 U302 ( .A(n144), .B(n157), .C(n147), .Y(n142) );
  XNOR2X1 U303 ( .A(B[8]), .B(B[7]), .Y(n215) );
  NAND2X2 U304 ( .A(n215), .B(n135), .Y(n625) );
  XOR2X1 U305 ( .A(B[9]), .B(B[8]), .Y(n135) );
  OAI22X1 U306 ( .A0(n1077), .A1(n411), .B0(n6), .B1(n356), .Y(n385) );
  NAND2X2 U307 ( .A(n320), .B(n567), .Y(n1205) );
  INVXL U308 ( .A(n1333), .Y(n1238) );
  NAND2XL U309 ( .A(n1235), .B(n1237), .Y(n1240) );
  INVXL U310 ( .A(n1157), .Y(n150) );
  INVXL U311 ( .A(n1330), .Y(n1237) );
  XNOR2XL U312 ( .A(n746), .B(A[6]), .Y(n161) );
  NOR2XL U313 ( .A(n1240), .B(n1334), .Y(n1295) );
  NOR2XL U314 ( .A(n1294), .B(n1322), .Y(n1299) );
  INVXL U315 ( .A(n1324), .Y(n1272) );
  OAI21XL U316 ( .A0(n1303), .A1(n1242), .B0(n1241), .Y(n1276) );
  INVXL U317 ( .A(n1300), .Y(n1241) );
  XNOR2X1 U318 ( .A(n659), .B(n658), .Y(PRODUCT[20]) );
  OAI21XL U319 ( .A0(n664), .A1(n660), .B0(n661), .Y(n659) );
  XNOR2X1 U320 ( .A(n146), .B(n442), .Y(PRODUCT[32]) );
  XNOR2X1 U321 ( .A(n313), .B(n312), .Y(PRODUCT[34]) );
  NAND2XL U322 ( .A(n1235), .B(n1333), .Y(n312) );
  CMPR32X1 U323 ( .A(n461), .B(n460), .C(n459), .CO(n446), .S(n498) );
  OAI22XL U324 ( .A0(n1205), .A1(n457), .B0(n5), .B1(n416), .Y(n461) );
  XNOR2XL U325 ( .A(n1210), .B(n776), .Y(n569) );
  XNOR2XL U326 ( .A(n585), .B(n668), .Y(n568) );
  XNOR2XL U327 ( .A(n777), .B(n1026), .Y(n715) );
  NOR2X1 U328 ( .A(n1046), .B(n721), .Y(n1091) );
  XNOR2X1 U329 ( .A(n1185), .B(A[6]), .Y(n1081) );
  ADDFX2 U330 ( .A(n386), .B(n385), .CI(n384), .CO(n367), .S(n429) );
  NOR2XL U331 ( .A(n1046), .B(n354), .Y(n386) );
  OAI22XL U332 ( .A0(n1187), .A1(n376), .B0(n5), .B1(n363), .Y(n381) );
  OAI22XL U333 ( .A0(n1088), .A1(n377), .B0(n1086), .B1(n361), .Y(n383) );
  NAND2XL U334 ( .A(n1295), .B(n1299), .Y(n1302) );
  NOR2XL U335 ( .A(n1046), .B(n1202), .Y(n1213) );
  INVXL U336 ( .A(n1203), .Y(n1204) );
  OAI22XL U337 ( .A0(n1056), .A1(n597), .B0(n9), .B1(n929), .Y(n963) );
  INVXL U338 ( .A(n385), .Y(n408) );
  NAND2XL U339 ( .A(n74), .B(n75), .Y(n72) );
  NAND2XL U340 ( .A(n76), .B(n77), .Y(n73) );
  INVXL U341 ( .A(n375), .Y(n74) );
  OAI22XL U342 ( .A0(n1049), .A1(n414), .B0(n8), .B1(n380), .Y(n405) );
  NOR2XL U343 ( .A(n1046), .B(n378), .Y(n407) );
  OAI22XL U344 ( .A0(n1218), .A1(n412), .B0(n1219), .B1(n379), .Y(n406) );
  OAI22XL U345 ( .A0(n1218), .A1(n1211), .B0(n1219), .B1(n1216), .Y(n1222) );
  OAI22XL U346 ( .A0(n1187), .A1(n1031), .B0(n5), .B1(n620), .Y(n1032) );
  OAI22X1 U347 ( .A0(n1077), .A1(n1027), .B0(n6), .B1(n618), .Y(n1034) );
  OAI22X2 U348 ( .A0(n1218), .A1(n1029), .B0(n1219), .B1(n619), .Y(n1033) );
  OAI22X1 U349 ( .A0(n1077), .A1(n1075), .B0(n6), .B1(n1027), .Y(n1084) );
  OAI22X2 U350 ( .A0(n1218), .A1(n1078), .B0(n1219), .B1(n1029), .Y(n1083) );
  ADDFX2 U351 ( .A(n1062), .B(n1061), .CI(n1060), .CO(n1063), .S(n1105) );
  NAND2XL U352 ( .A(n191), .B(n190), .Y(n1287) );
  AOI21XL U353 ( .A0(n1310), .A1(n1311), .B0(n184), .Y(n1289) );
  INVXL U354 ( .A(n1309), .Y(n184) );
  NAND2XL U355 ( .A(n200), .B(n199), .Y(n1291) );
  NOR2X1 U356 ( .A(n1346), .B(n1344), .Y(n654) );
  NOR2X1 U357 ( .A(n1369), .B(n1368), .Y(n562) );
  NOR2X1 U358 ( .A(n562), .B(n1342), .Y(n289) );
  NOR2XL U359 ( .A(n1328), .B(n1326), .Y(n1269) );
  NAND2X1 U360 ( .A(n81), .B(n79), .Y(n556) );
  NOR2BX1 U361 ( .AN(n1343), .B(n80), .Y(n79) );
  NAND2X1 U362 ( .A(n563), .B(n289), .Y(n81) );
  NOR2X1 U363 ( .A(n651), .B(n1342), .Y(n80) );
  AOI21X1 U364 ( .A0(n119), .A1(n654), .B0(n653), .Y(n664) );
  NAND2X1 U365 ( .A(n1371), .B(n1370), .Y(n316) );
  NAND2X1 U366 ( .A(n1368), .B(n1369), .Y(n651) );
  INVXL U367 ( .A(n562), .Y(n652) );
  NAND3BX1 U368 ( .AN(n650), .B(n144), .C(n652), .Y(n138) );
  INVXL U369 ( .A(n561), .Y(n650) );
  INVXL U370 ( .A(n1342), .Y(n566) );
  INVXL U371 ( .A(n556), .Y(n307) );
  NAND2X1 U372 ( .A(n1366), .B(n1367), .Y(n558) );
  INVXL U373 ( .A(n547), .Y(n559) );
  AOI21XL U374 ( .A0(n556), .A1(n559), .B0(n548), .Y(n549) );
  INVXL U375 ( .A(n558), .Y(n548) );
  NAND2XL U376 ( .A(n1364), .B(n1365), .Y(n552) );
  INVXL U377 ( .A(n551), .Y(n553) );
  XNOR2XL U378 ( .A(n585), .B(n798), .Y(n226) );
  XNOR2XL U379 ( .A(n777), .B(n776), .Y(n815) );
  XNOR2XL U380 ( .A(n777), .B(n920), .Y(n778) );
  XNOR2XL U381 ( .A(n777), .B(n1030), .Y(n816) );
  NAND2BXL U382 ( .AN(n1154), .B(n799), .Y(n267) );
  XNOR2XL U383 ( .A(n746), .B(A[15]), .Y(n675) );
  XNOR2XL U384 ( .A(n777), .B(n1035), .Y(n727) );
  XNOR2XL U385 ( .A(n777), .B(A[25]), .Y(n403) );
  XNOR2X1 U386 ( .A(n585), .B(n732), .Y(n227) );
  NAND2XL U387 ( .A(n1248), .B(n1329), .Y(n1245) );
  AOI21XL U388 ( .A0(n1276), .A1(n1269), .B0(n1273), .Y(n1260) );
  NAND2XL U389 ( .A(n1270), .B(n1269), .Y(n1261) );
  INVXL U390 ( .A(n1294), .Y(n1275) );
  NAND2XL U391 ( .A(n1251), .B(n1327), .Y(n1252) );
  NAND2XL U392 ( .A(n1237), .B(n1331), .Y(n350) );
  OAI22XL U393 ( .A0(n690), .A1(n222), .B0(n1051), .B1(n249), .Y(n251) );
  INVXL U394 ( .A(n1185), .Y(n749) );
  INVXL U395 ( .A(n337), .Y(n338) );
  XNOR2XL U396 ( .A(n916), .B(n1183), .Y(n449) );
  OAI22XL U397 ( .A0(n1049), .A1(n510), .B0(n8), .B1(n458), .Y(n495) );
  OAI22XL U398 ( .A0(n1088), .A1(n509), .B0(n1086), .B1(n456), .Y(n496) );
  XNOR2XL U399 ( .A(n916), .B(A[19]), .Y(n509) );
  INVXL U400 ( .A(n918), .Y(n518) );
  XNOR2X1 U401 ( .A(n799), .B(A[14]), .Y(n925) );
  XNOR2X1 U402 ( .A(n1210), .B(n772), .Y(n1079) );
  XNOR2X1 U403 ( .A(n1210), .B(n1043), .Y(n667) );
  NOR2XL U404 ( .A(n1046), .B(n321), .Y(n332) );
  INVXL U405 ( .A(n323), .Y(n324) );
  OAI22XL U406 ( .A0(n1049), .A1(n329), .B0(n8), .B1(n327), .Y(n333) );
  OAI22XL U407 ( .A0(n1187), .A1(n352), .B0(n5), .B1(n326), .Y(n334) );
  OAI22XL U408 ( .A0(n1218), .A1(n328), .B0(n1219), .B1(n325), .Y(n335) );
  INVXL U409 ( .A(n1049), .Y(n77) );
  OAI22XL U410 ( .A0(n1049), .A1(n421), .B0(n8), .B1(n414), .Y(n448) );
  AOI21XL U411 ( .A0(n1300), .A1(n1299), .B0(n1298), .Y(n1301) );
  AOI21XL U412 ( .A0(n1276), .A1(n1275), .B0(n1274), .Y(n1277) );
  INVXL U413 ( .A(n1297), .Y(n1274) );
  NAND2XL U414 ( .A(n1270), .B(n1275), .Y(n1278) );
  INVXL U415 ( .A(n1322), .Y(n1279) );
  OAI22XL U416 ( .A0(n1187), .A1(n339), .B0(n5), .B1(n1186), .Y(n1190) );
  OAI22XL U417 ( .A0(n1218), .A1(n340), .B0(n1219), .B1(n1182), .Y(n1189) );
  NOR2XL U418 ( .A(n1046), .B(n1184), .Y(n1199) );
  INVXL U419 ( .A(n1214), .Y(n1198) );
  OAI22XL U420 ( .A0(n1218), .A1(n1182), .B0(n1219), .B1(n1197), .Y(n1200) );
  INVX1 U421 ( .A(n897), .Y(n91) );
  INVXL U422 ( .A(n451), .Y(n452) );
  OAI21XL U423 ( .A0(n1086), .A1(n449), .B0(n101), .Y(n488) );
  OR2X2 U424 ( .A(n456), .B(n1088), .Y(n101) );
  OAI22XL U425 ( .A0(n1077), .A1(n489), .B0(n6), .B1(n455), .Y(n492) );
  OAI22X1 U426 ( .A0(n1218), .A1(n491), .B0(n1219), .B1(n454), .Y(n493) );
  CMPR32X1 U427 ( .A(n914), .B(n913), .C(n912), .CO(n527), .S(n940) );
  OAI22XL U428 ( .A0(n1053), .A1(n575), .B0(n1051), .B1(n595), .Y(n593) );
  OAI22XL U429 ( .A0(n1187), .A1(n588), .B0(n5), .B1(n947), .Y(n984) );
  OAI22X1 U430 ( .A0(n1077), .A1(n586), .B0(n6), .B1(n943), .Y(n986) );
  OAI22XL U431 ( .A0(n1187), .A1(n570), .B0(n5), .B1(n588), .Y(n582) );
  OAI22X1 U432 ( .A0(n1077), .A1(n568), .B0(n6), .B1(n586), .Y(n584) );
  OAI22X1 U433 ( .A0(n1218), .A1(n569), .B0(n1219), .B1(n587), .Y(n583) );
  XNOR2X1 U434 ( .A(n1210), .B(n1028), .Y(n1078) );
  XNOR2XL U435 ( .A(n585), .B(n1026), .Y(n1075) );
  OAI22X1 U436 ( .A0(n1056), .A1(n715), .B0(n9), .B1(n1055), .Y(n1115) );
  OAI22X1 U437 ( .A0(n1088), .A1(n714), .B0(n1086), .B1(n1087), .Y(n1116) );
  ADDFX2 U438 ( .A(n1122), .B(n1121), .CI(n1120), .CO(n1126), .S(n1123) );
  XOR2X1 U439 ( .A(n387), .B(n112), .Y(n428) );
  NOR2BXL U440 ( .AN(n1154), .B(n1051), .Y(n182) );
  OAI22XL U441 ( .A0(n808), .A1(n179), .B0(n185), .B1(n1153), .Y(n183) );
  OAI22XL U442 ( .A0(n1053), .A1(n189), .B0(n1051), .B1(n188), .Y(n190) );
  NAND2BXL U443 ( .AN(n1154), .B(n774), .Y(n188) );
  NOR2BXL U444 ( .AN(n1154), .B(n9), .Y(n207) );
  OAI22XL U445 ( .A0(n808), .A1(n193), .B0(n192), .B1(n1153), .Y(n206) );
  OAI22XL U446 ( .A0(n1053), .A1(n195), .B0(n1051), .B1(n194), .Y(n205) );
  OAI22XL U447 ( .A0(n1053), .A1(n194), .B0(n1051), .B1(n174), .Y(n204) );
  XNOR2XL U448 ( .A(n777), .B(n1154), .Y(n176) );
  OAI22XL U449 ( .A0(n1053), .A1(n174), .B0(n1051), .B1(n166), .Y(n173) );
  BUFX3 U450 ( .A(A[0]), .Y(n1154) );
  NOR2X1 U451 ( .A(n285), .B(n284), .Y(n871) );
  INVXL U452 ( .A(n1216), .Y(n1217) );
  NOR2X1 U453 ( .A(n1046), .B(n1215), .Y(n1221) );
  NOR2XL U454 ( .A(n1046), .B(n1209), .Y(n1232) );
  INVXL U455 ( .A(n1222), .Y(n1231) );
  OAI21XL U456 ( .A0(n906), .A1(n907), .B0(n905), .Y(n116) );
  OAI2BB1X1 U457 ( .A0N(n1001), .A1N(n1000), .B0(n82), .Y(n1004) );
  OAI21XL U458 ( .A0(n1000), .A1(n1001), .B0(n999), .Y(n82) );
  XOR3X2 U459 ( .A(n1001), .B(n1000), .C(n999), .Y(n1014) );
  INVX1 U460 ( .A(n1065), .Y(n87) );
  XNOR2X1 U461 ( .A(n1063), .B(n89), .Y(n1109) );
  OAI22XL U462 ( .A0(n808), .A1(n1154), .B0(n179), .B1(n1153), .Y(n1283) );
  NAND2XL U463 ( .A(n181), .B(n808), .Y(n1282) );
  NAND2BXL U464 ( .AN(n1154), .B(n746), .Y(n181) );
  NAND2XL U465 ( .A(n1283), .B(n1282), .Y(n1284) );
  NAND2XL U466 ( .A(n183), .B(n182), .Y(n1309) );
  INVXL U467 ( .A(n1284), .Y(n1311) );
  INVXL U468 ( .A(n1291), .Y(n201) );
  NOR2XL U469 ( .A(n209), .B(n208), .Y(n1313) );
  NAND2XL U470 ( .A(n209), .B(n208), .Y(n1314) );
  INVXL U471 ( .A(n1254), .Y(n1267) );
  NOR2X1 U472 ( .A(n304), .B(n301), .Y(n306) );
  NOR2X1 U473 ( .A(n1361), .B(n1360), .Y(n304) );
  OAI21XL U474 ( .A0(n1303), .A1(n1334), .B0(n1335), .Y(n348) );
  INVXL U475 ( .A(n1276), .Y(n1243) );
  INVXL U476 ( .A(n1270), .Y(n1244) );
  INVXL U477 ( .A(n1328), .Y(n1248) );
  INVXL U478 ( .A(n1295), .Y(n1242) );
  NAND2XL U479 ( .A(n1269), .B(n1272), .Y(n1294) );
  NAND2XL U480 ( .A(n306), .B(n305), .Y(n60) );
  AOI2BB1X1 U481 ( .A0N(n304), .A1N(n543), .B0(n145), .Y(n143) );
  AND2X2 U482 ( .A(n302), .B(n306), .Y(n147) );
  AOI21XL U483 ( .A0(n1276), .A1(n1248), .B0(n1247), .Y(n1249) );
  INVXL U484 ( .A(n1329), .Y(n1247) );
  NAND2XL U485 ( .A(n1270), .B(n1248), .Y(n1250) );
  INVXL U486 ( .A(n1326), .Y(n1251) );
  INVXL U487 ( .A(n1347), .Y(n297) );
  AOI21XL U488 ( .A0(n556), .A1(n302), .B0(n305), .Y(n541) );
  INVXL U489 ( .A(n301), .Y(n544) );
  INVXL U490 ( .A(n438), .Y(n473) );
  INVXL U491 ( .A(n436), .Y(n437) );
  INVXL U492 ( .A(n1338), .Y(n474) );
  NAND2XL U493 ( .A(n398), .B(n1335), .Y(n399) );
  INVXL U494 ( .A(n1334), .Y(n398) );
  AOI21XL U495 ( .A0(n438), .A1(n474), .B0(n439), .Y(n440) );
  INVXL U496 ( .A(n1339), .Y(n439) );
  AND2XL U497 ( .A(n436), .B(n474), .Y(n59) );
  INVXL U498 ( .A(n1336), .Y(n441) );
  NAND2XL U499 ( .A(n347), .B(n1235), .Y(n349) );
  AOI21XL U500 ( .A0(n348), .A1(n1235), .B0(n1238), .Y(n154) );
  XNOR2XL U501 ( .A(n777), .B(n1028), .Y(n248) );
  XNOR2X1 U502 ( .A(n585), .B(n1043), .Y(n247) );
  XNOR2XL U503 ( .A(n777), .B(n772), .Y(n218) );
  XNOR2XL U504 ( .A(n799), .B(n1154), .Y(n279) );
  NAND2BXL U505 ( .AN(n1154), .B(n1185), .Y(n748) );
  XNOR2XL U506 ( .A(n746), .B(n1026), .Y(n747) );
  XNOR2X1 U507 ( .A(n1185), .B(n732), .Y(n796) );
  XNOR2XL U508 ( .A(n1185), .B(n1154), .Y(n797) );
  OAI22XL U509 ( .A0(n808), .A1(n224), .B0(n253), .B1(n1153), .Y(n252) );
  CMPR32X1 U510 ( .A(n274), .B(n273), .C(n272), .CO(n880), .S(n270) );
  XNOR2XL U511 ( .A(n1044), .B(n1026), .Y(n418) );
  XNOR2XL U512 ( .A(n1185), .B(n668), .Y(n457) );
  XNOR2XL U513 ( .A(n746), .B(A[24]), .Y(n919) );
  XNOR2XL U514 ( .A(n908), .B(A[15]), .Y(n1054) );
  XNOR2XL U515 ( .A(n1210), .B(n1154), .Y(n678) );
  XNOR2XL U516 ( .A(n1185), .B(n798), .Y(n733) );
  XNOR2XL U517 ( .A(n1044), .B(n719), .Y(n321) );
  XNOR2XL U518 ( .A(n585), .B(A[25]), .Y(n356) );
  INVXL U519 ( .A(n356), .Y(n357) );
  XNOR2X1 U520 ( .A(n1036), .B(n1030), .Y(n683) );
  XNOR2XL U521 ( .A(n1185), .B(n1043), .Y(n685) );
  XNOR2XL U522 ( .A(n799), .B(n719), .Y(n458) );
  XNOR2XL U523 ( .A(n799), .B(A[19]), .Y(n421) );
  XNOR2XL U524 ( .A(n1185), .B(n915), .Y(n416) );
  XNOR2XL U525 ( .A(n585), .B(n1154), .Y(n164) );
  XNOR2XL U526 ( .A(n777), .B(n1043), .Y(n219) );
  OAI22XL U527 ( .A0(n808), .A1(n161), .B0(n225), .B1(n1153), .Y(n221) );
  OAI22XL U528 ( .A0(n1077), .A1(n355), .B0(n6), .B1(n159), .Y(n220) );
  NAND2BXL U529 ( .AN(n1154), .B(n585), .Y(n159) );
  XNOR2XL U530 ( .A(n777), .B(n798), .Y(n165) );
  AOI21XL U531 ( .A0(n1238), .A1(n1237), .B0(n1236), .Y(n1239) );
  INVXL U532 ( .A(n1331), .Y(n1236) );
  INVXL U533 ( .A(n1325), .Y(n1271) );
  OAI21XL U534 ( .A0(n868), .A1(n1318), .B0(n1319), .Y(n822) );
  OAI21XL U535 ( .A0(n868), .A1(n1350), .B0(n1355), .Y(n788) );
  NAND2XL U536 ( .A(n755), .B(n1347), .Y(n756) );
  NAND2XL U537 ( .A(n317), .B(n316), .Y(n318) );
  AOI21XL U538 ( .A0(n144), .A1(n150), .B0(n149), .Y(n148) );
  XOR2X1 U539 ( .A(n156), .B(n55), .Y(PRODUCT[23]) );
  AND2XL U540 ( .A(n652), .B(n651), .Y(n55) );
  XNOR2X1 U541 ( .A(n137), .B(n58), .Y(PRODUCT[24]) );
  AND2XL U542 ( .A(n566), .B(n1343), .Y(n58) );
  NAND2XL U543 ( .A(n553), .B(n552), .Y(n554) );
  NAND2XL U544 ( .A(n502), .B(n1341), .Y(n503) );
  CMPR32X1 U545 ( .A(n236), .B(n235), .C(n234), .CO(n259), .S(n237) );
  OAI22XL U546 ( .A0(n690), .A1(n217), .B0(n1051), .B1(n222), .Y(n236) );
  OAI22X1 U547 ( .A0(n1056), .A1(n219), .B0(n9), .B1(n218), .Y(n235) );
  ADDFX2 U548 ( .A(n230), .B(n229), .CI(n228), .CO(n250), .S(n239) );
  OAI22XL U549 ( .A0(n808), .A1(n225), .B0(n224), .B1(n1153), .Y(n229) );
  ADDFX2 U550 ( .A(n771), .B(n770), .CI(n769), .CO(n766), .S(n825) );
  OAI22X1 U551 ( .A0(n808), .A1(n747), .B0(n731), .B1(n1153), .Y(n770) );
  OAI22XL U552 ( .A0(n1187), .A1(n796), .B0(n5), .B1(n733), .Y(n769) );
  ADDFX2 U553 ( .A(n846), .B(n845), .CI(n844), .CO(n883), .S(n878) );
  OAI22XL U554 ( .A0(n1053), .A1(n280), .B0(n1051), .B1(n814), .Y(n844) );
  OAI22XL U555 ( .A0(n1049), .A1(n279), .B0(n8), .B1(n810), .Y(n845) );
  OAI22XL U556 ( .A0(n1077), .A1(n278), .B0(n6), .B1(n812), .Y(n846) );
  OAI22XL U557 ( .A0(n1049), .A1(n810), .B0(n8), .B1(n809), .Y(n836) );
  OAI22XL U558 ( .A0(n808), .A1(n807), .B0(n806), .B1(n1153), .Y(n837) );
  OAI22XL U559 ( .A0(n1056), .A1(n816), .B0(n9), .B1(n815), .Y(n850) );
  OAI22XL U560 ( .A0(n1077), .A1(n812), .B0(n6), .B1(n811), .Y(n852) );
  OAI22XL U561 ( .A0(n1053), .A1(n814), .B0(n1051), .B1(n813), .Y(n851) );
  OAI22XL U562 ( .A0(n1056), .A1(n815), .B0(n9), .B1(n778), .Y(n829) );
  OAI22X1 U563 ( .A0(n1088), .A1(n832), .B0(n1086), .B1(n773), .Y(n831) );
  XNOR2XL U564 ( .A(n1185), .B(A[25]), .Y(n1203) );
  XNOR2XL U565 ( .A(n1044), .B(n1201), .Y(n1202) );
  XNOR2XL U566 ( .A(n1185), .B(A[24]), .Y(n1186) );
  XNOR2XL U567 ( .A(n1210), .B(n1201), .Y(n1182) );
  XNOR2XL U568 ( .A(n1044), .B(n1183), .Y(n1184) );
  CMPR32X1 U569 ( .A(n781), .B(n780), .C(n779), .CO(n794), .S(n823) );
  OAI22XL U570 ( .A0(n1088), .A1(n773), .B0(n1086), .B1(n737), .Y(n781) );
  OAI22XL U571 ( .A0(n1056), .A1(n778), .B0(n9), .B1(n743), .Y(n803) );
  OAI22XL U572 ( .A0(n1077), .A1(n795), .B0(n6), .B1(n744), .Y(n802) );
  ADDFX2 U573 ( .A(n828), .B(n827), .CI(n826), .CO(n840), .S(n855) );
  OAI22XL U574 ( .A0(n1049), .A1(n809), .B0(n8), .B1(n800), .Y(n826) );
  OAI22XL U575 ( .A0(n1077), .A1(n811), .B0(n6), .B1(n795), .Y(n828) );
  OAI22XL U576 ( .A0(n1056), .A1(n263), .B0(n9), .B1(n816), .Y(n849) );
  XNOR2XL U577 ( .A(n916), .B(n596), .Y(n456) );
  XNOR2XL U578 ( .A(n585), .B(n1201), .Y(n455) );
  XNOR2XL U579 ( .A(n1044), .B(n1035), .Y(n490) );
  XNOR2XL U580 ( .A(n669), .B(n1183), .Y(n595) );
  XNOR2XL U581 ( .A(n916), .B(A[15]), .Y(n598) );
  NOR2X1 U582 ( .A(n1046), .B(n571), .Y(n580) );
  XNOR2XL U583 ( .A(n1044), .B(A[6]), .Y(n571) );
  NOR2X1 U584 ( .A(n1046), .B(n579), .Y(n601) );
  XNOR2XL U585 ( .A(n1044), .B(n1030), .Y(n579) );
  XNOR2X1 U586 ( .A(n1210), .B(n920), .Y(n587) );
  XNOR2XL U587 ( .A(n585), .B(n915), .Y(n586) );
  XNOR2XL U588 ( .A(n1185), .B(n1035), .Y(n588) );
  XNOR2XL U589 ( .A(n746), .B(A[19]), .Y(n1041) );
  ADDFX2 U590 ( .A(n608), .B(n607), .CI(n606), .CO(n617), .S(n642) );
  OAI22XL U591 ( .A0(n1053), .A1(n604), .B0(n1051), .B1(n575), .Y(n607) );
  OAI22XL U592 ( .A0(n1049), .A1(n603), .B0(n8), .B1(n574), .Y(n608) );
  ADDFX2 U593 ( .A(n634), .B(n633), .CI(n632), .CO(n643), .S(n1067) );
  OAI22XL U594 ( .A0(n1053), .A1(n630), .B0(n1051), .B1(n604), .Y(n633) );
  OAI22XL U595 ( .A0(n1049), .A1(n629), .B0(n8), .B1(n603), .Y(n634) );
  XNOR2X1 U596 ( .A(n777), .B(A[14]), .Y(n1055) );
  NAND2BXL U597 ( .AN(n1154), .B(n1210), .Y(n670) );
  NOR2BXL U598 ( .AN(n1154), .B(n1046), .Y(n681) );
  OAI22X1 U599 ( .A0(n1218), .A1(n677), .B0(n1219), .B1(n676), .Y(n679) );
  OAI22XL U600 ( .A0(n1056), .A1(n694), .B0(n9), .B1(n715), .Y(n711) );
  OAI22XL U601 ( .A0(n1053), .A1(n688), .B0(n1051), .B1(n687), .Y(n712) );
  XNOR2X1 U602 ( .A(n1210), .B(n798), .Y(n676) );
  XNOR2XL U603 ( .A(n1044), .B(n732), .Y(n665) );
  OAI22XL U604 ( .A0(n808), .A1(n674), .B0(n720), .B1(n1153), .Y(n723) );
  NOR2XL U605 ( .A(n1046), .B(n666), .Y(n722) );
  NAND2BXL U606 ( .AN(n1154), .B(n1044), .Y(n666) );
  XNOR2XL U607 ( .A(n1185), .B(n719), .Y(n415) );
  XNOR2XL U608 ( .A(n916), .B(n1208), .Y(n377) );
  XNOR2X1 U609 ( .A(n1185), .B(A[19]), .Y(n376) );
  INVXL U610 ( .A(n380), .Y(n76) );
  INVXL U611 ( .A(n8), .Y(n75) );
  XNOR2XL U612 ( .A(n1210), .B(n915), .Y(n379) );
  XNOR2XL U613 ( .A(n1044), .B(A[15]), .Y(n378) );
  XNOR2XL U614 ( .A(n799), .B(n1183), .Y(n380) );
  XNOR2XL U615 ( .A(n799), .B(n596), .Y(n414) );
  ADDFX2 U616 ( .A(n366), .B(n365), .CI(n364), .CO(n360), .S(n391) );
  OAI22XL U617 ( .A0(n1049), .A1(n375), .B0(n8), .B1(n329), .Y(n365) );
  INVXL U618 ( .A(n331), .Y(n364) );
  CMPR32X1 U619 ( .A(n765), .B(n764), .C(n763), .CO(n762), .S(n819) );
  OAI22XL U620 ( .A0(n1077), .A1(n744), .B0(n6), .B1(n698), .Y(n763) );
  OAI22XL U621 ( .A0(n690), .A1(n739), .B0(n1051), .B1(n689), .Y(n765) );
  OAI22XL U622 ( .A0(n1049), .A1(n738), .B0(n8), .B1(n696), .Y(n764) );
  OAI22XL U623 ( .A0(n1077), .A1(n698), .B0(n6), .B1(n697), .Y(n702) );
  OAI22XL U624 ( .A0(n1056), .A1(n727), .B0(n9), .B1(n694), .Y(n704) );
  OAI22XL U625 ( .A0(n1088), .A1(n449), .B0(n1086), .B1(n413), .Y(n425) );
  OAI22XL U626 ( .A0(n1077), .A1(n419), .B0(n6), .B1(n411), .Y(n427) );
  OAI2BB1XL U627 ( .A0N(n9), .A1N(n1056), .B0(n404), .Y(n422) );
  INVXL U628 ( .A(n403), .Y(n404) );
  XNOR2XL U629 ( .A(n746), .B(n798), .Y(n185) );
  XNOR2XL U630 ( .A(n746), .B(n1043), .Y(n193) );
  XNOR2XL U631 ( .A(n777), .B(n732), .Y(n175) );
  OAI22XL U632 ( .A0(n808), .A1(n192), .B0(n167), .B1(n1153), .Y(n178) );
  NAND2BXL U633 ( .AN(n1154), .B(n777), .Y(n169) );
  OAI22X1 U634 ( .A0(n808), .A1(n167), .B0(n161), .B1(n1153), .Y(n170) );
  INVXL U635 ( .A(n170), .Y(n107) );
  NAND2XL U636 ( .A(n1272), .B(n1325), .Y(n1262) );
  NOR2XL U637 ( .A(n1046), .B(n336), .Y(n1181) );
  OAI2BB1XL U638 ( .A0N(n8), .A1N(n71), .B0(n338), .Y(n1179) );
  XNOR2XL U639 ( .A(n1044), .B(n596), .Y(n336) );
  ADDFX2 U640 ( .A(n794), .B(n793), .CI(n792), .CO(n782), .S(n858) );
  OAI22XL U641 ( .A0(n1088), .A1(n933), .B0(n1086), .B1(n917), .Y(n953) );
  OAI22XL U642 ( .A0(n1056), .A1(n928), .B0(n9), .B1(n909), .Y(n950) );
  OAI22XL U643 ( .A0(n1056), .A1(n909), .B0(n9), .B1(n505), .Y(n520) );
  INVXL U644 ( .A(n507), .Y(n519) );
  OAI22XL U645 ( .A0(n1187), .A1(n911), .B0(n5), .B1(n504), .Y(n521) );
  OAI22XL U646 ( .A0(n1088), .A1(n917), .B0(n1086), .B1(n509), .Y(n524) );
  OAI22XL U647 ( .A0(n1049), .A1(n516), .B0(n8), .B1(n510), .Y(n523) );
  OAI2BB1XL U648 ( .A0N(n1153), .A1N(n808), .B0(n518), .Y(n930) );
  OAI22XL U649 ( .A0(n1049), .A1(n924), .B0(n8), .B1(n516), .Y(n932) );
  OAI22XL U650 ( .A0(n1053), .A1(n926), .B0(n1051), .B1(n517), .Y(n931) );
  CMPR32X1 U651 ( .A(n977), .B(n976), .C(n975), .CO(n978), .S(n1002) );
  OAI22XL U652 ( .A0(n1056), .A1(n929), .B0(n9), .B1(n928), .Y(n966) );
  OAI22XL U653 ( .A0(n1053), .A1(n927), .B0(n1051), .B1(n926), .Y(n967) );
  NOR2BXL U654 ( .AN(n626), .B(n84), .Y(n609) );
  OAI22X1 U655 ( .A0(n1077), .A1(n618), .B0(n6), .B1(n568), .Y(n623) );
  OAI22XL U656 ( .A0(n1187), .A1(n620), .B0(n5), .B1(n570), .Y(n621) );
  OAI22X2 U657 ( .A0(n1218), .A1(n619), .B0(n1219), .B1(n569), .Y(n622) );
  OAI22XL U658 ( .A0(n625), .A1(n1037), .B0(n1086), .B1(n624), .Y(n637) );
  XNOR2X1 U659 ( .A(n1210), .B(n1030), .Y(n619) );
  XNOR2X1 U660 ( .A(n585), .B(A[15]), .Y(n618) );
  XNOR2XL U661 ( .A(n1185), .B(n920), .Y(n620) );
  XNOR2X1 U662 ( .A(n1210), .B(A[6]), .Y(n1029) );
  XNOR2X1 U663 ( .A(n585), .B(A[14]), .Y(n1027) );
  XNOR2XL U664 ( .A(n1185), .B(n776), .Y(n1031) );
  INVX1 U665 ( .A(n65), .Y(n66) );
  OAI22X1 U666 ( .A0(n1077), .A1(n1076), .B0(n6), .B1(n1075), .Y(n1119) );
  OAI22XL U667 ( .A0(n1187), .A1(n1081), .B0(n5), .B1(n1080), .Y(n1117) );
  ADDFX2 U668 ( .A(n1095), .B(n1094), .CI(n1093), .CO(n1131), .S(n1138) );
  OAI22XL U669 ( .A0(n1053), .A1(n687), .B0(n1051), .B1(n1052), .Y(n1093) );
  NOR2XL U670 ( .A(n1046), .B(n319), .Y(n342) );
  INVXL U671 ( .A(n1180), .Y(n341) );
  OAI22XL U672 ( .A0(n1218), .A1(n325), .B0(n1219), .B1(n340), .Y(n343) );
  OAI22XL U673 ( .A0(n1187), .A1(n326), .B0(n5), .B1(n339), .Y(n346) );
  NOR2XL U674 ( .A(n1046), .B(n353), .Y(n368) );
  OAI22XL U675 ( .A0(n1187), .A1(n363), .B0(n5), .B1(n352), .Y(n369) );
  XNOR2XL U676 ( .A(n1044), .B(n915), .Y(n353) );
  CMPR32X1 U677 ( .A(n392), .B(n391), .C(n390), .CO(n393), .S(n431) );
  ADDFX2 U678 ( .A(n784), .B(n783), .CI(n782), .CO(n758), .S(n789) );
  NAND2XL U679 ( .A(n487), .B(n488), .Y(n139) );
  OAI21XL U680 ( .A0(n487), .A1(n488), .B0(n486), .Y(n140) );
  ADDFX2 U681 ( .A(n64), .B(n241), .CI(n240), .CO(n243), .S(n213) );
  NAND2XL U682 ( .A(n109), .B(n170), .Y(n105) );
  INVXL U683 ( .A(n1304), .Y(n1305) );
  OR2XL U684 ( .A(n1296), .B(n1302), .Y(n1306) );
  NAND2XL U685 ( .A(n1279), .B(n1323), .Y(n1280) );
  NAND2BX1 U686 ( .AN(n244), .B(n94), .Y(n902) );
  OAI22XL U687 ( .A0(n1218), .A1(n1197), .B0(n1219), .B1(n1211), .Y(n1229) );
  OAI21XL U688 ( .A0(n104), .A1(n103), .B0(n102), .Y(n753) );
  OAI21XL U689 ( .A0(n758), .A1(n759), .B0(n757), .Y(n102) );
  XNOR3X2 U690 ( .A(n134), .B(n789), .C(n790), .Y(n821) );
  ADDFX2 U691 ( .A(n858), .B(n857), .CI(n856), .CO(n820), .S(n865) );
  INVXL U692 ( .A(mult_x_1_n306), .Y(n869) );
  OR2X2 U693 ( .A(n865), .B(n864), .Y(n1156) );
  NOR2XL U694 ( .A(n871), .B(n890), .Y(n873) );
  XOR2XL U695 ( .A(n487), .B(n488), .Y(n100) );
  ADDFX2 U696 ( .A(n956), .B(n955), .CI(n954), .CO(n905), .S(n957) );
  ADDFX2 U697 ( .A(n962), .B(n961), .CI(n960), .CO(n956), .S(n983) );
  INVX1 U698 ( .A(n983), .Y(n123) );
  ADDFX2 U699 ( .A(n752), .B(n751), .CI(n750), .CO(n1151), .S(n757) );
  NAND2XL U700 ( .A(n388), .B(n389), .Y(n110) );
  OR2X2 U701 ( .A(n790), .B(n791), .Y(n133) );
  XOR3X2 U702 ( .A(n759), .B(n758), .C(n757), .Y(n786) );
  NOR2XL U703 ( .A(n1175), .B(n1174), .Y(mult_x_1_n136) );
  NOR2XL U704 ( .A(n1234), .B(n1233), .Y(mult_x_1_n109) );
  NOR2BXL U705 ( .AN(n1154), .B(n1153), .Y(n1401) );
  NAND2XL U706 ( .A(n902), .B(n901), .Y(n903) );
  NAND2XL U707 ( .A(n1226), .B(n1225), .Y(mult_x_1_n58) );
  NAND2XL U708 ( .A(n1224), .B(n1223), .Y(n1225) );
  NAND2XL U709 ( .A(n1234), .B(n1233), .Y(mult_x_1_n110) );
  NOR2XL U710 ( .A(n1207), .B(n1206), .Y(mult_x_1_n120) );
  NAND2XL U711 ( .A(n1207), .B(n1206), .Y(mult_x_1_n121) );
  NOR2XL U712 ( .A(n1192), .B(n1191), .Y(mult_x_1_n129) );
  NAND2XL U713 ( .A(n1192), .B(n1191), .Y(mult_x_1_n130) );
  NAND2XL U714 ( .A(n57), .B(n1173), .Y(mult_x_1_n85) );
  OAI21XL U715 ( .A0(n123), .A1(n122), .B0(n121), .Y(mult_x_1_n521) );
  OAI21XL U716 ( .A0(n982), .A1(n983), .B0(n981), .Y(n121) );
  XNOR3X2 U717 ( .A(n123), .B(n982), .C(n981), .Y(mult_x_1_n522) );
  NAND2X1 U718 ( .A(n114), .B(n113), .Y(n1006) );
  NAND2XL U719 ( .A(n1016), .B(n1015), .Y(n113) );
  NAND2X1 U720 ( .A(n115), .B(n1014), .Y(n114) );
  XOR3X2 U721 ( .A(n1015), .B(n1014), .C(n1016), .Y(n1017) );
  NAND2X1 U722 ( .A(n1064), .B(n1065), .Y(n85) );
  OAI21XL U723 ( .A0(n1136), .A1(n1137), .B0(n1135), .Y(n125) );
  INVX1 U724 ( .A(n1137), .Y(n126) );
  NAND2XL U725 ( .A(n1310), .B(n1309), .Y(n1312) );
  NAND2XL U726 ( .A(n1288), .B(n1287), .Y(n1290) );
  INVXL U727 ( .A(n1286), .Y(n1288) );
  NAND2XL U728 ( .A(n198), .B(n1291), .Y(n1293) );
  NAND2XL U729 ( .A(n1315), .B(n1314), .Y(n1317) );
  INVXL U730 ( .A(n1313), .Y(n1315) );
  NAND2XL U731 ( .A(n1266), .B(n1265), .Y(n1268) );
  INVXL U732 ( .A(n1264), .Y(n1266) );
  NAND2XL U733 ( .A(n1257), .B(n1256), .Y(n1258) );
  CLKINVX3 U734 ( .A(B[9]), .Y(n322) );
  INVX4 U735 ( .A(n322), .Y(n1036) );
  AND2X2 U736 ( .A(n60), .B(n143), .Y(n54) );
  OR2X2 U737 ( .A(n1167), .B(n1166), .Y(n57) );
  OAI21XL U738 ( .A0(n551), .A1(n558), .B0(n552), .Y(n305) );
  NOR2X1 U739 ( .A(n1373), .B(n1372), .Y(n1157) );
  NOR2X1 U740 ( .A(n1157), .B(n315), .Y(n561) );
  NAND2X1 U741 ( .A(n561), .B(n289), .Y(n557) );
  INVX1 U742 ( .A(n557), .Y(n157) );
  XNOR2X1 U743 ( .A(n1136), .B(n126), .Y(n61) );
  XOR3X2 U744 ( .A(n907), .B(n906), .C(n905), .Y(n62) );
  INVXL U745 ( .A(n242), .Y(n63) );
  XNOR2X1 U746 ( .A(n1044), .B(n798), .Y(n721) );
  CMPR22X1 U747 ( .A(n1092), .B(n1091), .CO(n1099), .S(n1121) );
  OAI22X1 U748 ( .A0(n808), .A1(n720), .B0(n1042), .B1(n1040), .Y(n1092) );
  NOR2X1 U749 ( .A(n6), .B(n10), .Y(n109) );
  AOI21X1 U750 ( .A0(n904), .A1(n902), .B0(n896), .Y(n900) );
  XNOR2X2 U751 ( .A(B[6]), .B(B[5]), .Y(n160) );
  CMPR22X1 U752 ( .A(n1039), .B(n1038), .CO(n635), .S(n1061) );
  OAI22X1 U753 ( .A0(n808), .A1(n1041), .B0(n627), .B1(n1153), .Y(n1039) );
  NOR2X1 U754 ( .A(n1046), .B(n628), .Y(n1038) );
  INVXL U755 ( .A(n1100), .Y(n65) );
  CMPR22X1 U756 ( .A(n805), .B(n804), .CO(n801), .S(n843) );
  NOR2X1 U757 ( .A(n1359), .B(n1358), .Y(n536) );
  INVXL U758 ( .A(n610), .Y(n67) );
  INVX1 U759 ( .A(n67), .Y(n68) );
  INVXL U760 ( .A(n767), .Y(n69) );
  INVX1 U761 ( .A(n69), .Y(n70) );
  CMPR22X1 U762 ( .A(n835), .B(n834), .CO(n876), .S(n847) );
  OAI22X1 U763 ( .A0(n1049), .A1(n268), .B0(n8), .B1(n267), .Y(n834) );
  CMPR22X1 U764 ( .A(n936), .B(n935), .CO(n952), .S(n970) );
  OAI22X1 U765 ( .A0(n808), .A1(n578), .B0(n599), .B1(n1153), .Y(n602) );
  OAI22X1 U766 ( .A0(n1088), .A1(n361), .B0(n1086), .B1(n323), .Y(n331) );
  NOR2X1 U767 ( .A(n155), .B(n308), .Y(n1303) );
  CMPR22X1 U768 ( .A(n197), .B(n196), .CO(n199), .S(n191) );
  OAI22X1 U769 ( .A0(n690), .A1(n186), .B0(n1051), .B1(n195), .Y(n196) );
  XOR2X1 U770 ( .A(n1307), .B(n538), .Y(PRODUCT[29]) );
  XOR2X1 U771 ( .A(n148), .B(n318), .Y(PRODUCT[22]) );
  XNOR2X1 U772 ( .A(n555), .B(n554), .Y(PRODUCT[26]) );
  OAI21X1 U773 ( .A0(n626), .A1(n84), .B0(n83), .Y(n636) );
  OAI21XL U774 ( .A0(n573), .A1(n1046), .B0(n626), .Y(n83) );
  INVXL U775 ( .A(n77), .Y(n71) );
  XOR2X1 U776 ( .A(n170), .B(n109), .Y(n108) );
  NAND2X1 U777 ( .A(n72), .B(n73), .Y(n389) );
  XOR2X1 U778 ( .A(n388), .B(n389), .Y(n112) );
  OAI2BB1X1 U779 ( .A0N(n59), .A1N(n78), .B0(n440), .Y(n146) );
  OR2X2 U780 ( .A(n573), .B(n1046), .Y(n84) );
  XNOR2X2 U781 ( .A(n1064), .B(n1065), .Y(n89) );
  AOI21X1 U782 ( .A0(n896), .A1(n898), .B0(n91), .Y(n92) );
  INVX1 U783 ( .A(n874), .Y(n894) );
  OAI21X2 U784 ( .A0(n895), .A1(n93), .B0(n92), .Y(n874) );
  OAI21XL U785 ( .A0(n1255), .A1(n1265), .B0(n1256), .Y(n95) );
  AND2X2 U786 ( .A(n214), .B(n1254), .Y(n96) );
  AOI21X4 U787 ( .A0(n99), .A1(n1036), .B0(n98), .Y(n97) );
  NOR2X2 U788 ( .A(n223), .B(n1086), .Y(n98) );
  OR2X2 U789 ( .A(n1016), .B(n1015), .Y(n115) );
  OAI21X1 U790 ( .A0(n655), .A1(n661), .B0(n656), .Y(n128) );
  NAND2X1 U791 ( .A(n1374), .B(n1375), .Y(n656) );
  NOR2X2 U792 ( .A(n1374), .B(n1375), .Y(n655) );
  AOI2BB1X2 U793 ( .A0N(n296), .A1N(n1346), .B0(n297), .Y(n300) );
  XOR2X1 U794 ( .A(n756), .B(n296), .Y(PRODUCT[17]) );
  NAND2X4 U795 ( .A(n266), .B(n120), .Y(n1049) );
  XNOR2X2 U796 ( .A(B[10]), .B(B[9]), .Y(n266) );
  OAI21X4 U797 ( .A0(n129), .A1(n296), .B0(n127), .Y(n144) );
  OAI21X1 U798 ( .A0(n1347), .A1(n1344), .B0(n1345), .Y(n653) );
  NAND2X1 U799 ( .A(n130), .B(n654), .Y(n129) );
  NOR2X2 U800 ( .A(n655), .B(n660), .Y(n130) );
  XNOR2X1 U801 ( .A(n136), .B(n295), .Y(PRODUCT[28]) );
  OAI21XL U802 ( .A0(n1159), .A1(n293), .B0(n292), .Y(n136) );
  INVX1 U803 ( .A(n144), .Y(n1159) );
  AND2X2 U804 ( .A(n565), .B(n138), .Y(n137) );
  OAI21XL U805 ( .A0(n1307), .A1(n437), .B0(n473), .Y(n476) );
  INVX8 U806 ( .A(n355), .Y(n585) );
  NOR2X2 U807 ( .A(n1376), .B(n1377), .Y(n660) );
  AOI21XL U808 ( .A0(n556), .A1(n291), .B0(n290), .Y(n292) );
  ADDFX2 U809 ( .A(n527), .B(n526), .CI(n525), .CO(n514), .S(n955) );
  XNOR2X1 U810 ( .A(B[16]), .B(B[15]), .Y(n417) );
  INVX8 U811 ( .A(n672), .Y(n1210) );
  AOI21XL U812 ( .A0(n1273), .A1(n1272), .B0(n1271), .Y(n1297) );
  XNOR2XL U813 ( .A(n669), .B(n719), .Y(n630) );
  XNOR2X1 U814 ( .A(n1210), .B(n668), .Y(n412) );
  OAI22X1 U815 ( .A0(n1077), .A1(n164), .B0(n6), .B1(n227), .Y(n232) );
  XNOR2XL U816 ( .A(n1185), .B(n745), .Y(n947) );
  XNOR2XL U817 ( .A(n1185), .B(n1030), .Y(n1080) );
  XNOR2XL U818 ( .A(n1185), .B(n772), .Y(n684) );
  ADDFX2 U819 ( .A(n693), .B(n692), .CI(n691), .CO(n700), .S(n761) );
  BUFX4 U820 ( .A(B[1]), .Y(n746) );
  XNOR2X1 U821 ( .A(n746), .B(n1030), .Y(n225) );
  BUFX3 U822 ( .A(n1040), .Y(n1153) );
  XOR2X1 U823 ( .A(B[6]), .B(B[7]), .Y(n158) );
  XNOR2X1 U824 ( .A(n746), .B(n1028), .Y(n167) );
  XOR2X1 U825 ( .A(B[4]), .B(B[5]), .Y(n162) );
  XNOR2X1 U826 ( .A(B[4]), .B(B[3]), .Y(n168) );
  NAND2X2 U827 ( .A(n162), .B(n168), .Y(n728) );
  CLKINVX3 U828 ( .A(B[5]), .Y(n402) );
  XOR2X1 U829 ( .A(B[2]), .B(B[3]), .Y(n163) );
  XNOR2X1 U830 ( .A(B[2]), .B(B[1]), .Y(n187) );
  CLKINVX3 U831 ( .A(n189), .Y(n774) );
  XNOR2X1 U832 ( .A(n774), .B(n772), .Y(n166) );
  XNOR2X1 U833 ( .A(n774), .B(n1028), .Y(n217) );
  OAI22X1 U834 ( .A0(n1053), .A1(n166), .B0(n1051), .B1(n217), .Y(n233) );
  XNOR2X1 U835 ( .A(n746), .B(n772), .Y(n192) );
  OAI22XL U836 ( .A0(n1056), .A1(n402), .B0(n9), .B1(n169), .Y(n177) );
  XNOR2X1 U837 ( .A(n774), .B(n798), .Y(n194) );
  OAI22XL U838 ( .A0(n728), .A1(n176), .B0(n9), .B1(n175), .Y(n203) );
  ADDHXL U839 ( .A(n178), .B(n177), .CO(n172), .S(n202) );
  OAI22X1 U840 ( .A0(n808), .A1(n185), .B0(n193), .B1(n1153), .Y(n197) );
  XNOR2XL U841 ( .A(n774), .B(n732), .Y(n195) );
  BUFX3 U842 ( .A(n187), .Y(n1051) );
  NOR2XL U843 ( .A(n191), .B(n190), .Y(n1286) );
  OAI21XL U844 ( .A0(n1289), .A1(n1286), .B0(n1287), .Y(n1292) );
  AOI21XL U845 ( .A0(n1292), .A1(n198), .B0(n201), .Y(n1316) );
  CMPR32X1 U846 ( .A(n204), .B(n203), .C(n202), .CO(n210), .S(n209) );
  CMPR32X1 U847 ( .A(n207), .B(n206), .C(n205), .CO(n208), .S(n200) );
  OAI21XL U848 ( .A0(n1316), .A1(n1313), .B0(n1314), .Y(n1254) );
  OAI22X1 U849 ( .A0(n1077), .A1(n226), .B0(n6), .B1(n247), .Y(n257) );
  XNOR2X1 U850 ( .A(n1036), .B(n1154), .Y(n216) );
  XNOR2X1 U851 ( .A(n1036), .B(n732), .Y(n254) );
  OAI22XL U852 ( .A0(n728), .A1(n218), .B0(n9), .B1(n248), .Y(n255) );
  XNOR2X1 U853 ( .A(n774), .B(A[6]), .Y(n222) );
  ADDHXL U854 ( .A(n221), .B(n220), .CO(n234), .S(n242) );
  XNOR2X1 U855 ( .A(n774), .B(n1030), .Y(n249) );
  XNOR2X1 U856 ( .A(n746), .B(n776), .Y(n224) );
  XNOR2X1 U857 ( .A(n746), .B(n920), .Y(n253) );
  NAND2BX1 U858 ( .AN(n1154), .B(n1036), .Y(n223) );
  OAI22XL U859 ( .A0(n718), .A1(n227), .B0(n6), .B1(n226), .Y(n228) );
  CMPR32X1 U860 ( .A(n239), .B(n238), .C(n237), .CO(n245), .S(n244) );
  NAND2XL U861 ( .A(n246), .B(n245), .Y(n897) );
  OAI22X1 U862 ( .A0(n1077), .A1(n247), .B0(n6), .B1(n278), .Y(n277) );
  XNOR2X1 U863 ( .A(n777), .B(A[6]), .Y(n263) );
  OAI22X1 U864 ( .A0(n1056), .A1(n248), .B0(n9), .B1(n263), .Y(n276) );
  XNOR2X1 U865 ( .A(n774), .B(n776), .Y(n280) );
  XNOR2XL U866 ( .A(n746), .B(A[10]), .Y(n265) );
  OAI22XL U867 ( .A0(n808), .A1(n253), .B0(n265), .B1(n1153), .Y(n273) );
  XNOR2X1 U868 ( .A(n1036), .B(n798), .Y(n264) );
  OAI22XL U869 ( .A0(n625), .A1(n254), .B0(n1086), .B1(n264), .Y(n272) );
  CMPR32X1 U870 ( .A(n257), .B(n256), .C(n255), .CO(n269), .S(n260) );
  ADDFHX1 U871 ( .A(n260), .B(n259), .CI(n258), .CO(n261), .S(n246) );
  NOR2X1 U872 ( .A(n262), .B(n261), .Y(n890) );
  OAI21X1 U873 ( .A0(n894), .A1(n890), .B0(n891), .Y(n288) );
  OAI22XL U874 ( .A0(n625), .A1(n264), .B0(n1086), .B1(n833), .Y(n848) );
  OAI22X1 U875 ( .A0(n808), .A1(n265), .B0(n807), .B1(n1153), .Y(n835) );
  INVX8 U876 ( .A(n268), .Y(n799) );
  XNOR2X1 U877 ( .A(n585), .B(n1028), .Y(n812) );
  XNOR2X1 U878 ( .A(n799), .B(n732), .Y(n810) );
  XNOR2X1 U879 ( .A(n774), .B(n920), .Y(n814) );
  CMPR32X1 U880 ( .A(n283), .B(n282), .C(n281), .CO(n284), .S(n262) );
  INVXL U881 ( .A(n871), .Y(n286) );
  NAND2XL U882 ( .A(n286), .B(n870), .Y(n287) );
  XNOR2X1 U883 ( .A(n288), .B(n287), .Y(n1390) );
  INVXL U884 ( .A(n302), .Y(n539) );
  NOR2X1 U885 ( .A(n1362), .B(n1363), .Y(n301) );
  NOR2XL U886 ( .A(n539), .B(n301), .Y(n291) );
  NAND2XL U887 ( .A(n291), .B(n157), .Y(n293) );
  INVXL U888 ( .A(n305), .Y(n540) );
  NAND2X1 U889 ( .A(n1362), .B(n1363), .Y(n543) );
  OAI21XL U890 ( .A0(n540), .A1(n301), .B0(n543), .Y(n290) );
  INVXL U891 ( .A(n304), .Y(n294) );
  NAND2X1 U892 ( .A(n1360), .B(n1361), .Y(n303) );
  NAND2X1 U893 ( .A(n294), .B(n303), .Y(n295) );
  INVXL U894 ( .A(n1344), .Y(n298) );
  NAND2XL U895 ( .A(n298), .B(n1345), .Y(n299) );
  XOR2X1 U896 ( .A(n300), .B(n299), .Y(PRODUCT[18]) );
  NOR2XL U897 ( .A(n536), .B(n1340), .Y(n436) );
  NOR2XL U898 ( .A(n1338), .B(n1336), .Y(n309) );
  NAND2XL U899 ( .A(n436), .B(n309), .Y(n1296) );
  NOR2XL U900 ( .A(n1296), .B(n1334), .Y(n347) );
  INVXL U901 ( .A(n347), .Y(n311) );
  NAND2X1 U902 ( .A(n1359), .B(n1358), .Y(n537) );
  OAI21XL U903 ( .A0(n1340), .A1(n537), .B0(n1341), .Y(n438) );
  OAI21XL U904 ( .A0(n1336), .A1(n1339), .B0(n1337), .Y(n308) );
  INVXL U905 ( .A(n348), .Y(n310) );
  OAI21XL U906 ( .A0(n1307), .A1(n311), .B0(n310), .Y(n313) );
  INVXL U907 ( .A(n315), .Y(n317) );
  BUFX12 U908 ( .A(n673), .Y(n1218) );
  CLKINVX3 U909 ( .A(B[15]), .Y(n672) );
  XNOR2X1 U910 ( .A(n1210), .B(n596), .Y(n325) );
  XNOR2X1 U911 ( .A(n1210), .B(n1183), .Y(n340) );
  XNOR2X1 U912 ( .A(n799), .B(A[24]), .Y(n327) );
  XNOR2X1 U913 ( .A(n799), .B(A[25]), .Y(n337) );
  OAI22X1 U914 ( .A0(n1049), .A1(n327), .B0(n8), .B1(n337), .Y(n1180) );
  CLKBUFX8 U915 ( .A(n1205), .Y(n1187) );
  BUFX8 U916 ( .A(B[13]), .Y(n1185) );
  XNOR2X1 U917 ( .A(n1185), .B(n1201), .Y(n326) );
  XNOR2X1 U918 ( .A(n1185), .B(n1208), .Y(n339) );
  CLKINVX3 U919 ( .A(n322), .Y(n916) );
  XNOR2XL U920 ( .A(n916), .B(A[24]), .Y(n361) );
  XNOR2X1 U921 ( .A(n1036), .B(A[25]), .Y(n323) );
  XNOR2X1 U922 ( .A(n1210), .B(A[19]), .Y(n328) );
  XNOR2X1 U923 ( .A(n1185), .B(n1183), .Y(n352) );
  XNOR2X1 U924 ( .A(n799), .B(n1208), .Y(n329) );
  XNOR2X1 U925 ( .A(n1210), .B(n719), .Y(n362) );
  OAI22XL U926 ( .A0(n673), .A1(n362), .B0(n1219), .B1(n328), .Y(n366) );
  XNOR2X1 U927 ( .A(n799), .B(n1201), .Y(n375) );
  CMPR32X1 U928 ( .A(n332), .B(n331), .C(n330), .CO(n345), .S(n359) );
  CMPR32X1 U929 ( .A(n335), .B(n334), .C(n333), .CO(n344), .S(n358) );
  CMPR32X1 U930 ( .A(n343), .B(n342), .C(n341), .CO(n1188), .S(n372) );
  CMPR32X1 U931 ( .A(n346), .B(n345), .C(n344), .CO(n1176), .S(n371) );
  NAND2XL U932 ( .A(n1175), .B(n1174), .Y(mult_x_1_n137) );
  XNOR2X1 U933 ( .A(n351), .B(n350), .Y(PRODUCT[35]) );
  XNOR2X1 U934 ( .A(n1185), .B(n596), .Y(n363) );
  XNOR2X1 U935 ( .A(n585), .B(A[24]), .Y(n411) );
  CMPR32X1 U936 ( .A(n360), .B(n359), .C(n358), .CO(n370), .S(n394) );
  OAI22XL U937 ( .A0(n673), .A1(n379), .B0(n1219), .B1(n362), .Y(n382) );
  CMPR32X1 U938 ( .A(n369), .B(n368), .C(n367), .CO(n395), .S(n390) );
  CMPR32X1 U939 ( .A(n372), .B(n371), .C(n370), .CO(n1175), .S(n373) );
  NOR2XL U940 ( .A(n374), .B(n373), .Y(mult_x_1_n151) );
  NAND2XL U941 ( .A(n374), .B(n373), .Y(mult_x_1_n152) );
  OAI22X1 U942 ( .A0(n1205), .A1(n415), .B0(n5), .B1(n376), .Y(n410) );
  OAI22X2 U943 ( .A0(n1088), .A1(n413), .B0(n1086), .B1(n377), .Y(n409) );
  CMPR32X1 U944 ( .A(n383), .B(n382), .C(n381), .CO(n392), .S(n430) );
  CMPR32X1 U945 ( .A(n395), .B(n394), .C(n393), .CO(n374), .S(n396) );
  NOR2XL U946 ( .A(n397), .B(n396), .Y(mult_x_1_n160) );
  NAND2XL U947 ( .A(n397), .B(n396), .Y(mult_x_1_n161) );
  XNOR2X1 U948 ( .A(n400), .B(n399), .Y(PRODUCT[33]) );
  XNOR2XL U949 ( .A(n1044), .B(A[14]), .Y(n401) );
  NOR2XL U950 ( .A(n1046), .B(n401), .Y(n424) );
  CLKINVX3 U951 ( .A(n402), .Y(n908) );
  XNOR2X1 U952 ( .A(n908), .B(A[24]), .Y(n453) );
  OAI22X2 U953 ( .A0(n1056), .A1(n453), .B0(n9), .B1(n403), .Y(n423) );
  CMPR32X1 U954 ( .A(n407), .B(n406), .C(n405), .CO(n387), .S(n444) );
  XNOR2X1 U955 ( .A(n585), .B(n1208), .Y(n419) );
  XNOR2X1 U956 ( .A(n1210), .B(A[15]), .Y(n420) );
  OAI22XL U957 ( .A0(n1218), .A1(n420), .B0(n1219), .B1(n412), .Y(n426) );
  OAI22XL U958 ( .A0(n1205), .A1(n416), .B0(n5), .B1(n415), .Y(n447) );
  NOR2XL U959 ( .A(n1046), .B(n418), .Y(n460) );
  INVXL U960 ( .A(n423), .Y(n459) );
  OAI22X1 U961 ( .A0(n1077), .A1(n455), .B0(n6), .B1(n419), .Y(n464) );
  OAI22X1 U962 ( .A0(n1218), .A1(n454), .B0(n1219), .B1(n420), .Y(n463) );
  OAI22X1 U963 ( .A0(n1049), .A1(n458), .B0(n8), .B1(n421), .Y(n462) );
  CMPR32X1 U964 ( .A(n427), .B(n426), .C(n425), .CO(n467), .S(n480) );
  CMPR32X1 U965 ( .A(n430), .B(n429), .C(n428), .CO(n432), .S(n468) );
  CMPR32X1 U966 ( .A(n433), .B(n432), .C(n431), .CO(n397), .S(n434) );
  NOR2XL U967 ( .A(n435), .B(n434), .Y(mult_x_1_n169) );
  NAND2XL U968 ( .A(n435), .B(n434), .Y(mult_x_1_n170) );
  CMPR32X1 U969 ( .A(n445), .B(n444), .C(n443), .CO(n470), .S(n479) );
  CMPR32X1 U970 ( .A(n448), .B(n447), .C(n446), .CO(n466), .S(n485) );
  XNOR2XL U971 ( .A(n1044), .B(n745), .Y(n450) );
  NOR2XL U972 ( .A(n1046), .B(n450), .Y(n508) );
  CLKINVX3 U973 ( .A(n189), .Y(n669) );
  XNOR2X1 U974 ( .A(n669), .B(A[24]), .Y(n517) );
  XNOR2X1 U975 ( .A(n774), .B(A[25]), .Y(n451) );
  OAI22X2 U976 ( .A0(n1053), .A1(n517), .B0(n1051), .B1(n451), .Y(n507) );
  XNOR2X1 U977 ( .A(n908), .B(n1208), .Y(n505) );
  OAI22X1 U978 ( .A0(n1056), .A1(n505), .B0(n9), .B1(n453), .Y(n494) );
  XNOR2X1 U979 ( .A(n1185), .B(A[15]), .Y(n504) );
  XNOR2X1 U980 ( .A(n799), .B(n915), .Y(n510) );
  ADDFHX1 U981 ( .A(n467), .B(n466), .CI(n465), .CO(n469), .S(n477) );
  CMPR32X1 U982 ( .A(n470), .B(n469), .C(n468), .CO(n435), .S(n471) );
  NOR2XL U983 ( .A(n472), .B(n471), .Y(mult_x_1_n176) );
  NAND2XL U984 ( .A(n472), .B(n471), .Y(mult_x_1_n177) );
  ADDFHX1 U985 ( .A(n479), .B(n478), .CI(n477), .CO(n472), .S(n501) );
  CMPR32X1 U986 ( .A(n482), .B(n481), .C(n480), .CO(n465), .S(n533) );
  CMPR32X1 U987 ( .A(n485), .B(n484), .C(n483), .CO(n478), .S(n532) );
  XNOR2X1 U988 ( .A(n585), .B(n596), .Y(n511) );
  NOR2X1 U989 ( .A(n1046), .B(n490), .Y(n913) );
  NOR2XL U990 ( .A(n501), .B(n500), .Y(mult_x_1_n183) );
  NAND2XL U991 ( .A(n501), .B(n500), .Y(mult_x_1_n184) );
  INVXL U992 ( .A(n1340), .Y(n502) );
  XNOR2X1 U993 ( .A(n1185), .B(A[14]), .Y(n911) );
  XNOR2X1 U994 ( .A(n908), .B(n1201), .Y(n909) );
  XNOR2X1 U995 ( .A(n916), .B(n719), .Y(n917) );
  XNOR2X1 U996 ( .A(n799), .B(n668), .Y(n516) );
  XNOR2X1 U997 ( .A(n585), .B(A[19]), .Y(n942) );
  OAI22X1 U998 ( .A0(n1077), .A1(n942), .B0(n6), .B1(n511), .Y(n923) );
  XNOR2X1 U999 ( .A(n1210), .B(n1035), .Y(n944) );
  OR2X2 U1000 ( .A(n923), .B(n922), .Y(n522) );
  XNOR2X1 U1001 ( .A(n799), .B(A[15]), .Y(n924) );
  XNOR2X1 U1002 ( .A(n669), .B(n1208), .Y(n926) );
  XNOR2X1 U1003 ( .A(n746), .B(A[25]), .Y(n918) );
  CMPR32X1 U1004 ( .A(n521), .B(n520), .C(n519), .CO(n530), .S(n961) );
  CMPR32X1 U1005 ( .A(n524), .B(n523), .C(n522), .CO(n528), .S(n960) );
  CMPR32X1 U1006 ( .A(n530), .B(n529), .C(n528), .CO(n907), .S(n954) );
  ADDFHX1 U1007 ( .A(n533), .B(n532), .CI(n531), .CO(n500), .S(n534) );
  NOR2XL U1008 ( .A(n535), .B(n534), .Y(mult_x_1_n194) );
  NAND2XL U1009 ( .A(n535), .B(n534), .Y(mult_x_1_n195) );
  NAND2XL U1010 ( .A(n157), .B(n302), .Y(n542) );
  OAI21XL U1011 ( .A0(n1159), .A1(n542), .B0(n541), .Y(n546) );
  NAND2X1 U1012 ( .A(n544), .B(n543), .Y(n545) );
  NAND2XL U1013 ( .A(n157), .B(n559), .Y(n550) );
  OAI21XL U1014 ( .A0(n1159), .A1(n550), .B0(n549), .Y(n555) );
  OAI21XL U1015 ( .A0(n1159), .A1(n557), .B0(n307), .Y(n560) );
  INVXL U1016 ( .A(n651), .Y(n564) );
  AOI21XL U1017 ( .A0(n563), .A1(n652), .B0(n564), .Y(n565) );
  XNOR2X1 U1018 ( .A(n1185), .B(A[10]), .Y(n570) );
  XNOR2X1 U1019 ( .A(n1036), .B(n1026), .Y(n624) );
  XNOR2X1 U1020 ( .A(n1036), .B(A[14]), .Y(n577) );
  OAI22X1 U1021 ( .A0(n1088), .A1(n624), .B0(n1086), .B1(n577), .Y(n611) );
  XNOR2X1 U1022 ( .A(n746), .B(n1183), .Y(n572) );
  XNOR2X1 U1023 ( .A(n746), .B(n1201), .Y(n578) );
  OAI22XL U1024 ( .A0(n180), .A1(n572), .B0(n578), .B1(n1153), .Y(n581) );
  XNOR2XL U1025 ( .A(n746), .B(n596), .Y(n627) );
  XNOR2X1 U1026 ( .A(n1044), .B(n1028), .Y(n573) );
  XNOR2X1 U1027 ( .A(n799), .B(n1035), .Y(n603) );
  XNOR2X1 U1028 ( .A(n799), .B(n745), .Y(n574) );
  XNOR2X1 U1029 ( .A(n669), .B(A[19]), .Y(n604) );
  XNOR2X1 U1030 ( .A(n669), .B(n596), .Y(n575) );
  XNOR2X1 U1031 ( .A(n908), .B(n719), .Y(n576) );
  OAI22XL U1032 ( .A0(n1056), .A1(n605), .B0(n9), .B1(n576), .Y(n606) );
  XNOR2XL U1033 ( .A(n908), .B(A[19]), .Y(n597) );
  OAI22XL U1034 ( .A0(n1056), .A1(n576), .B0(n9), .B1(n597), .Y(n592) );
  OAI22XL U1035 ( .A0(n1088), .A1(n577), .B0(n1086), .B1(n598), .Y(n591) );
  XNOR2XL U1036 ( .A(n746), .B(n1208), .Y(n599) );
  ADDHXL U1037 ( .A(n581), .B(n580), .CO(n589), .S(n610) );
  XNOR2X1 U1038 ( .A(n585), .B(n719), .Y(n943) );
  XNOR2X1 U1039 ( .A(n1210), .B(A[10]), .Y(n945) );
  CMPR32X1 U1040 ( .A(n591), .B(n590), .C(n589), .CO(n1008), .S(n615) );
  CMPR32X1 U1041 ( .A(n594), .B(n593), .C(n592), .CO(n995), .S(n616) );
  XNOR2X1 U1042 ( .A(n669), .B(n1201), .Y(n927) );
  OAI22X1 U1043 ( .A0(n1053), .A1(n595), .B0(n1051), .B1(n927), .Y(n964) );
  XNOR2XL U1044 ( .A(n916), .B(n668), .Y(n934) );
  OAI22XL U1045 ( .A0(n1088), .A1(n598), .B0(n1086), .B1(n934), .Y(n992) );
  OAI22XL U1046 ( .A0(n808), .A1(n599), .B0(n919), .B1(n1153), .Y(n938) );
  XNOR2XL U1047 ( .A(n1044), .B(n776), .Y(n600) );
  NOR2XL U1048 ( .A(n1046), .B(n600), .Y(n937) );
  CMPR22X1 U1049 ( .A(n602), .B(n601), .CO(n990), .S(n590) );
  XNOR2X1 U1050 ( .A(n799), .B(A[10]), .Y(n629) );
  XNOR2XL U1051 ( .A(n908), .B(n668), .Y(n631) );
  OAI22XL U1052 ( .A0(n1056), .A1(n631), .B0(n9), .B1(n605), .Y(n632) );
  XNOR2X1 U1053 ( .A(n1036), .B(n745), .Y(n1037) );
  XNOR2XL U1054 ( .A(n1044), .B(n772), .Y(n628) );
  XNOR2X1 U1055 ( .A(n799), .B(n920), .Y(n1047) );
  OAI22X1 U1056 ( .A0(n1049), .A1(n1047), .B0(n8), .B1(n629), .Y(n1059) );
  XNOR2X1 U1057 ( .A(n669), .B(n915), .Y(n1050) );
  OAI22X1 U1058 ( .A0(n1053), .A1(n1050), .B0(n1051), .B1(n630), .Y(n1058) );
  CMPR32X1 U1059 ( .A(n637), .B(n636), .C(n635), .CO(n638), .S(n1066) );
  CMPR32X1 U1060 ( .A(n643), .B(n642), .C(n641), .CO(n646), .S(n1069) );
  CMPR32X1 U1061 ( .A(n646), .B(n645), .C(n644), .CO(n1020), .S(n1023) );
  NOR2XL U1062 ( .A(n648), .B(n647), .Y(mult_x_1_n244) );
  NAND2XL U1063 ( .A(n648), .B(n647), .Y(mult_x_1_n245) );
  INVXL U1064 ( .A(n563), .Y(n649) );
  INVXL U1065 ( .A(n655), .Y(n657) );
  NAND2XL U1066 ( .A(n657), .B(n656), .Y(n658) );
  INVXL U1067 ( .A(n660), .Y(n662) );
  NAND2XL U1068 ( .A(n662), .B(n661), .Y(n663) );
  OAI22X1 U1069 ( .A0(n1218), .A1(n676), .B0(n1219), .B1(n667), .Y(n707) );
  NOR2XL U1070 ( .A(n1046), .B(n665), .Y(n706) );
  XNOR2XL U1071 ( .A(n1185), .B(n1028), .Y(n716) );
  OAI22XL U1072 ( .A0(n1187), .A1(n684), .B0(n5), .B1(n716), .Y(n705) );
  XNOR2X1 U1073 ( .A(n585), .B(A[10]), .Y(n697) );
  XNOR2XL U1074 ( .A(n585), .B(n1035), .Y(n717) );
  OAI22XL U1075 ( .A0(n718), .A1(n697), .B0(n6), .B1(n717), .Y(n710) );
  OAI22XL U1076 ( .A0(n1088), .A1(n682), .B0(n1086), .B1(n714), .Y(n709) );
  XNOR2X1 U1077 ( .A(n746), .B(n668), .Y(n674) );
  XNOR2X1 U1078 ( .A(n746), .B(n915), .Y(n720) );
  XNOR2X1 U1079 ( .A(n799), .B(n1030), .Y(n686) );
  XNOR2X1 U1080 ( .A(n799), .B(n776), .Y(n1048) );
  OAI22XL U1081 ( .A0(n1049), .A1(n686), .B0(n8), .B1(n1048), .Y(n1095) );
  OAI22X1 U1082 ( .A0(n1218), .A1(n667), .B0(n1219), .B1(n1079), .Y(n1094) );
  XNOR2X1 U1083 ( .A(n669), .B(A[15]), .Y(n687) );
  OAI22XL U1084 ( .A0(n180), .A1(n731), .B0(n675), .B1(n1153), .Y(n730) );
  OAI22X1 U1085 ( .A0(n673), .A1(n672), .B0(n671), .B1(n670), .Y(n729) );
  OAI22XL U1086 ( .A0(n808), .A1(n675), .B0(n674), .B1(n1040), .Y(n680) );
  XNOR2X1 U1087 ( .A(n1210), .B(n732), .Y(n677) );
  XNOR2X1 U1088 ( .A(n1036), .B(A[6]), .Y(n737) );
  OAI22X1 U1089 ( .A0(n1218), .A1(n678), .B0(n1219), .B1(n677), .Y(n741) );
  OAI22XL U1090 ( .A0(n1187), .A1(n733), .B0(n5), .B1(n685), .Y(n740) );
  CMPR32X1 U1091 ( .A(n681), .B(n680), .C(n679), .CO(n701), .S(n735) );
  XNOR2X1 U1092 ( .A(n774), .B(n1026), .Y(n689) );
  XNOR2X1 U1093 ( .A(n774), .B(A[14]), .Y(n688) );
  OAI22X1 U1094 ( .A0(n1053), .A1(n689), .B0(n1051), .B1(n688), .Y(n692) );
  OAI22XL U1095 ( .A0(n1187), .A1(n685), .B0(n5), .B1(n684), .Y(n691) );
  XNOR2X1 U1096 ( .A(n799), .B(A[6]), .Y(n695) );
  XNOR2X1 U1097 ( .A(n777), .B(n745), .Y(n694) );
  XNOR2X1 U1098 ( .A(n774), .B(n745), .Y(n739) );
  XNOR2X1 U1099 ( .A(n799), .B(n772), .Y(n738) );
  XNOR2X1 U1100 ( .A(n799), .B(n1028), .Y(n696) );
  XNOR2X1 U1101 ( .A(n585), .B(n920), .Y(n698) );
  OAI22XL U1102 ( .A0(n1049), .A1(n696), .B0(n8), .B1(n695), .Y(n703) );
  CMPR32X1 U1103 ( .A(n704), .B(n703), .C(n702), .CO(n726), .S(n760) );
  CMPR32X1 U1104 ( .A(n707), .B(n706), .C(n705), .CO(n1140), .S(n725) );
  CMPR32X1 U1105 ( .A(n710), .B(n709), .C(n708), .CO(n1139), .S(n724) );
  CMPR32X1 U1106 ( .A(n713), .B(n712), .C(n711), .CO(n1125), .S(n699) );
  XNOR2X1 U1107 ( .A(n1036), .B(A[10]), .Y(n1087) );
  OAI22XL U1108 ( .A0(n1187), .A1(n716), .B0(n5), .B1(n1081), .Y(n1114) );
  XNOR2X1 U1109 ( .A(n585), .B(n745), .Y(n1076) );
  OAI22XL U1110 ( .A0(n718), .A1(n717), .B0(n6), .B1(n1076), .Y(n1122) );
  XNOR2XL U1111 ( .A(n746), .B(n719), .Y(n1042) );
  ADDHXL U1112 ( .A(n723), .B(n722), .CO(n1120), .S(n708) );
  XNOR2X1 U1113 ( .A(n777), .B(A[10]), .Y(n743) );
  OAI22X1 U1114 ( .A0(n728), .A1(n743), .B0(n9), .B1(n727), .Y(n768) );
  ADDHXL U1115 ( .A(n730), .B(n729), .CO(n736), .S(n767) );
  ADDFHX1 U1116 ( .A(n736), .B(n735), .CI(n734), .CO(n752), .S(n783) );
  XNOR2X1 U1117 ( .A(n1036), .B(n1028), .Y(n773) );
  XNOR2X1 U1118 ( .A(n799), .B(n1043), .Y(n800) );
  OAI22XL U1119 ( .A0(n1049), .A1(n800), .B0(n8), .B1(n738), .Y(n780) );
  XNOR2XL U1120 ( .A(n774), .B(n1035), .Y(n775) );
  OAI22XL U1121 ( .A0(n1053), .A1(n775), .B0(n1051), .B1(n739), .Y(n779) );
  XNOR2X1 U1122 ( .A(n585), .B(n1030), .Y(n795) );
  XNOR2X1 U1123 ( .A(n746), .B(n745), .Y(n806) );
  OAI22X1 U1124 ( .A0(n808), .A1(n806), .B0(n747), .B1(n1153), .Y(n805) );
  OAI22X1 U1125 ( .A0(n1205), .A1(n749), .B0(n5), .B1(n748), .Y(n804) );
  NAND2XL U1126 ( .A(n754), .B(n753), .Y(mult_x_1_n282) );
  CMPR32X1 U1127 ( .A(n762), .B(n761), .C(n760), .CO(n750), .S(n791) );
  XNOR2X1 U1128 ( .A(n1036), .B(n772), .Y(n832) );
  XNOR2XL U1129 ( .A(n774), .B(A[10]), .Y(n813) );
  OAI22XL U1130 ( .A0(n1053), .A1(n813), .B0(n1051), .B1(n775), .Y(n830) );
  NOR2XL U1131 ( .A(n786), .B(n785), .Y(mult_x_1_n286) );
  NAND2XL U1132 ( .A(n786), .B(n785), .Y(mult_x_1_n287) );
  INVX1 U1133 ( .A(n1356), .Y(n868) );
  NAND2XL U1134 ( .A(n13), .B(n1349), .Y(n787) );
  XNOR2X1 U1135 ( .A(n585), .B(A[6]), .Y(n811) );
  XNOR2X1 U1136 ( .A(n799), .B(n798), .Y(n809) );
  CMPR32X1 U1137 ( .A(n803), .B(n802), .C(n801), .CO(n792), .S(n839) );
  NOR2XL U1138 ( .A(n821), .B(n820), .Y(mult_x_1_n292) );
  NAND2XL U1139 ( .A(n821), .B(n820), .Y(mult_x_1_n293) );
  CMPR32X1 U1140 ( .A(n831), .B(n830), .C(n829), .CO(n824), .S(n854) );
  OAI22X1 U1141 ( .A0(n1088), .A1(n833), .B0(n1086), .B1(n832), .Y(n877) );
  CMPR32X1 U1142 ( .A(n849), .B(n848), .C(n847), .CO(n882), .S(n886) );
  CMPR32X1 U1143 ( .A(n852), .B(n851), .C(n850), .CO(n841), .S(n881) );
  CMPR32X1 U1144 ( .A(n855), .B(n854), .C(n853), .CO(n860), .S(n1160) );
  NAND2XL U1145 ( .A(n1156), .B(n869), .Y(mult_x_1_n295) );
  INVXL U1146 ( .A(n1155), .Y(n866) );
  XOR2X1 U1147 ( .A(n1357), .B(n1353), .Y(PRODUCT[13]) );
  XNOR2X1 U1148 ( .A(n1320), .B(n1354), .Y(PRODUCT[12]) );
  OAI21XL U1149 ( .A0(n871), .A1(n891), .B0(n870), .Y(n872) );
  INVXL U1150 ( .A(n1172), .Y(mult_x_1_n321) );
  CMPR32X1 U1151 ( .A(n880), .B(n879), .C(n878), .CO(n1164), .S(n884) );
  ADDFHX1 U1152 ( .A(n883), .B(n882), .CI(n881), .CO(n1161), .S(n1163) );
  AOI21XL U1153 ( .A0(mult_x_1_n321), .A1(n887), .B0(n1169), .Y(mult_x_1_n316)
         );
  INVXL U1154 ( .A(n890), .Y(n892) );
  NAND2XL U1155 ( .A(n892), .B(n891), .Y(n893) );
  XOR2X1 U1156 ( .A(n894), .B(n893), .Y(n1391) );
  XOR2X1 U1157 ( .A(n900), .B(n899), .Y(n1392) );
  XNOR2X1 U1158 ( .A(n908), .B(n1183), .Y(n928) );
  XNOR2X1 U1159 ( .A(n1044), .B(A[10]), .Y(n910) );
  NOR2XL U1160 ( .A(n1046), .B(n910), .Y(n949) );
  OAI22XL U1161 ( .A0(n1187), .A1(n946), .B0(n5), .B1(n911), .Y(n948) );
  XNOR2X1 U1162 ( .A(n916), .B(n915), .Y(n933) );
  OAI22X1 U1163 ( .A0(n180), .A1(n919), .B0(n918), .B1(n1153), .Y(n936) );
  XNOR2XL U1164 ( .A(n1044), .B(n920), .Y(n921) );
  CMPR32X1 U1165 ( .A(n932), .B(n931), .C(n930), .CO(n962), .S(n973) );
  OAI22XL U1166 ( .A0(n1088), .A1(n934), .B0(n1086), .B1(n933), .Y(n971) );
  ADDHXL U1167 ( .A(n938), .B(n937), .CO(n969), .S(n991) );
  OAI22X1 U1168 ( .A0(n1077), .A1(n943), .B0(n6), .B1(n942), .Y(n989) );
  OAI22X1 U1169 ( .A0(n1218), .A1(n945), .B0(n1219), .B1(n944), .Y(n988) );
  OAI22XL U1170 ( .A0(n1187), .A1(n947), .B0(n5), .B1(n946), .Y(n987) );
  CMPR32X1 U1171 ( .A(n950), .B(n949), .C(n948), .CO(n941), .S(n976) );
  CMPR32X1 U1172 ( .A(n953), .B(n952), .C(n951), .CO(n939), .S(n975) );
  CMPR32X1 U1173 ( .A(n968), .B(n967), .C(n966), .CO(n974), .S(n1000) );
  CMPR32X1 U1174 ( .A(n971), .B(n970), .C(n969), .CO(n972), .S(n999) );
  ADDFHX1 U1175 ( .A(n986), .B(n985), .CI(n984), .CO(n998), .S(n1009) );
  CMPR32X1 U1176 ( .A(n992), .B(n990), .C(n991), .CO(n996), .S(n993) );
  CMPR32X1 U1177 ( .A(n995), .B(n994), .C(n993), .CO(n1016), .S(n1011) );
  CMPR32X1 U1178 ( .A(n998), .B(n997), .C(n996), .CO(n1007), .S(n1015) );
  ADDFX2 U1179 ( .A(n1010), .B(n1009), .CI(n1008), .CO(n1019), .S(n1012) );
  ADDFHX1 U1180 ( .A(n1022), .B(n1021), .CI(n1020), .CO(mult_x_1_n569), .S(
        n648) );
  ADDFHX1 U1181 ( .A(n1025), .B(n1024), .CI(n1023), .CO(n647), .S(
        mult_x_1_n586) );
  OAI22XL U1182 ( .A0(n1187), .A1(n1080), .B0(n5), .B1(n1031), .Y(n1082) );
  OAI22XL U1183 ( .A0(n1088), .A1(n1085), .B0(n1086), .B1(n1037), .Y(n1062) );
  OAI22XL U1184 ( .A0(n808), .A1(n1042), .B0(n1041), .B1(n1040), .Y(n1090) );
  XNOR2XL U1185 ( .A(n1044), .B(n1043), .Y(n1045) );
  NOR2XL U1186 ( .A(n1046), .B(n1045), .Y(n1089) );
  OAI22X1 U1187 ( .A0(n1049), .A1(n1048), .B0(n8), .B1(n1047), .Y(n1098) );
  OAI22X1 U1188 ( .A0(n1053), .A1(n1052), .B0(n1051), .B1(n1050), .Y(n1097) );
  OAI22X1 U1189 ( .A0(n1056), .A1(n1055), .B0(n9), .B1(n1054), .Y(n1096) );
  CMPR32X1 U1190 ( .A(n1068), .B(n1067), .C(n1066), .CO(n1071), .S(n1108) );
  CMPR32X1 U1191 ( .A(n1071), .B(n1070), .C(n1069), .CO(n1024), .S(n1072) );
  CMPR32X1 U1192 ( .A(n1074), .B(n1073), .C(n1072), .CO(mult_x_1_n601), .S(
        mult_x_1_n602) );
  OAI22X2 U1193 ( .A0(n1218), .A1(n1079), .B0(n1219), .B1(n1078), .Y(n1118) );
  OAI22XL U1194 ( .A0(n1088), .A1(n1087), .B0(n1086), .B1(n1085), .Y(n1101) );
  ADDHXL U1195 ( .A(n1090), .B(n1089), .CO(n1060), .S(n1100) );
  CMPR32X1 U1196 ( .A(n1098), .B(n1097), .C(n1096), .CO(n1107), .S(n1130) );
  CMPR32X1 U1197 ( .A(n1101), .B(n66), .C(n1099), .CO(n1102), .S(n1129) );
  CMPR32X1 U1198 ( .A(n1104), .B(n1103), .C(n1102), .CO(n1113), .S(n1133) );
  ADDFHX1 U1199 ( .A(n1110), .B(n1109), .CI(n1108), .CO(n1073), .S(n1111) );
  ADDFHX1 U1200 ( .A(n1113), .B(n1112), .CI(n1111), .CO(mult_x_1_n617), .S(
        mult_x_1_n618) );
  CMPR32X1 U1201 ( .A(n1116), .B(n1115), .C(n1114), .CO(n1128), .S(n1124) );
  ADDFX2 U1202 ( .A(n1128), .B(n1127), .CI(n1126), .CO(n1137), .S(n1145) );
  CMPR32X1 U1203 ( .A(n1131), .B(n1130), .C(n1129), .CO(n1134), .S(n1144) );
  CMPR32X1 U1204 ( .A(n1140), .B(n1139), .C(n1138), .CO(n1149), .S(n1152) );
  CMPR32X1 U1205 ( .A(n1149), .B(n1148), .C(n1147), .CO(mult_x_1_n649), .S(
        mult_x_1_n650) );
  NAND2XL U1206 ( .A(n1156), .B(n1155), .Y(mult_x_1_n83) );
  NAND2XL U1207 ( .A(n150), .B(n314), .Y(n1158) );
  ADDFHX1 U1208 ( .A(n1162), .B(n1161), .CI(n1160), .CO(n862), .S(n1167) );
  NAND2XL U1209 ( .A(n57), .B(n887), .Y(n1171) );
  NAND2XL U1210 ( .A(n1167), .B(n1166), .Y(n1173) );
  INVXL U1211 ( .A(n1173), .Y(n1168) );
  AOI21XL U1212 ( .A0(n57), .A1(n1169), .B0(n1168), .Y(n1170) );
  OAI21XL U1213 ( .A0(n1172), .A1(n1171), .B0(n1170), .Y(mult_x_1_n309) );
  CMPR32X1 U1214 ( .A(n1178), .B(n1177), .C(n1176), .CO(n1192), .S(n1174) );
  CMPR32X1 U1215 ( .A(n1181), .B(n1180), .C(n1179), .CO(n1196), .S(n1178) );
  XNOR2X1 U1216 ( .A(n1210), .B(n1208), .Y(n1197) );
  OAI22X1 U1217 ( .A0(n1187), .A1(n1186), .B0(n5), .B1(n1203), .Y(n1214) );
  CMPR32X1 U1218 ( .A(n1190), .B(n1189), .C(n1188), .CO(n1194), .S(n1177) );
  NAND2XL U1219 ( .A(n887), .B(n1193), .Y(mult_x_1_n86) );
  CMPR32X1 U1220 ( .A(n1196), .B(n1195), .C(n1194), .CO(n1207), .S(n1191) );
  CMPR32X1 U1221 ( .A(n1200), .B(n1199), .C(n1198), .CO(n1228), .S(n1195) );
  CMPR32X1 U1222 ( .A(n1214), .B(n1213), .C(n1212), .CO(n1230), .S(n1227) );
  OAI2BB1X1 U1223 ( .A0N(n1219), .A1N(n1218), .B0(n1217), .Y(n1220) );
  XOR3X2 U1224 ( .A(n1222), .B(n1221), .C(n1220), .Y(n1223) );
  CMPR32X1 U1225 ( .A(n1229), .B(n1228), .C(n1227), .CO(n1234), .S(n1206) );
  CMPR32X1 U1226 ( .A(n1232), .B(n1231), .C(n1230), .CO(n1224), .S(n1233) );
  OAI21XL U1227 ( .A0(n1240), .A1(n1335), .B0(n1239), .Y(n1300) );
  OAI21XL U1228 ( .A0(n1307), .A1(n1244), .B0(n1243), .Y(n1246) );
  OAI21XL U1229 ( .A0(n1307), .A1(n1250), .B0(n1249), .Y(n1253) );
  OAI21XL U1230 ( .A0(n1267), .A1(n1264), .B0(n1265), .Y(n1259) );
  INVXL U1231 ( .A(n1255), .Y(n1257) );
  OAI21XL U1232 ( .A0(n1326), .A1(n1329), .B0(n1327), .Y(n1273) );
  OAI21XL U1233 ( .A0(n1307), .A1(n1261), .B0(n1260), .Y(n1263) );
  OAI21XL U1234 ( .A0(n1307), .A1(n1278), .B0(n1277), .Y(n1281) );
  XOR2XL U1235 ( .A(n1290), .B(n1289), .Y(n1398) );
  XNOR2XL U1236 ( .A(n1293), .B(n1292), .Y(n1397) );
  OAI21XL U1237 ( .A0(n1297), .A1(n1322), .B0(n1323), .Y(n1298) );
  OAI21XL U1238 ( .A0(n1303), .A1(n1302), .B0(n1301), .Y(n1304) );
  OAI21XL U1239 ( .A0(n1307), .A1(n1306), .B0(n1305), .Y(n1308) );
  XNOR2XL U1240 ( .A(n1308), .B(n1321), .Y(PRODUCT[40]) );
  XNOR2XL U1241 ( .A(n1312), .B(n1311), .Y(n1399) );
  XOR2XL U1242 ( .A(n1317), .B(n1316), .Y(n1396) );
endmodule


module FFT2048_DW02_mult_2_stage_J1_8 ( A, B, TC, CLK, PRODUCT );
  input [25:0] A;
  input [16:0] B;
  output [42:0] PRODUCT;
  input TC, CLK;
  wire   n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, mult_x_1_n633, mult_x_1_n618, mult_x_1_n617,
         mult_x_1_n602, mult_x_1_n601, mult_x_1_n586, mult_x_1_n569,
         mult_x_1_n554, mult_x_1_n537, mult_x_1_n522, mult_x_1_n316,
         mult_x_1_n309, mult_x_1_n307, mult_x_1_n306, mult_x_1_n296,
         mult_x_1_n295, mult_x_1_n293, mult_x_1_n292, mult_x_1_n287,
         mult_x_1_n286, mult_x_1_n282, mult_x_1_n281, mult_x_1_n277,
         mult_x_1_n276, mult_x_1_n274, mult_x_1_n273, mult_x_1_n245,
         mult_x_1_n244, mult_x_1_n227, mult_x_1_n226, mult_x_1_n207,
         mult_x_1_n206, mult_x_1_n198, mult_x_1_n197, mult_x_1_n195,
         mult_x_1_n194, mult_x_1_n184, mult_x_1_n183, mult_x_1_n177,
         mult_x_1_n176, mult_x_1_n170, mult_x_1_n169, mult_x_1_n161,
         mult_x_1_n160, mult_x_1_n152, mult_x_1_n151, mult_x_1_n137,
         mult_x_1_n136, mult_x_1_n130, mult_x_1_n129, mult_x_1_n121,
         mult_x_1_n120, mult_x_1_n110, mult_x_1_n109, mult_x_1_n85,
         mult_x_1_n84, mult_x_1_n83, mult_x_1_n58, n5, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299;

  DFFHQXL mult_x_1_clk_r_REG9_S1 ( .D(mult_x_1_n195), .CK(CLK), .Q(n1264) );
  DFFHQX4 mult_x_1_clk_r_REG38_S1 ( .D(mult_x_1_n633), .CK(CLK), .Q(n1299) );
  DFFHQX4 mult_x_1_clk_r_REG37_S1 ( .D(mult_x_1_n618), .CK(CLK), .Q(n1298) );
  DFFHQX4 mult_x_1_clk_r_REG36_S1 ( .D(mult_x_1_n617), .CK(CLK), .Q(n1297) );
  DFFHQX4 mult_x_1_clk_r_REG35_S1 ( .D(mult_x_1_n602), .CK(CLK), .Q(n1296) );
  DFFHQX4 mult_x_1_clk_r_REG34_S1 ( .D(mult_x_1_n601), .CK(CLK), .Q(n1295) );
  DFFHQX4 mult_x_1_clk_r_REG33_S1 ( .D(mult_x_1_n586), .CK(CLK), .Q(n1294) );
  DFFHQX4 mult_x_1_clk_r_REG30_S1 ( .D(mult_x_1_n569), .CK(CLK), .Q(n1293) );
  DFFHQX4 mult_x_1_clk_r_REG0_S1 ( .D(mult_x_1_n554), .CK(CLK), .Q(n1292) );
  DFFHQX4 mult_x_1_clk_r_REG3_S1 ( .D(mult_x_1_n537), .CK(CLK), .Q(n1291) );
  DFFHQX4 mult_x_1_clk_r_REG4_S1 ( .D(mult_x_1_n522), .CK(CLK), .Q(n1290) );
  DFFHQX4 mult_x_1_clk_r_REG56_S1 ( .D(mult_x_1_n309), .CK(CLK), .Q(n1288) );
  DFFHQX4 mult_x_1_clk_r_REG50_S1 ( .D(mult_x_1_n296), .CK(CLK), .Q(n1287) );
  DFFHQXL mult_x_1_clk_r_REG49_S1 ( .D(mult_x_1_n83), .CK(CLK), .Q(n1284) );
  DFFHQX4 mult_x_1_clk_r_REG51_S1 ( .D(mult_x_1_n295), .CK(CLK), .Q(n1283) );
  DFFHQX4 mult_x_1_clk_r_REG48_S1 ( .D(mult_x_1_n292), .CK(CLK), .Q(n1281) );
  DFFHQX4 mult_x_1_clk_r_REG45_S1 ( .D(mult_x_1_n287), .CK(CLK), .Q(n1280) );
  DFFHQX4 mult_x_1_clk_r_REG46_S1 ( .D(mult_x_1_n286), .CK(CLK), .Q(n1279) );
  DFFHQX4 mult_x_1_clk_r_REG44_S1 ( .D(mult_x_1_n281), .CK(CLK), .Q(n1277) );
  DFFHQX4 mult_x_1_clk_r_REG41_S1 ( .D(mult_x_1_n277), .CK(CLK), .Q(n1276) );
  DFFHQX4 mult_x_1_clk_r_REG42_S1 ( .D(mult_x_1_n276), .CK(CLK), .Q(n1275) );
  DFFHQX4 mult_x_1_clk_r_REG40_S1 ( .D(mult_x_1_n273), .CK(CLK), .Q(n1273) );
  DFFHQXL mult_x_1_clk_r_REG31_S1 ( .D(mult_x_1_n245), .CK(CLK), .Q(n1272) );
  DFFHQXL mult_x_1_clk_r_REG5_S1 ( .D(mult_x_1_n207), .CK(CLK), .Q(n1268) );
  DFFHQXL clk_r_REG57_S1 ( .D(n1313), .CK(CLK), .Q(PRODUCT[12]) );
  DFFHQXL clk_r_REG59_S1 ( .D(n1314), .CK(CLK), .Q(PRODUCT[11]) );
  DFFHQXL mult_x_1_clk_r_REG13_S1 ( .D(mult_x_1_n177), .CK(CLK), .Q(n1260) );
  DFFHQXL clk_r_REG61_S1 ( .D(n1316), .CK(CLK), .Q(PRODUCT[9]) );
  DFFHQXL mult_x_1_clk_r_REG11_S1 ( .D(mult_x_1_n184), .CK(CLK), .Q(n1262) );
  DFFHQXL mult_x_1_clk_r_REG17_S1 ( .D(mult_x_1_n161), .CK(CLK), .Q(n1256) );
  DFFHQXL mult_x_1_clk_r_REG15_S1 ( .D(mult_x_1_n170), .CK(CLK), .Q(n1258) );
  DFFHQXL clk_r_REG60_S1 ( .D(n1315), .CK(CLK), .Q(PRODUCT[10]) );
  DFFHQXL mult_x_1_clk_r_REG1_S1 ( .D(mult_x_1_n227), .CK(CLK), .Q(n1270) );
  DFFHQX4 mult_x_1_clk_r_REG47_S1 ( .D(mult_x_1_n293), .CK(CLK), .Q(n1282) );
  DFFHQXL clk_r_REG62_S1 ( .D(n1317), .CK(CLK), .Q(PRODUCT[8]) );
  DFFHQXL clk_r_REG64_S1 ( .D(n1319), .CK(CLK), .Q(PRODUCT[6]) );
  DFFHQXL clk_r_REG66_S1 ( .D(n1321), .CK(CLK), .Q(PRODUCT[4]) );
  DFFHQXL clk_r_REG69_S1 ( .D(n1324), .CK(CLK), .Q(PRODUCT[1]) );
  DFFHQXL clk_r_REG70_S1 ( .D(n1325), .CK(CLK), .Q(PRODUCT[0]) );
  DFFHQXL mult_x_1_clk_r_REG58_S1 ( .D(mult_x_1_n316), .CK(CLK), .Q(n1289) );
  DFFHQXL mult_x_1_clk_r_REG52_S1 ( .D(mult_x_1_n84), .CK(CLK), .Q(n1285) );
  DFFHQXL mult_x_1_clk_r_REG7_S1 ( .D(mult_x_1_n198), .CK(CLK), .Q(n1266) );
  DFFHQXL mult_x_1_clk_r_REG10_S1 ( .D(mult_x_1_n194), .CK(CLK), .Q(n1263) );
  DFFHQXL mult_x_1_clk_r_REG19_S1 ( .D(mult_x_1_n152), .CK(CLK), .Q(n1254) );
  DFFHQXL mult_x_1_clk_r_REG21_S1 ( .D(mult_x_1_n137), .CK(CLK), .Q(n1252) );
  DFFHQXL mult_x_1_clk_r_REG23_S1 ( .D(mult_x_1_n130), .CK(CLK), .Q(n1250) );
  DFFHQXL mult_x_1_clk_r_REG24_S1 ( .D(mult_x_1_n129), .CK(CLK), .Q(n1249) );
  DFFHQXL mult_x_1_clk_r_REG25_S1 ( .D(mult_x_1_n121), .CK(CLK), .Q(n1248) );
  DFFHQXL mult_x_1_clk_r_REG26_S1 ( .D(mult_x_1_n120), .CK(CLK), .Q(n1247) );
  DFFHQXL mult_x_1_clk_r_REG27_S1 ( .D(mult_x_1_n110), .CK(CLK), .Q(n1246) );
  DFFHQXL mult_x_1_clk_r_REG28_S1 ( .D(mult_x_1_n109), .CK(CLK), .Q(n1245) );
  DFFHQXL mult_x_1_clk_r_REG29_S1 ( .D(mult_x_1_n58), .CK(CLK), .Q(n1244) );
  DFFHQXL mult_x_1_clk_r_REG53_S1 ( .D(mult_x_1_n307), .CK(CLK), .Q(n1243) );
  DFFHQXL mult_x_1_clk_r_REG54_S1 ( .D(mult_x_1_n306), .CK(CLK), .Q(n1242) );
  DFFHQXL mult_x_1_clk_r_REG8_S1 ( .D(mult_x_1_n197), .CK(CLK), .Q(n1265) );
  DFFHQXL clk_r_REG68_S1 ( .D(n1323), .CK(CLK), .Q(PRODUCT[2]) );
  DFFHQXL clk_r_REG67_S1 ( .D(n1322), .CK(CLK), .Q(PRODUCT[3]) );
  DFFHQXL clk_r_REG65_S1 ( .D(n1320), .CK(CLK), .Q(PRODUCT[5]) );
  DFFHQXL clk_r_REG63_S1 ( .D(n1318), .CK(CLK), .Q(PRODUCT[7]) );
  DFFHQXL mult_x_1_clk_r_REG22_S1 ( .D(mult_x_1_n136), .CK(CLK), .Q(n1251) );
  DFFHQXL mult_x_1_clk_r_REG20_S1 ( .D(mult_x_1_n151), .CK(CLK), .Q(n1253) );
  DFFHQXL mult_x_1_clk_r_REG18_S1 ( .D(mult_x_1_n160), .CK(CLK), .Q(n1255) );
  DFFHQXL mult_x_1_clk_r_REG12_S1 ( .D(mult_x_1_n183), .CK(CLK), .Q(n1261) );
  DFFHQXL mult_x_1_clk_r_REG16_S1 ( .D(mult_x_1_n169), .CK(CLK), .Q(n1257) );
  DFFHQXL mult_x_1_clk_r_REG14_S1 ( .D(mult_x_1_n176), .CK(CLK), .Q(n1259) );
  DFFHQX2 mult_x_1_clk_r_REG43_S1 ( .D(mult_x_1_n282), .CK(CLK), .Q(n1278) );
  DFFHQXL mult_x_1_clk_r_REG55_S1 ( .D(mult_x_1_n85), .CK(CLK), .Q(n1286) );
  DFFHQX1 mult_x_1_clk_r_REG39_S1 ( .D(mult_x_1_n274), .CK(CLK), .Q(n1274) );
  DFFHQX1 mult_x_1_clk_r_REG32_S1 ( .D(mult_x_1_n244), .CK(CLK), .Q(n1271) );
  DFFHQX1 mult_x_1_clk_r_REG6_S1 ( .D(mult_x_1_n206), .CK(CLK), .Q(n1267) );
  DFFHQX2 mult_x_1_clk_r_REG2_S1 ( .D(mult_x_1_n226), .CK(CLK), .Q(n1269) );
  ADDFHX1 U1 ( .A(n1021), .B(n1020), .CI(n1019), .CO(n382), .S(mult_x_1_n522)
         );
  ADDFHX1 U2 ( .A(n1027), .B(n1026), .CI(n1025), .CO(n459), .S(mult_x_1_n554)
         );
  ADDFHX1 U3 ( .A(n653), .B(n652), .CI(n651), .CO(n646), .S(n685) );
  ADDFHX1 U4 ( .A(n693), .B(n692), .CI(n691), .CO(n684), .S(n722) );
  ADDFHX2 U5 ( .A(n428), .B(n427), .CI(n426), .CO(n1020), .S(n1022) );
  ADDFHX2 U6 ( .A(n502), .B(n501), .CI(n500), .CO(n1026), .S(n1028) );
  ADDFHX2 U7 ( .A(n683), .B(n682), .CI(n681), .CO(n652), .S(n691) );
  ADDFHX2 U8 ( .A(n458), .B(n457), .CI(n456), .CO(n1023), .S(n1025) );
  ADDFHX1 U9 ( .A(n327), .B(n326), .CI(n325), .CO(n320), .S(n340) );
  ADDFHX1 U10 ( .A(n280), .B(n279), .CI(n278), .CO(n282), .S(n307) );
  ADDFHX2 U11 ( .A(n720), .B(n719), .CI(n718), .CO(n692), .S(n724) );
  ADDFX2 U12 ( .A(n324), .B(n323), .CI(n322), .CO(n304), .S(n341) );
  CMPR32X1 U13 ( .A(n455), .B(n454), .C(n453), .CO(n458), .S(n500) );
  CMPR32X1 U14 ( .A(n642), .B(n641), .C(n640), .CO(n645), .S(n681) );
  ADDFX2 U15 ( .A(n496), .B(n495), .CI(n494), .CO(n1030), .S(n530) );
  ADDFX2 U16 ( .A(n572), .B(n571), .CI(n570), .CO(n1072), .S(n644) );
  ADDFHX1 U17 ( .A(n821), .B(n820), .CI(n819), .CO(n824), .S(n823) );
  ADDFHX1 U18 ( .A(n818), .B(n817), .CI(n816), .CO(n776), .S(n825) );
  CMPR32X1 U19 ( .A(n121), .B(n120), .C(n119), .CO(n303), .S(n137) );
  CMPR32X1 U20 ( .A(n271), .B(n270), .C(n269), .CO(n324), .S(n301) );
  CMPR32X1 U21 ( .A(n114), .B(n113), .C(n112), .CO(n298), .S(n138) );
  CMPR32X1 U22 ( .A(n268), .B(n267), .C(n266), .CO(n295), .S(n302) );
  OAI22XL U23 ( .A0(n1121), .A1(n265), .B0(n5), .B1(n264), .Y(n296) );
  ADDFHX1 U24 ( .A(n696), .B(n695), .CI(n694), .CO(n682), .S(n726) );
  ADDFX2 U25 ( .A(n528), .B(n527), .CI(n526), .CO(n531), .S(n1052) );
  ADDFHX1 U26 ( .A(n479), .B(n478), .CI(n477), .CO(n452), .S(n495) );
  ADDFHX1 U27 ( .A(n995), .B(n994), .CI(n993), .CO(n850), .S(n1000) );
  ADDFX2 U28 ( .A(n1051), .B(n1050), .CI(n1049), .CO(n1054), .S(n1064) );
  ADDFHX1 U29 ( .A(n1036), .B(n1035), .CI(n1034), .CO(n1048), .S(n1059) );
  ADDFHX1 U30 ( .A(n594), .B(n593), .CI(n592), .CO(n1060), .S(n571) );
  ADDFHX1 U31 ( .A(n848), .B(n847), .CI(n846), .CO(n832), .S(n993) );
  ADDFHX1 U32 ( .A(n781), .B(n780), .CI(n779), .CO(n773), .S(n821) );
  CMPR32X1 U33 ( .A(n815), .B(n814), .C(n813), .CO(n820), .S(n831) );
  NOR2BX2 U34 ( .AN(A[0]), .B(n698), .Y(n738) );
  BUFX3 U35 ( .A(B[16]), .Y(n1141) );
  ADDFHX1 U36 ( .A(n973), .B(n972), .CI(n971), .CO(n994), .S(n996) );
  ADDFHX1 U37 ( .A(n982), .B(n981), .CI(n980), .CO(n997), .S(n983) );
  CLKBUFX8 U38 ( .A(n93), .Y(n1121) );
  CMPR32X1 U39 ( .A(n976), .B(n975), .C(n974), .CO(n972), .S(n985) );
  ADDFX2 U40 ( .A(n950), .B(n949), .CI(n948), .CO(n957), .S(n955) );
  BUFX3 U41 ( .A(n171), .Y(n5) );
  NAND2X2 U42 ( .A(n106), .B(n62), .Y(n575) );
  NAND2X4 U43 ( .A(n101), .B(n410), .Y(n409) );
  BUFX3 U44 ( .A(n410), .Y(n837) );
  ADDFHX1 U45 ( .A(n944), .B(n943), .CI(n942), .CO(n949), .S(n951) );
  ADDHXL U46 ( .A(n923), .B(n922), .CO(n945), .S(n953) );
  BUFX3 U47 ( .A(n916), .Y(n921) );
  BUFX3 U48 ( .A(n933), .Y(n930) );
  BUFX3 U49 ( .A(n938), .Y(n855) );
  BUFX3 U50 ( .A(n670), .Y(n8) );
  BUFX4 U51 ( .A(n100), .Y(n932) );
  CLKBUFX8 U52 ( .A(B[9]), .Y(n928) );
  NAND2X1 U53 ( .A(n94), .B(n45), .Y(n916) );
  XNOR2X1 U54 ( .A(B[6]), .B(B[5]), .Y(n556) );
  XNOR2X1 U55 ( .A(B[4]), .B(B[3]), .Y(n94) );
  NAND2X1 U56 ( .A(n534), .B(n83), .Y(n462) );
  NOR2X2 U57 ( .A(n547), .B(n542), .Y(n534) );
  OAI21XL U58 ( .A0(n1273), .A1(n1276), .B0(n1274), .Y(n19) );
  NOR2X2 U59 ( .A(n1293), .B(n1292), .Y(n463) );
  OAI21X1 U60 ( .A0(n1277), .A1(n1280), .B0(n1278), .Y(n553) );
  NOR2X1 U61 ( .A(n1291), .B(n1290), .Y(n348) );
  OAI21X2 U62 ( .A0(n542), .A1(n548), .B0(n543), .Y(n535) );
  NOR2X1 U63 ( .A(n538), .B(n1271), .Y(n15) );
  NOR2BX1 U64 ( .AN(n1272), .B(n15), .Y(n14) );
  NOR2X2 U65 ( .A(n463), .B(n1269), .Y(n347) );
  AOI21XL U66 ( .A0(n85), .A1(n385), .B0(n84), .Y(n82) );
  XNOR2XL U67 ( .A(n926), .B(A[10]), .Y(n838) );
  XNOR2XL U68 ( .A(n442), .B(A[6]), .Y(n841) );
  XNOR2XL U69 ( .A(n926), .B(A[13]), .Y(n715) );
  XNOR2XL U70 ( .A(B[3]), .B(A[0]), .Y(n881) );
  XNOR2XL U71 ( .A(n1141), .B(A[16]), .Y(n184) );
  XNOR2XL U72 ( .A(n1123), .B(A[1]), .Y(n664) );
  XNOR2XL U73 ( .A(n1107), .B(A[3]), .Y(n666) );
  XNOR2XL U74 ( .A(B[1]), .B(A[22]), .Y(n438) );
  XNOR2XL U75 ( .A(n926), .B(A[19]), .Y(n584) );
  XNOR2XL U76 ( .A(n802), .B(A[8]), .Y(n578) );
  XNOR2XL U77 ( .A(n442), .B(A[25]), .Y(n248) );
  XNOR2XL U78 ( .A(n1209), .B(n1208), .Y(PRODUCT[39]) );
  XNOR2XL U79 ( .A(n1123), .B(A[20]), .Y(n202) );
  XNOR2XL U80 ( .A(n802), .B(A[22]), .Y(n223) );
  XNOR2XL U81 ( .A(n442), .B(A[23]), .Y(n105) );
  XNOR2XL U82 ( .A(n1123), .B(A[9]), .Y(n430) );
  XNOR2XL U83 ( .A(n1107), .B(A[5]), .Y(n615) );
  ADDFX2 U84 ( .A(n297), .B(n296), .CI(n295), .CO(n305), .S(n327) );
  ADDFX2 U85 ( .A(n797), .B(n796), .CI(n795), .CO(n817), .S(n819) );
  XNOR2XL U86 ( .A(n1182), .B(n1181), .Y(n1318) );
  XOR2XL U87 ( .A(n1191), .B(n1190), .Y(n1319) );
  XOR2XL U88 ( .A(n1011), .B(n1010), .Y(n1315) );
  XOR2X1 U89 ( .A(n1018), .B(n1017), .Y(n1316) );
  NAND2XL U90 ( .A(n685), .B(n684), .Y(mult_x_1_n277) );
  INVX1 U91 ( .A(n1001), .Y(n1076) );
  XNOR2X1 U92 ( .A(n1176), .B(n1175), .Y(n1317) );
  INVX1 U93 ( .A(n957), .Y(n22) );
  NOR2X1 U94 ( .A(n1143), .B(n562), .Y(n618) );
  NOR2X1 U95 ( .A(n1143), .B(n183), .Y(n200) );
  NOR2X1 U96 ( .A(n1143), .B(n1118), .Y(n1126) );
  NOR2X1 U97 ( .A(n1143), .B(n1122), .Y(n1140) );
  NOR2X1 U98 ( .A(n1143), .B(n247), .Y(n274) );
  NOR2X1 U99 ( .A(n1143), .B(n184), .Y(n234) );
  NOR2X1 U100 ( .A(n1143), .B(n226), .Y(n252) );
  XNOR2XL U101 ( .A(n1141), .B(A[21]), .Y(n1106) );
  INVXL U102 ( .A(n946), .Y(n25) );
  INVX1 U103 ( .A(n552), .Y(n7) );
  NAND2X1 U104 ( .A(n539), .B(n538), .Y(n540) );
  NAND2X1 U105 ( .A(n289), .B(n1260), .Y(n290) );
  NAND2X1 U106 ( .A(n355), .B(n1268), .Y(n356) );
  INVX1 U107 ( .A(n463), .Y(n391) );
  INVX1 U108 ( .A(n1288), .Y(n829) );
  ADDFHX1 U109 ( .A(n1033), .B(n1032), .CI(n1031), .CO(n532), .S(mult_x_1_n586) );
  INVX1 U110 ( .A(n1005), .Y(n28) );
  NAND2XL U111 ( .A(n725), .B(n726), .Y(n49) );
  ADDFHX1 U112 ( .A(n341), .B(n340), .CI(n339), .CO(n331), .S(n342) );
  NAND2X1 U113 ( .A(n1000), .B(n999), .Y(n1001) );
  NAND2X1 U114 ( .A(n851), .B(n850), .Y(n1074) );
  ADDFHX1 U115 ( .A(n303), .B(n302), .CI(n301), .CO(n325), .S(n328) );
  INVX1 U116 ( .A(n1173), .Y(n1014) );
  NOR2X1 U117 ( .A(n1143), .B(n1106), .Y(n1116) );
  NOR2X1 U118 ( .A(n1143), .B(n1086), .Y(n1104) );
  NOR2X1 U119 ( .A(n1143), .B(n203), .Y(n1092) );
  NOR2X1 U120 ( .A(n1143), .B(n187), .Y(n208) );
  NAND2X1 U121 ( .A(n906), .B(n905), .Y(n1188) );
  NAND2XL U122 ( .A(n947), .B(n946), .Y(n23) );
  OAI2BB1XL U123 ( .A0N(n883), .A1N(n8), .B0(n98), .Y(n102) );
  XOR2X1 U124 ( .A(n61), .B(n91), .Y(PRODUCT[35]) );
  XNOR2X1 U125 ( .A(n222), .B(n221), .Y(PRODUCT[34]) );
  XNOR2X1 U126 ( .A(n1186), .B(n1185), .Y(PRODUCT[38]) );
  NOR2BXL U127 ( .AN(n89), .B(n75), .Y(n61) );
  XNOR2X1 U128 ( .A(n1165), .B(n1164), .Y(PRODUCT[36]) );
  XNOR2X1 U129 ( .A(n1172), .B(n1171), .Y(PRODUCT[37]) );
  OAI21XL U130 ( .A0(n1236), .A1(n220), .B0(n219), .Y(n222) );
  XNOR2X1 U131 ( .A(n466), .B(n465), .Y(PRODUCT[25]) );
  XOR2X1 U132 ( .A(B[2]), .B(B[3]), .Y(n95) );
  INVX1 U133 ( .A(n392), .Y(n461) );
  NOR2X1 U134 ( .A(n1225), .B(n1161), .Y(n1198) );
  NAND2X2 U135 ( .A(n16), .B(n14), .Y(n392) );
  XNOR2X1 U136 ( .A(n752), .B(n751), .Y(PRODUCT[16]) );
  XOR2X1 U137 ( .A(n1285), .B(n829), .Y(PRODUCT[14]) );
  NAND2X1 U138 ( .A(n554), .B(n21), .Y(n20) );
  INVX1 U139 ( .A(n467), .Y(n539) );
  INVXL U140 ( .A(n1284), .Y(n17) );
  INVXL U141 ( .A(n1279), .Y(n687) );
  XOR2X1 U142 ( .A(n1289), .B(n1286), .Y(PRODUCT[13]) );
  CLKINVX3 U143 ( .A(n1281), .Y(n12) );
  INVX1 U144 ( .A(n1255), .Y(n1154) );
  XOR2X1 U145 ( .A(n1002), .B(n46), .Y(n1313) );
  XOR2X1 U146 ( .A(n1007), .B(n35), .Y(n1314) );
  AOI2BB1X2 U147 ( .A0N(n1004), .A1N(n1009), .B0(n28), .Y(n27) );
  AND2X2 U148 ( .A(n1006), .B(n1005), .Y(n1007) );
  ADDFHX2 U149 ( .A(n1072), .B(n1071), .CI(n1070), .CO(mult_x_1_n633), .S(n647) );
  NOR2X1 U150 ( .A(n1004), .B(n1008), .Y(n30) );
  NAND2X1 U151 ( .A(n1016), .B(n1014), .Y(n959) );
  INVXL U152 ( .A(n1008), .Y(n37) );
  OAI21XL U153 ( .A0(n725), .A1(n726), .B0(n724), .Y(n50) );
  INVXL U154 ( .A(n1082), .Y(n826) );
  NAND2XL U155 ( .A(n345), .B(n346), .Y(mult_x_1_n198) );
  INVXL U156 ( .A(n1000), .Y(n47) );
  NAND2X1 U157 ( .A(n823), .B(n822), .Y(mult_x_1_n307) );
  ADDFHX2 U158 ( .A(n1024), .B(n1023), .CI(n1022), .CO(mult_x_1_n537), .S(n460) );
  ADDFHX2 U159 ( .A(n1030), .B(n1029), .CI(n1028), .CO(mult_x_1_n569), .S(n533) );
  ADDFHX1 U160 ( .A(n338), .B(n337), .CI(n336), .CO(n343), .S(n345) );
  NOR2X1 U161 ( .A(n823), .B(n822), .Y(mult_x_1_n306) );
  NAND2BX2 U162 ( .AN(n956), .B(n22), .Y(n1016) );
  ADDFHX2 U163 ( .A(n360), .B(n359), .CI(n358), .CO(n346), .S(n383) );
  OR2XL U164 ( .A(n1151), .B(n1150), .Y(n1153) );
  INVXL U165 ( .A(n1052), .Y(n64) );
  ADDFHX2 U166 ( .A(n833), .B(n832), .CI(n831), .CO(n822), .S(n851) );
  INVXL U167 ( .A(n999), .Y(n48) );
  OAI2BB1XL U168 ( .A0N(n602), .A1N(n41), .B0(n39), .Y(n1045) );
  INVXL U169 ( .A(n1064), .Y(n68) );
  NAND2XL U170 ( .A(n40), .B(n603), .Y(n39) );
  ADDFHX1 U171 ( .A(n139), .B(n138), .CI(n137), .CO(n329), .S(n180) );
  ADDFHX2 U172 ( .A(n735), .B(n734), .CI(n733), .CO(n747), .S(n774) );
  NAND2BXL U173 ( .AN(n603), .B(n42), .Y(n41) );
  INVXL U174 ( .A(n42), .Y(n40) );
  OAI2BB1XL U175 ( .A0N(n5), .A1N(n1121), .B0(n1120), .Y(n1125) );
  ADDFHX1 U176 ( .A(n970), .B(n969), .CI(n968), .CO(n980), .S(n988) );
  ADDFHX1 U177 ( .A(n434), .B(n433), .CI(n432), .CO(n422), .S(n451) );
  ADDFHX1 U178 ( .A(n403), .B(n402), .CI(n401), .CO(n378), .S(n421) );
  ADDFHX1 U179 ( .A(n508), .B(n507), .CI(n506), .CO(n496), .S(n524) );
  XNOR2XL U180 ( .A(n1141), .B(A[22]), .Y(n1118) );
  NAND2BXL U181 ( .AN(n947), .B(n25), .Y(n24) );
  AND2XL U182 ( .A(n1222), .B(n1221), .Y(n1324) );
  OR2XL U183 ( .A(n1220), .B(n1219), .Y(n1222) );
  XNOR2X1 U184 ( .A(n357), .B(n356), .Y(PRODUCT[28]) );
  BUFX3 U185 ( .A(n556), .Y(n9) );
  NAND2X1 U186 ( .A(B[1]), .B(n559), .Y(n714) );
  CLKINVX3 U187 ( .A(n349), .Y(n551) );
  AOI21X1 U188 ( .A0(n7), .A1(n554), .B0(n553), .Y(n650) );
  OR2X2 U189 ( .A(n462), .B(n86), .Y(n80) );
  NAND2X2 U190 ( .A(n85), .B(n347), .Y(n86) );
  NAND2X1 U191 ( .A(n535), .B(n83), .Y(n16) );
  NAND2X1 U192 ( .A(n1296), .B(n1297), .Y(n543) );
  INVXL U193 ( .A(n1265), .Y(n344) );
  INVXL U194 ( .A(A[6]), .Y(n60) );
  INVX1 U195 ( .A(n1288), .Y(n10) );
  NOR2X1 U196 ( .A(n1279), .B(n1277), .Y(n554) );
  AOI21X4 U197 ( .A0(n13), .A1(n12), .B0(n11), .Y(n552) );
  OAI21X2 U198 ( .A0(n1281), .A1(n1287), .B0(n1282), .Y(n11) );
  NOR2X2 U199 ( .A(n10), .B(n1283), .Y(n13) );
  OAI22X1 U200 ( .A0(n409), .A1(n440), .B0(n837), .B1(n411), .Y(n446) );
  NAND2X1 U201 ( .A(n749), .B(n748), .Y(mult_x_1_n287) );
  OAI22X1 U202 ( .A0(n1146), .A1(n664), .B0(n698), .B1(n624), .Y(n660) );
  XNOR2X1 U203 ( .A(n911), .B(A[17]), .Y(n429) );
  XNOR2X1 U204 ( .A(n1123), .B(A[11]), .Y(n170) );
  OAI22X1 U205 ( .A0(n409), .A1(n485), .B0(n837), .B1(n440), .Y(n490) );
  XNOR2X1 U206 ( .A(n1141), .B(A[12]), .Y(n96) );
  OAI22X1 U207 ( .A0(n932), .A1(n663), .B0(n930), .B1(n625), .Y(n677) );
  XNOR2X1 U208 ( .A(n1107), .B(A[8]), .Y(n597) );
  OAI22X1 U209 ( .A0(n409), .A1(n155), .B0(n837), .B1(n128), .Y(n160) );
  OAI22X1 U210 ( .A0(n1121), .A1(n145), .B0(n5), .B1(n117), .Y(n133) );
  XNOR2X1 U211 ( .A(n1107), .B(A[9]), .Y(n503) );
  XNOR2X1 U212 ( .A(n911), .B(A[21]), .Y(n107) );
  NOR2X2 U213 ( .A(n348), .B(n1267), .Y(n85) );
  NOR2X2 U214 ( .A(n467), .B(n1271), .Y(n83) );
  NOR2X1 U215 ( .A(n1294), .B(n1295), .Y(n467) );
  NAND2X2 U216 ( .A(n1299), .B(n1298), .Y(n548) );
  NOR2X4 U217 ( .A(n1296), .B(n1297), .Y(n542) );
  XOR2X1 U218 ( .A(n778), .B(n17), .Y(PRODUCT[15]) );
  OAI21X4 U219 ( .A0(n552), .A1(n20), .B0(n18), .Y(n349) );
  AOI21X2 U220 ( .A0(n553), .A1(n21), .B0(n19), .Y(n18) );
  NOR2X1 U221 ( .A(n1273), .B(n1275), .Y(n21) );
  OAI2BB1X1 U222 ( .A0N(n24), .A1N(n945), .B0(n23), .Y(n987) );
  XOR2X1 U223 ( .A(n945), .B(n26), .Y(n948) );
  XOR2X1 U224 ( .A(n947), .B(n946), .Y(n26) );
  NAND2X1 U225 ( .A(n29), .B(n27), .Y(n1002) );
  NAND2X1 U226 ( .A(n991), .B(n992), .Y(n1005) );
  NAND2X1 U227 ( .A(n1003), .B(n30), .Y(n29) );
  NAND2X2 U228 ( .A(n72), .B(n73), .Y(n1003) );
  OAI2BB1X1 U229 ( .A0N(n32), .A1N(n977), .B0(n31), .Y(n984) );
  NAND2X1 U230 ( .A(n978), .B(n979), .Y(n31) );
  NAND2BX1 U231 ( .AN(n978), .B(n33), .Y(n32) );
  INVXL U232 ( .A(n979), .Y(n33) );
  XOR2X1 U233 ( .A(n977), .B(n34), .Y(n986) );
  XOR2X1 U234 ( .A(n978), .B(n979), .Y(n34) );
  NAND2X1 U235 ( .A(n990), .B(n989), .Y(n1009) );
  NOR2X1 U236 ( .A(n992), .B(n991), .Y(n1004) );
  INVX1 U237 ( .A(n1003), .Y(n1011) );
  NAND2X1 U238 ( .A(n36), .B(n1009), .Y(n35) );
  NAND2X1 U239 ( .A(n1003), .B(n37), .Y(n36) );
  OAI22X2 U240 ( .A0(n595), .A1(n9), .B0(n855), .B1(n38), .Y(n1036) );
  OAI22X1 U241 ( .A0(n558), .A1(n855), .B0(n9), .B1(n38), .Y(n594) );
  XNOR2X1 U242 ( .A(n911), .B(A[13]), .Y(n38) );
  INVX1 U243 ( .A(n1002), .Y(n1080) );
  XNOR3X2 U244 ( .A(n603), .B(n42), .C(n602), .Y(n590) );
  AOI2BB2X2 U245 ( .B0(n44), .B1(n43), .A0N(n409), .A1N(n578), .Y(n42) );
  INVX1 U246 ( .A(n837), .Y(n43) );
  INVX1 U247 ( .A(n577), .Y(n44) );
  NOR2X1 U248 ( .A(n906), .B(n905), .Y(n1187) );
  XOR2X1 U249 ( .A(B[4]), .B(B[5]), .Y(n45) );
  AND2X2 U250 ( .A(n55), .B(n1001), .Y(n46) );
  NAND2X1 U251 ( .A(n48), .B(n47), .Y(n55) );
  NAND2X1 U252 ( .A(n50), .B(n49), .Y(n721) );
  XOR2X1 U253 ( .A(n51), .B(n724), .Y(n749) );
  XNOR2X1 U254 ( .A(n725), .B(n52), .Y(n51) );
  INVX1 U255 ( .A(n726), .Y(n52) );
  XOR2X1 U256 ( .A(B[12]), .B(B[13]), .Y(n92) );
  CLKINVX3 U257 ( .A(B[13]), .Y(n717) );
  BUFX3 U258 ( .A(n94), .Y(n919) );
  NOR2XL U259 ( .A(n1225), .B(n1257), .Y(n217) );
  NAND2XL U260 ( .A(n1154), .B(n1156), .Y(n1159) );
  INVXL U261 ( .A(n1251), .Y(n1167) );
  XNOR2XL U262 ( .A(n928), .B(A[24]), .Y(n193) );
  BUFX1 U263 ( .A(A[7]), .Y(n852) );
  XNOR2XL U264 ( .A(n928), .B(A[22]), .Y(n260) );
  XNOR2X1 U265 ( .A(n1123), .B(A[14]), .Y(n126) );
  XNOR2XL U266 ( .A(n911), .B(A[22]), .Y(n125) );
  BUFX3 U267 ( .A(B[7]), .Y(n911) );
  NOR2XL U268 ( .A(n1261), .B(n1259), .Y(n88) );
  NOR2XL U269 ( .A(n1265), .B(n1263), .Y(n312) );
  NOR2XL U270 ( .A(n1159), .B(n1257), .Y(n1224) );
  NOR2XL U271 ( .A(n1223), .B(n1245), .Y(n1228) );
  OAI21XL U272 ( .A0(n1232), .A1(n1161), .B0(n1160), .Y(n1204) );
  INVXL U273 ( .A(n1229), .Y(n1160) );
  INVXL U274 ( .A(n1223), .Y(n1203) );
  XOR2X1 U275 ( .A(B[14]), .B(B[15]), .Y(n62) );
  XNOR2XL U276 ( .A(n928), .B(A[13]), .Y(n509) );
  XNOR2XL U277 ( .A(n911), .B(A[15]), .Y(n505) );
  NAND2X2 U278 ( .A(n74), .B(n556), .Y(n938) );
  XOR2X1 U279 ( .A(B[6]), .B(B[7]), .Y(n74) );
  NAND2XL U280 ( .A(n1224), .B(n1228), .Y(n1231) );
  INVXL U281 ( .A(n1119), .Y(n1120) );
  OAI22XL U282 ( .A0(n8), .A1(n869), .B0(n671), .B1(n859), .Y(n868) );
  OAI22XL U283 ( .A0(n8), .A1(n889), .B0(n671), .B1(n869), .Y(n899) );
  OAI22XL U284 ( .A0(n1146), .A1(n1124), .B0(n106), .B1(n1144), .Y(n1149) );
  NAND2BXL U285 ( .AN(A[0]), .B(n928), .Y(n929) );
  INVXL U286 ( .A(n1256), .Y(n1157) );
  NOR2XL U287 ( .A(n1236), .B(n90), .Y(n75) );
  INVXL U288 ( .A(n1253), .Y(n1156) );
  AOI21XL U289 ( .A0(n392), .A1(n347), .B0(n385), .Y(n71) );
  INVXL U290 ( .A(n1261), .Y(n316) );
  INVXL U291 ( .A(n1252), .Y(n1166) );
  NAND2XL U292 ( .A(n1198), .B(n1167), .Y(n1169) );
  INVXL U293 ( .A(n1249), .Y(n1170) );
  XNOR2XL U294 ( .A(n928), .B(A[1]), .Y(n913) );
  XNOR2XL U295 ( .A(n911), .B(A[3]), .Y(n912) );
  XNOR2XL U296 ( .A(n911), .B(A[4]), .Y(n840) );
  XNOR2XL U297 ( .A(n911), .B(A[10]), .Y(n633) );
  XNOR2XL U298 ( .A(n928), .B(A[8]), .Y(n625) );
  XNOR2XL U299 ( .A(n928), .B(A[5]), .Y(n739) );
  XNOR2XL U300 ( .A(n911), .B(A[6]), .Y(n770) );
  XNOR2XL U301 ( .A(n911), .B(n852), .Y(n759) );
  XNOR2XL U302 ( .A(n911), .B(A[9]), .Y(n674) );
  XNOR2XL U303 ( .A(n911), .B(A[8]), .Y(n713) );
  XNOR2XL U304 ( .A(n928), .B(A[4]), .Y(n788) );
  XNOR2XL U305 ( .A(n928), .B(A[3]), .Y(n807) );
  NAND2BXL U306 ( .AN(A[0]), .B(n802), .Y(n790) );
  XNOR2XL U307 ( .A(n911), .B(A[20]), .Y(n108) );
  XNOR2XL U308 ( .A(n928), .B(A[17]), .Y(n161) );
  XNOR2XL U309 ( .A(n1123), .B(A[3]), .Y(n613) );
  XNOR2XL U310 ( .A(n1141), .B(A[14]), .Y(n247) );
  XNOR2XL U311 ( .A(n911), .B(A[23]), .Y(n257) );
  XNOR2XL U312 ( .A(n928), .B(A[21]), .Y(n261) );
  XNOR2XL U313 ( .A(n928), .B(A[20]), .Y(n115) );
  OAI22XL U314 ( .A0(n921), .A1(n105), .B0(n919), .B1(n124), .Y(n114) );
  NAND2BXL U315 ( .AN(A[0]), .B(n442), .Y(n861) );
  XNOR2X1 U316 ( .A(n442), .B(A[4]), .Y(n918) );
  XNOR2XL U317 ( .A(n911), .B(A[2]), .Y(n936) );
  NAND2BXL U318 ( .AN(A[0]), .B(n911), .Y(n853) );
  XNOR2X1 U319 ( .A(n442), .B(A[3]), .Y(n920) );
  XNOR2XL U320 ( .A(n911), .B(A[1]), .Y(n937) );
  NAND2XL U321 ( .A(n391), .B(n464), .Y(n465) );
  OAI21XL U322 ( .A0(n551), .A1(n462), .B0(n461), .Y(n466) );
  XNOR2X1 U323 ( .A(n318), .B(n317), .Y(PRODUCT[31]) );
  NAND2XL U324 ( .A(n316), .B(n1262), .Y(n317) );
  OAI21XL U325 ( .A0(n1236), .A1(n315), .B0(n314), .Y(n318) );
  XNOR2X1 U326 ( .A(n335), .B(n334), .Y(PRODUCT[30]) );
  NAND2XL U327 ( .A(n333), .B(n1264), .Y(n334) );
  OAI21XL U328 ( .A0(n1236), .A1(n1265), .B0(n1266), .Y(n335) );
  AND2XL U329 ( .A(n246), .B(n1258), .Y(n54) );
  NAND2XL U330 ( .A(n1167), .B(n1252), .Y(n1164) );
  XOR2X1 U331 ( .A(n650), .B(n649), .Y(PRODUCT[19]) );
  NAND2XL U332 ( .A(n648), .B(n1276), .Y(n649) );
  XOR2X1 U333 ( .A(n79), .B(n56), .Y(PRODUCT[20]) );
  AND2XL U334 ( .A(n555), .B(n1274), .Y(n56) );
  OAI21XL U335 ( .A0(n650), .A1(n1275), .B0(n1276), .Y(n79) );
  OAI22XL U336 ( .A0(n409), .A1(n262), .B0(n410), .B1(n228), .Y(n250) );
  OAI22XL U337 ( .A0(n1146), .A1(n258), .B0(n698), .B1(n227), .Y(n251) );
  ADDFX2 U338 ( .A(n255), .B(n254), .CI(n253), .CO(n236), .S(n292) );
  OAI22X1 U339 ( .A0(n932), .A1(n260), .B0(n930), .B1(n225), .Y(n254) );
  OAI22XL U340 ( .A0(n1121), .A1(n264), .B0(n5), .B1(n224), .Y(n255) );
  XNOR2XL U341 ( .A(n1141), .B(A[20]), .Y(n1086) );
  OAI2BB1XL U342 ( .A0N(n9), .A1N(n855), .B0(n186), .Y(n232) );
  INVXL U343 ( .A(n185), .Y(n186) );
  OAI22XL U344 ( .A0(n409), .A1(n192), .B0(n410), .B1(n204), .Y(n209) );
  OAI22XL U345 ( .A0(n1146), .A1(n190), .B0(n106), .B1(n202), .Y(n211) );
  INVXL U346 ( .A(n188), .Y(n189) );
  XNOR2X1 U347 ( .A(n1107), .B(A[14]), .Y(n145) );
  XNOR2X1 U348 ( .A(n1107), .B(A[15]), .Y(n117) );
  XNOR2XL U349 ( .A(n928), .B(A[18]), .Y(n149) );
  XNOR2XL U350 ( .A(n911), .B(A[19]), .Y(n169) );
  XNOR2XL U351 ( .A(n928), .B(A[16]), .Y(n404) );
  OAI22XL U352 ( .A0(n875), .A1(n407), .B0(n164), .B1(n559), .Y(n406) );
  XNOR2XL U353 ( .A(n911), .B(A[18]), .Y(n398) );
  XNOR2XL U354 ( .A(n928), .B(A[15]), .Y(n435) );
  XNOR2XL U355 ( .A(n928), .B(A[14]), .Y(n480) );
  OAI22XL U356 ( .A0(n875), .A1(n483), .B0(n438), .B1(n559), .Y(n482) );
  XNOR2XL U357 ( .A(n1123), .B(A[8]), .Y(n475) );
  XNOR2XL U358 ( .A(n911), .B(A[16]), .Y(n474) );
  XNOR2X1 U359 ( .A(n1123), .B(A[4]), .Y(n574) );
  XNOR2XL U360 ( .A(n911), .B(A[11]), .Y(n616) );
  OAI22XL U361 ( .A0(n875), .A1(n623), .B0(n561), .B1(n1073), .Y(n619) );
  NAND2BXL U362 ( .AN(A[0]), .B(B[16]), .Y(n562) );
  INVXL U363 ( .A(n97), .Y(n98) );
  AOI21XL U364 ( .A0(n1229), .A1(n1228), .B0(n1227), .Y(n1230) );
  INVXL U365 ( .A(n1226), .Y(n1202) );
  NAND2XL U366 ( .A(n1198), .B(n1203), .Y(n1206) );
  INVXL U367 ( .A(n1245), .Y(n1207) );
  NAND2XL U368 ( .A(n1200), .B(n1248), .Y(n1185) );
  OAI22XL U369 ( .A0(n8), .A1(n884), .B0(n883), .B1(n882), .Y(n885) );
  INVXL U370 ( .A(B[3]), .Y(n884) );
  NAND2BXL U371 ( .AN(A[0]), .B(B[3]), .Y(n882) );
  INVXL U372 ( .A(n1127), .Y(n1115) );
  OAI22XL U373 ( .A0(n1146), .A1(n1105), .B0(n106), .B1(n1114), .Y(n1117) );
  OAI22XL U374 ( .A0(n1146), .A1(n1090), .B0(n106), .B1(n1105), .Y(n1110) );
  CMPR32X1 U375 ( .A(n998), .B(n997), .C(n996), .CO(n999), .S(n992) );
  OAI22XL U376 ( .A0(n932), .A1(n607), .B0(n933), .B1(n509), .Y(n522) );
  ADDFX2 U377 ( .A(n606), .B(n605), .CI(n604), .CO(n1051), .S(n1044) );
  OAI22X1 U378 ( .A0(n8), .A1(n579), .B0(n883), .B1(n515), .Y(n605) );
  OAI22XL U379 ( .A0(n409), .A1(n577), .B0(n837), .B1(n514), .Y(n606) );
  ADDFX2 U380 ( .A(n519), .B(n518), .CI(n517), .CO(n528), .S(n1050) );
  OAI22XL U381 ( .A0(n921), .A1(n516), .B0(n919), .B1(n487), .Y(n517) );
  OAI22X1 U382 ( .A0(n8), .A1(n515), .B0(n883), .B1(n486), .Y(n518) );
  OAI22XL U383 ( .A0(n409), .A1(n514), .B0(n837), .B1(n485), .Y(n519) );
  OAI22XL U384 ( .A0(n932), .A1(n608), .B0(n933), .B1(n607), .Y(n1042) );
  OAI22XL U385 ( .A0(n855), .A1(n595), .B0(n9), .B1(n505), .Y(n1037) );
  OAI22X1 U386 ( .A0(n698), .A1(n504), .B0(n1146), .B1(n59), .Y(n1038) );
  OAI22XL U387 ( .A0(n1121), .A1(n597), .B0(n5), .B1(n503), .Y(n1039) );
  AOI21XL U388 ( .A0(n910), .A1(n1177), .B0(n909), .Y(n1012) );
  NOR2XL U389 ( .A(n886), .B(n885), .Y(n1210) );
  NAND2XL U390 ( .A(n886), .B(n885), .Y(n1211) );
  AOI21XL U391 ( .A0(n1216), .A1(n1217), .B0(n879), .Y(n1213) );
  INVXL U392 ( .A(n1215), .Y(n879) );
  INVXL U393 ( .A(n1221), .Y(n1217) );
  NOR2XL U394 ( .A(n1143), .B(n1142), .Y(n1148) );
  XNOR2XL U395 ( .A(n1141), .B(A[24]), .Y(n1142) );
  INVXL U396 ( .A(n1144), .Y(n1145) );
  INVXL U397 ( .A(n1149), .Y(n1139) );
  XNOR2XL U398 ( .A(n1141), .B(A[23]), .Y(n1122) );
  NOR2X1 U399 ( .A(n1053), .B(n1054), .Y(n65) );
  XOR2X1 U400 ( .A(n1052), .B(n1054), .Y(n66) );
  CMPR32X1 U401 ( .A(n525), .B(n524), .C(n523), .CO(n1033), .S(n1053) );
  NAND2XL U402 ( .A(n1065), .B(n1066), .Y(n67) );
  NOR2X1 U403 ( .A(n1065), .B(n1066), .Y(n69) );
  OAI22XL U404 ( .A0(n875), .A1(A[0]), .B0(n874), .B1(n1073), .Y(n1220) );
  NAND2XL U405 ( .A(n876), .B(n875), .Y(n1219) );
  NAND2BXL U406 ( .AN(A[0]), .B(n926), .Y(n876) );
  NAND2XL U407 ( .A(n1220), .B(n1219), .Y(n1221) );
  NAND2XL U408 ( .A(n895), .B(n894), .Y(n1238) );
  INVXL U409 ( .A(n893), .Y(n1239) );
  NOR2XL U410 ( .A(n895), .B(n894), .Y(n893) );
  INVXL U411 ( .A(n1177), .Y(n1190) );
  INVXL U412 ( .A(n1224), .Y(n1161) );
  NAND2XL U413 ( .A(n1197), .B(n1200), .Y(n1223) );
  NOR2XL U414 ( .A(n1251), .B(n1249), .Y(n1197) );
  INVXL U415 ( .A(n1271), .Y(n471) );
  AOI21XL U416 ( .A0(n392), .A1(n391), .B0(n390), .Y(n393) );
  NAND2XL U417 ( .A(n389), .B(n391), .Y(n394) );
  INVXL U418 ( .A(n1269), .Y(n395) );
  AOI21XL U419 ( .A0(n392), .A1(n352), .B0(n351), .Y(n353) );
  INVXL U420 ( .A(n1267), .Y(n355) );
  INVXL U421 ( .A(n313), .Y(n314) );
  INVXL U422 ( .A(n312), .Y(n315) );
  INVXL U423 ( .A(n1263), .Y(n333) );
  INVXL U424 ( .A(n1257), .Y(n246) );
  INVXL U425 ( .A(n1262), .Y(n286) );
  NAND2XL U426 ( .A(n312), .B(n316), .Y(n288) );
  INVXL U427 ( .A(n1259), .Y(n289) );
  INVXL U428 ( .A(n1204), .Y(n1162) );
  INVXL U429 ( .A(n1198), .Y(n1163) );
  INVXL U430 ( .A(n1280), .Y(n686) );
  INVXL U431 ( .A(n1273), .Y(n555) );
  NAND2X1 U432 ( .A(n1295), .B(n1294), .Y(n538) );
  NOR2X2 U433 ( .A(n1298), .B(n1299), .Y(n547) );
  XNOR2XL U434 ( .A(n911), .B(A[25]), .Y(n185) );
  ADDFX2 U435 ( .A(n662), .B(n661), .CI(n660), .CO(n669), .S(n704) );
  OAI22X1 U436 ( .A0(n875), .A1(n657), .B0(n623), .B1(n1073), .Y(n661) );
  NOR2BXL U437 ( .AN(A[0]), .B(n182), .Y(n662) );
  XNOR2XL U438 ( .A(n928), .B(n852), .Y(n663) );
  XNOR2XL U439 ( .A(n928), .B(A[6]), .Y(n706) );
  NAND2BXL U440 ( .AN(A[0]), .B(n1123), .Y(n658) );
  OAI22X1 U441 ( .A0(n932), .A1(n931), .B0(n930), .B1(n929), .Y(n963) );
  INVXL U442 ( .A(n928), .Y(n931) );
  XNOR2XL U443 ( .A(n928), .B(A[2]), .Y(n839) );
  XNOR2XL U444 ( .A(n802), .B(A[20]), .Y(n262) );
  AOI21XL U445 ( .A0(n1157), .A1(n1156), .B0(n1155), .Y(n1158) );
  INVXL U446 ( .A(n1254), .Y(n1155) );
  AOI21XL U447 ( .A0(n1201), .A1(n1200), .B0(n1199), .Y(n1226) );
  INVXL U448 ( .A(n1248), .Y(n1199) );
  INVX1 U449 ( .A(n349), .Y(n81) );
  NAND2XL U450 ( .A(n1198), .B(n1197), .Y(n1184) );
  INVXL U451 ( .A(n1247), .Y(n1200) );
  NAND2XL U452 ( .A(n1154), .B(n1256), .Y(n221) );
  NAND2XL U453 ( .A(n1156), .B(n1254), .Y(n91) );
  OAI21XL U454 ( .A0(n829), .A1(n1242), .B0(n1243), .Y(n778) );
  XNOR2X1 U455 ( .A(n397), .B(n396), .Y(PRODUCT[26]) );
  NAND2XL U456 ( .A(n395), .B(n1270), .Y(n396) );
  OAI21XL U457 ( .A0(n551), .A1(n394), .B0(n393), .Y(n397) );
  XOR2X1 U458 ( .A(n70), .B(n53), .Y(PRODUCT[27]) );
  AND2XL U459 ( .A(n388), .B(n387), .Y(n53) );
  OAI21XL U460 ( .A0(n386), .A1(n551), .B0(n71), .Y(n70) );
  NAND2XL U461 ( .A(n1170), .B(n1250), .Y(n1171) );
  XOR2X1 U462 ( .A(n723), .B(n552), .Y(PRODUCT[17]) );
  NAND2XL U463 ( .A(n687), .B(n1280), .Y(n723) );
  OAI22XL U464 ( .A0(n8), .A1(n924), .B0(n671), .B1(n842), .Y(n974) );
  OAI22X1 U465 ( .A0(n936), .A1(n938), .B0(n912), .B1(n9), .Y(n970) );
  OAI22XL U466 ( .A0(n916), .A1(n918), .B0(n919), .B1(n915), .Y(n968) );
  OAI22X1 U467 ( .A0(n932), .A1(n914), .B0(n930), .B1(n913), .Y(n969) );
  OAI22XL U468 ( .A0(n875), .A1(n768), .B0(n715), .B1(n1073), .Y(n767) );
  NAND2BXL U469 ( .AN(A[0]), .B(n1107), .Y(n716) );
  ADDFX2 U470 ( .A(n845), .B(n844), .CI(n843), .CO(n848), .S(n971) );
  OAI22XL U471 ( .A0(n8), .A1(n842), .B0(n671), .B1(n805), .Y(n843) );
  CMPR32X1 U472 ( .A(n812), .B(n811), .C(n810), .CO(n798), .S(n846) );
  OAI22XL U473 ( .A0(n938), .A1(n801), .B0(n9), .B1(n770), .Y(n812) );
  OAI22X1 U474 ( .A0(n8), .A1(n805), .B0(n883), .B1(n771), .Y(n811) );
  OAI22XL U475 ( .A0(n916), .A1(n772), .B0(n919), .B1(n741), .Y(n785) );
  OAI22X1 U476 ( .A0(n932), .A1(n788), .B0(n930), .B1(n739), .Y(n787) );
  OAI22XL U477 ( .A0(n8), .A1(n771), .B0(n883), .B1(n740), .Y(n786) );
  OAI22XL U478 ( .A0(n932), .A1(n225), .B0(n930), .B1(n193), .Y(n231) );
  OAI22XL U479 ( .A0(n1121), .A1(n224), .B0(n5), .B1(n195), .Y(n229) );
  OAI22XL U480 ( .A0(n1146), .A1(n227), .B0(n106), .B1(n194), .Y(n230) );
  INVXL U481 ( .A(n207), .Y(n196) );
  OAI22XL U482 ( .A0(n1121), .A1(n627), .B0(n5), .B1(n615), .Y(n634) );
  OAI22XL U483 ( .A0(n938), .A1(n633), .B0(n9), .B1(n616), .Y(n639) );
  ADDFX2 U484 ( .A(n669), .B(n668), .CI(n667), .CO(n683), .S(n719) );
  OAI22XL U485 ( .A0(n938), .A1(n674), .B0(n9), .B1(n633), .Y(n678) );
  OAI22XL U486 ( .A0(n409), .A1(n673), .B0(n837), .B1(n632), .Y(n679) );
  OAI22XL U487 ( .A0(n921), .A1(n697), .B0(n919), .B1(n631), .Y(n680) );
  ADDFX2 U488 ( .A(n677), .B(n676), .CI(n675), .CO(n668), .S(n728) );
  OAI22X1 U489 ( .A0(n8), .A1(n672), .B0(n883), .B1(n626), .Y(n676) );
  OAI22XL U490 ( .A0(n1121), .A1(n666), .B0(n5), .B1(n627), .Y(n675) );
  CMPR32X1 U491 ( .A(n705), .B(n704), .C(n703), .CO(n720), .S(n746) );
  ADDFX2 U492 ( .A(n744), .B(n743), .CI(n742), .CO(n758), .S(n779) );
  OAI22XL U493 ( .A0(n8), .A1(n740), .B0(n671), .B1(n708), .Y(n742) );
  OAI22XL U494 ( .A0(n409), .A1(n762), .B0(n837), .B1(n707), .Y(n743) );
  OAI22XL U495 ( .A0(n932), .A1(n739), .B0(n930), .B1(n706), .Y(n744) );
  OAI22XL U496 ( .A0(n938), .A1(n770), .B0(n9), .B1(n759), .Y(n784) );
  OAI22XL U497 ( .A0(n409), .A1(n769), .B0(n837), .B1(n762), .Y(n782) );
  CMPR32X1 U498 ( .A(n765), .B(n764), .C(n763), .CO(n756), .S(n796) );
  OAI22XL U499 ( .A0(n938), .A1(n759), .B0(n9), .B1(n713), .Y(n764) );
  OAI22XL U500 ( .A0(n921), .A1(n741), .B0(n919), .B1(n712), .Y(n765) );
  OAI22XL U501 ( .A0(n938), .A1(n713), .B0(n9), .B1(n674), .Y(n730) );
  OAI22XL U502 ( .A0(n8), .A1(n708), .B0(n883), .B1(n672), .Y(n732) );
  ADDFX2 U503 ( .A(n962), .B(n961), .CI(n960), .CO(n847), .S(n998) );
  OAI22X1 U504 ( .A0(n932), .A1(n839), .B0(n930), .B1(n807), .Y(n961) );
  OAI22XL U505 ( .A0(n921), .A1(n841), .B0(n919), .B1(n806), .Y(n962) );
  OAI22XL U506 ( .A0(n932), .A1(n807), .B0(n933), .B1(n788), .Y(n836) );
  INVXL U507 ( .A(n151), .Y(n130) );
  CMPR32X1 U508 ( .A(n148), .B(n147), .C(n146), .CO(n139), .S(n167) );
  OAI22XL U509 ( .A0(n855), .A1(n108), .B0(n9), .B1(n107), .Y(n148) );
  OAI22XL U510 ( .A0(n575), .A1(n111), .B0(n698), .B1(n110), .Y(n146) );
  NOR2XL U511 ( .A(n182), .B(n109), .Y(n147) );
  OAI22XL U512 ( .A0(n932), .A1(n161), .B0(n930), .B1(n149), .Y(n178) );
  ADDFX2 U513 ( .A(n369), .B(n368), .CI(n367), .CO(n375), .S(n424) );
  OAI22X1 U514 ( .A0(n8), .A1(n365), .B0(n883), .B1(n156), .Y(n368) );
  OAI22XL U515 ( .A0(n409), .A1(n364), .B0(n837), .B1(n155), .Y(n369) );
  OAI22XL U516 ( .A0(n409), .A1(n411), .B0(n837), .B1(n364), .Y(n416) );
  OAI22XL U517 ( .A0(n8), .A1(n412), .B0(n883), .B1(n365), .Y(n415) );
  XNOR2XL U518 ( .A(n802), .B(A[12]), .Y(n440) );
  ADDFX2 U519 ( .A(n446), .B(n445), .CI(n444), .CO(n455), .S(n498) );
  OAI22XL U520 ( .A0(n921), .A1(n443), .B0(n919), .B1(n413), .Y(n444) );
  OAI22X1 U521 ( .A0(n8), .A1(n441), .B0(n883), .B1(n412), .Y(n445) );
  XNOR2XL U522 ( .A(n802), .B(A[10]), .Y(n514) );
  XNOR2XL U523 ( .A(n802), .B(A[11]), .Y(n485) );
  XNOR2XL U524 ( .A(n928), .B(A[12]), .Y(n607) );
  OAI22XL U525 ( .A0(n875), .A1(n584), .B0(n512), .B1(n559), .Y(n610) );
  XNOR2XL U526 ( .A(n928), .B(A[11]), .Y(n608) );
  XOR2X1 U527 ( .A(n1123), .B(n60), .Y(n59) );
  XNOR2XL U528 ( .A(n911), .B(A[14]), .Y(n595) );
  ADDFX2 U529 ( .A(n630), .B(n629), .CI(n628), .CO(n642), .S(n667) );
  OAI22XL U530 ( .A0(n921), .A1(n631), .B0(n919), .B1(n563), .Y(n628) );
  OAI22XL U531 ( .A0(n409), .A1(n632), .B0(n837), .B1(n573), .Y(n630) );
  OAI22X1 U532 ( .A0(n8), .A1(n626), .B0(n883), .B1(n576), .Y(n629) );
  OAI22XL U533 ( .A0(n8), .A1(n576), .B0(n883), .B1(n580), .Y(n620) );
  OAI22XL U534 ( .A0(n409), .A1(n573), .B0(n837), .B1(n578), .Y(n622) );
  OAI2BB1XL U535 ( .A0N(n919), .A1N(n921), .B0(n249), .Y(n272) );
  INVXL U536 ( .A(n248), .Y(n249) );
  OAI22XL U537 ( .A0(n932), .A1(n261), .B0(n930), .B1(n260), .Y(n275) );
  OAI22XL U538 ( .A0(n1146), .A1(n259), .B0(n106), .B1(n258), .Y(n276) );
  OAI22XL U539 ( .A0(n409), .A1(n127), .B0(n410), .B1(n263), .Y(n269) );
  OAI22XL U540 ( .A0(n932), .A1(n115), .B0(n930), .B1(n261), .Y(n300) );
  INVXL U541 ( .A(n442), .Y(n862) );
  NOR2BXL U542 ( .AN(A[0]), .B(n933), .Y(n941) );
  INVXL U543 ( .A(n911), .Y(n854) );
  OAI22XL U544 ( .A0(n921), .A1(n858), .B0(n919), .B1(n920), .Y(n942) );
  OAI22X1 U545 ( .A0(n8), .A1(n859), .B0(n883), .B1(n917), .Y(n944) );
  OAI22XL U546 ( .A0(n409), .A1(n228), .B0(n410), .B1(n223), .Y(n237) );
  OAI22XL U547 ( .A0(n875), .A1(n874), .B0(n880), .B1(n1073), .Y(n878) );
  NOR2BXL U548 ( .AN(A[0]), .B(n671), .Y(n877) );
  INVXL U549 ( .A(n1087), .Y(n1088) );
  INVXL U550 ( .A(n1103), .Y(n1091) );
  OAI22XL U551 ( .A0(n1146), .A1(n202), .B0(n106), .B1(n1090), .Y(n1093) );
  OAI22XL U552 ( .A0(n1121), .A1(n205), .B0(n5), .B1(n1089), .Y(n1096) );
  ADDFX2 U553 ( .A(n160), .B(n159), .CI(n158), .CO(n363), .S(n374) );
  OAI2BB1XL U554 ( .A0N(n1073), .A1N(n875), .B0(n130), .Y(n158) );
  OAI22XL U555 ( .A0(n8), .A1(n156), .B0(n883), .B1(n129), .Y(n159) );
  INVXL U556 ( .A(n103), .Y(n131) );
  OAI22XL U557 ( .A0(n932), .A1(n149), .B0(n930), .B1(n116), .Y(n136) );
  OR2XL U558 ( .A(n154), .B(n153), .Y(n134) );
  OAI22XL U559 ( .A0(n1121), .A1(n400), .B0(n5), .B1(n172), .Y(n401) );
  OAI22XL U560 ( .A0(n932), .A1(n435), .B0(n930), .B1(n404), .Y(n419) );
  ADDFX2 U561 ( .A(n375), .B(n374), .CI(n373), .CO(n381), .S(n427) );
  ADDFX2 U562 ( .A(n378), .B(n377), .CI(n376), .CO(n379), .S(n426) );
  OAI22XL U563 ( .A0(n1121), .A1(n431), .B0(n5), .B1(n400), .Y(n432) );
  OAI22XL U564 ( .A0(n932), .A1(n480), .B0(n930), .B1(n435), .Y(n449) );
  OAI22XL U565 ( .A0(n1121), .A1(n476), .B0(n5), .B1(n431), .Y(n477) );
  OAI22XL U566 ( .A0(n932), .A1(n509), .B0(n930), .B1(n480), .Y(n493) );
  ADDFX2 U567 ( .A(n490), .B(n489), .CI(n488), .CO(n499), .S(n527) );
  OAI22XL U568 ( .A0(n921), .A1(n487), .B0(n919), .B1(n443), .Y(n488) );
  OAI22X1 U569 ( .A0(n8), .A1(n486), .B0(n883), .B1(n441), .Y(n489) );
  ADDFX2 U570 ( .A(n499), .B(n498), .CI(n497), .CO(n502), .S(n529) );
  OAI22XL U571 ( .A0(n1121), .A1(n503), .B0(n5), .B1(n476), .Y(n506) );
  OAI22XL U572 ( .A0(n1121), .A1(n557), .B0(n5), .B1(n598), .Y(n592) );
  OAI22XL U573 ( .A0(n938), .A1(n616), .B0(n9), .B1(n558), .Y(n569) );
  ADDFX2 U574 ( .A(n566), .B(n565), .CI(n564), .CO(n572), .S(n641) );
  OAI22X1 U575 ( .A0(n921), .A1(n563), .B0(n919), .B1(n582), .Y(n565) );
  OAI22XL U576 ( .A0(n932), .A1(n617), .B0(n930), .B1(n583), .Y(n566) );
  OAI22XL U577 ( .A0(n1121), .A1(n615), .B0(n5), .B1(n557), .Y(n564) );
  OAI22XL U578 ( .A0(n714), .A1(n888), .B0(n887), .B1(n1073), .Y(n901) );
  NOR2BXL U579 ( .AN(A[0]), .B(n919), .Y(n902) );
  OAI22XL U580 ( .A0(n8), .A1(n890), .B0(n883), .B1(n889), .Y(n900) );
  INVXL U581 ( .A(n1233), .Y(n1234) );
  OR2XL U582 ( .A(n1225), .B(n1231), .Y(n1235) );
  NAND2XL U583 ( .A(n1207), .B(n1246), .Y(n1208) );
  AOI21XL U584 ( .A0(n1240), .A1(n1239), .B0(n896), .Y(n1195) );
  INVXL U585 ( .A(n1238), .Y(n896) );
  NAND2XL U586 ( .A(n878), .B(n877), .Y(n1215) );
  OAI22XL U587 ( .A0(n1146), .A1(n1114), .B0(n106), .B1(n1124), .Y(n1133) );
  INVXL U588 ( .A(mult_x_1_n306), .Y(n830) );
  NAND2XL U589 ( .A(n1016), .B(n1015), .Y(n1017) );
  NOR2XL U590 ( .A(n332), .B(n331), .Y(mult_x_1_n183) );
  NOR2XL U591 ( .A(n1098), .B(n1097), .Y(mult_x_1_n136) );
  NAND2XL U592 ( .A(n1180), .B(n1179), .Y(n1181) );
  INVXL U593 ( .A(n1178), .Y(n1180) );
  XOR2XL U594 ( .A(n1196), .B(n1195), .Y(n1320) );
  NAND2XL U595 ( .A(n1194), .B(n1193), .Y(n1196) );
  INVXL U596 ( .A(n1192), .Y(n1194) );
  NAND2XL U597 ( .A(n1212), .B(n1211), .Y(n1214) );
  INVXL U598 ( .A(n1210), .Y(n1212) );
  XNOR2XL U599 ( .A(n1218), .B(n1217), .Y(n1323) );
  NAND2XL U600 ( .A(n1216), .B(n1215), .Y(n1218) );
  NOR2X1 U601 ( .A(n346), .B(n345), .Y(mult_x_1_n197) );
  NAND2XL U602 ( .A(n1153), .B(n1152), .Y(mult_x_1_n58) );
  NAND2XL U603 ( .A(n1151), .B(n1150), .Y(n1152) );
  NOR2XL U604 ( .A(n1135), .B(n1134), .Y(mult_x_1_n109) );
  NAND2XL U605 ( .A(n1135), .B(n1134), .Y(mult_x_1_n110) );
  NOR2XL U606 ( .A(n1137), .B(n1136), .Y(mult_x_1_n120) );
  NAND2XL U607 ( .A(n1137), .B(n1136), .Y(mult_x_1_n121) );
  NOR2XL U608 ( .A(n1113), .B(n1112), .Y(mult_x_1_n129) );
  NAND2XL U609 ( .A(n1113), .B(n1112), .Y(mult_x_1_n130) );
  NAND2XL U610 ( .A(n1098), .B(n1097), .Y(mult_x_1_n137) );
  NAND2XL U611 ( .A(n828), .B(n1082), .Y(mult_x_1_n83) );
  AOI21XL U612 ( .A0(n828), .A1(n827), .B0(n826), .Y(mult_x_1_n296) );
  INVXL U613 ( .A(mult_x_1_n307), .Y(n827) );
  OAI21X1 U614 ( .A0(n65), .A1(n64), .B0(n63), .Y(n1032) );
  NAND2X1 U615 ( .A(n1053), .B(n1054), .Y(n63) );
  OAI21X1 U616 ( .A0(n69), .A1(n68), .B0(n67), .Y(n1056) );
  XOR2X1 U617 ( .A(n1053), .B(n66), .Y(n1055) );
  NOR2BXL U618 ( .AN(A[0]), .B(n1073), .Y(n1325) );
  NAND2XL U619 ( .A(n1239), .B(n1238), .Y(n1241) );
  NAND2XL U620 ( .A(n1189), .B(n1188), .Y(n1191) );
  INVXL U621 ( .A(n1187), .Y(n1189) );
  NAND2XL U622 ( .A(n1014), .B(n1174), .Y(n1175) );
  INVX1 U623 ( .A(B[1]), .Y(n150) );
  BUFX8 U624 ( .A(n106), .Y(n698) );
  AND2X1 U625 ( .A(n344), .B(n1266), .Y(n57) );
  XOR2X1 U626 ( .A(n76), .B(n54), .Y(PRODUCT[33]) );
  NOR2X1 U627 ( .A(n825), .B(n824), .Y(n1081) );
  XNOR2X1 U628 ( .A(n1236), .B(n57), .Y(PRODUCT[29]) );
  OAI21XL U629 ( .A0(n1236), .A1(n288), .B0(n287), .Y(n291) );
  OAI21XL U630 ( .A0(n1236), .A1(n1225), .B0(n1232), .Y(n76) );
  OAI22X1 U631 ( .A0(n855), .A1(n256), .B0(n9), .B1(n185), .Y(n233) );
  CMPR22X1 U632 ( .A(n437), .B(n436), .CO(n417), .S(n448) );
  CMPR22X1 U633 ( .A(n511), .B(n510), .CO(n491), .S(n521) );
  CMPR22X1 U634 ( .A(n588), .B(n587), .CO(n599), .S(n568) );
  CMPR22X1 U635 ( .A(n612), .B(n611), .CO(n1040), .S(n600) );
  ADDFX2 U636 ( .A(n175), .B(n174), .CI(n173), .CO(n168), .S(n377) );
  CMPR22X1 U637 ( .A(n873), .B(n872), .CO(n867), .S(n897) );
  CMPR22X1 U638 ( .A(n163), .B(n162), .CO(n177), .S(n371) );
  OAI22X1 U639 ( .A0(n875), .A1(n934), .B0(n927), .B1(n1073), .Y(n964) );
  OAI22X1 U640 ( .A0(n916), .A1(n712), .B0(n919), .B1(n697), .Y(n735) );
  OAI22X1 U641 ( .A0(n855), .A1(n854), .B0(n9), .B1(n853), .Y(n922) );
  CMPR22X1 U642 ( .A(n809), .B(n808), .CO(n835), .S(n960) );
  OAI22X1 U643 ( .A0(n409), .A1(n791), .B0(n837), .B1(n790), .Y(n808) );
  OAI22X1 U644 ( .A0(n932), .A1(n193), .B0(n930), .B1(n188), .Y(n207) );
  OAI22X2 U645 ( .A0(n8), .A1(n129), .B0(n883), .B1(n97), .Y(n103) );
  CMPR22X1 U646 ( .A(n702), .B(n701), .CO(n705), .S(n733) );
  NAND2X1 U647 ( .A(n544), .B(n543), .Y(n545) );
  NOR2X1 U648 ( .A(n182), .B(n123), .Y(n267) );
  OAI22X1 U649 ( .A0(n1146), .A1(n504), .B0(n698), .B1(n475), .Y(n507) );
  NOR2X1 U650 ( .A(n908), .B(n907), .Y(n1178) );
  OAI22X4 U651 ( .A0(n596), .A1(n1146), .B0(n698), .B1(n59), .Y(n1035) );
  XNOR2X4 U652 ( .A(B[14]), .B(B[13]), .Y(n106) );
  XOR3X2 U653 ( .A(n1064), .B(n1066), .C(n1065), .Y(n1067) );
  AOI21X1 U654 ( .A0(n7), .A1(n687), .B0(n686), .Y(n690) );
  OAI21XL U655 ( .A0(n551), .A1(n470), .B0(n469), .Y(n473) );
  XNOR2X1 U656 ( .A(n473), .B(n472), .Y(PRODUCT[24]) );
  NOR2X1 U657 ( .A(n990), .B(n989), .Y(n1008) );
  AOI21X1 U658 ( .A0(n1016), .A1(n1013), .B0(n958), .Y(n72) );
  OR2X2 U659 ( .A(n959), .B(n1012), .Y(n73) );
  NOR2X4 U660 ( .A(n78), .B(n77), .Y(n1236) );
  OAI21X2 U661 ( .A0(n461), .A1(n86), .B0(n82), .Y(n77) );
  NOR2X1 U662 ( .A(n81), .B(n80), .Y(n78) );
  OAI22X2 U663 ( .A0(n1146), .A1(n430), .B0(n698), .B1(n399), .Y(n433) );
  OAI22X2 U664 ( .A0(n1146), .A1(n475), .B0(n698), .B1(n430), .Y(n478) );
  OAI22X2 U665 ( .A0(n1146), .A1(n399), .B0(n698), .B1(n170), .Y(n402) );
  OAI22X2 U666 ( .A0(n1146), .A1(n574), .B0(n698), .B1(n596), .Y(n593) );
  OAI22X1 U667 ( .A0(n575), .A1(n613), .B0(n698), .B1(n574), .Y(n621) );
  OAI22X1 U668 ( .A0(n1146), .A1(n665), .B0(n698), .B1(n664), .Y(n710) );
  AOI21X1 U669 ( .A0(n313), .A1(n88), .B0(n87), .Y(n1232) );
  OAI21XL U670 ( .A0(n1263), .A1(n1266), .B0(n1264), .Y(n313) );
  XNOR2X2 U671 ( .A(B[16]), .B(B[15]), .Y(n182) );
  NAND2X1 U672 ( .A(n92), .B(n171), .Y(n93) );
  OAI22X1 U673 ( .A0(n409), .A1(n804), .B0(n837), .B1(n803), .Y(n844) );
  NOR2BX1 U674 ( .AN(A[0]), .B(n837), .Y(n967) );
  OAI22X1 U675 ( .A0(n855), .A1(n505), .B0(n9), .B1(n474), .Y(n508) );
  OAI22X1 U676 ( .A0(n855), .A1(n429), .B0(n9), .B1(n398), .Y(n434) );
  OAI22X1 U677 ( .A0(n855), .A1(n474), .B0(n9), .B1(n429), .Y(n479) );
  INVX8 U678 ( .A(n717), .Y(n1107) );
  XNOR2XL U679 ( .A(n928), .B(A[23]), .Y(n225) );
  XNOR2XL U680 ( .A(B[3]), .B(A[12]), .Y(n708) );
  XNOR2X1 U681 ( .A(n1107), .B(A[17]), .Y(n265) );
  OAI22X1 U682 ( .A0(n1121), .A1(n122), .B0(n5), .B1(n265), .Y(n268) );
  XNOR2XL U683 ( .A(B[3]), .B(A[3]), .Y(n869) );
  XNOR2XL U684 ( .A(n1141), .B(A[19]), .Y(n203) );
  XNOR2XL U685 ( .A(n928), .B(A[19]), .Y(n116) );
  OAI22X1 U686 ( .A0(n855), .A1(n398), .B0(n9), .B1(n169), .Y(n403) );
  XOR2XL U687 ( .A(n1214), .B(n1213), .Y(n1322) );
  NAND2X1 U688 ( .A(n1292), .B(n1293), .Y(n464) );
  OAI21XL U689 ( .A0(n1269), .A1(n464), .B0(n1270), .Y(n385) );
  NAND2XL U690 ( .A(n1290), .B(n1291), .Y(n387) );
  OAI21XL U691 ( .A0(n1267), .A1(n387), .B0(n1268), .Y(n84) );
  NAND2XL U692 ( .A(n312), .B(n88), .Y(n1225) );
  NAND2XL U693 ( .A(n217), .B(n1154), .Y(n90) );
  OAI21XL U694 ( .A0(n1259), .A1(n1262), .B0(n1260), .Y(n87) );
  OAI21XL U695 ( .A0(n1232), .A1(n1257), .B0(n1258), .Y(n218) );
  AOI21XL U696 ( .A0(n218), .A1(n1154), .B0(n1157), .Y(n89) );
  XNOR2X1 U697 ( .A(B[12]), .B(B[11]), .Y(n171) );
  BUFX3 U698 ( .A(B[5]), .Y(n442) );
  XNOR2X1 U699 ( .A(n442), .B(A[22]), .Y(n143) );
  OAI22XL U700 ( .A0(n921), .A1(n143), .B0(n919), .B1(n105), .Y(n132) );
  XNOR2X1 U701 ( .A(B[2]), .B(B[1]), .Y(n671) );
  NAND2X1 U702 ( .A(n95), .B(n671), .Y(n670) );
  XNOR2X1 U703 ( .A(B[3]), .B(A[24]), .Y(n129) );
  BUFX3 U704 ( .A(n671), .Y(n883) );
  XNOR2X1 U705 ( .A(B[3]), .B(A[25]), .Y(n97) );
  NOR2XL U706 ( .A(n182), .B(n96), .Y(n104) );
  XOR2X1 U707 ( .A(B[8]), .B(B[9]), .Y(n99) );
  XNOR2X1 U708 ( .A(B[8]), .B(B[7]), .Y(n933) );
  NAND2X1 U709 ( .A(n99), .B(n933), .Y(n100) );
  XOR2X1 U710 ( .A(B[10]), .B(B[11]), .Y(n101) );
  XNOR2X2 U711 ( .A(B[10]), .B(B[9]), .Y(n410) );
  INVX4 U712 ( .A(B[11]), .Y(n791) );
  XNOR2X1 U713 ( .A(n802), .B(A[16]), .Y(n128) );
  XNOR2XL U714 ( .A(n802), .B(A[17]), .Y(n118) );
  OAI22XL U715 ( .A0(n409), .A1(n128), .B0(n837), .B1(n118), .Y(n135) );
  OAI22XL U716 ( .A0(n855), .A1(n169), .B0(n9), .B1(n108), .Y(n154) );
  BUFX12 U717 ( .A(n575), .Y(n1146) );
  INVX4 U718 ( .A(B[15]), .Y(n659) );
  INVX8 U719 ( .A(n659), .Y(n1123) );
  XNOR2X1 U720 ( .A(n1123), .B(A[12]), .Y(n111) );
  OAI22X1 U721 ( .A0(n1146), .A1(n170), .B0(n698), .B1(n111), .Y(n153) );
  ADDFHX1 U722 ( .A(n104), .B(n103), .CI(n102), .CO(n299), .S(n141) );
  XNOR2X1 U723 ( .A(n442), .B(A[24]), .Y(n124) );
  XNOR2X1 U724 ( .A(n1123), .B(A[13]), .Y(n110) );
  OAI22X1 U725 ( .A0(n1146), .A1(n110), .B0(n698), .B1(n126), .Y(n113) );
  OAI22XL U726 ( .A0(n855), .A1(n107), .B0(n9), .B1(n125), .Y(n112) );
  XNOR2XL U727 ( .A(B[16]), .B(A[11]), .Y(n109) );
  OAI22XL U728 ( .A0(n932), .A1(n116), .B0(n930), .B1(n115), .Y(n121) );
  XNOR2X1 U729 ( .A(n1107), .B(A[16]), .Y(n122) );
  OAI22X1 U730 ( .A0(n1121), .A1(n117), .B0(n5), .B1(n122), .Y(n120) );
  XNOR2XL U731 ( .A(n802), .B(A[18]), .Y(n127) );
  OAI22XL U732 ( .A0(n409), .A1(n118), .B0(n410), .B1(n127), .Y(n119) );
  XNOR2XL U733 ( .A(n1141), .B(A[13]), .Y(n123) );
  OAI22X1 U734 ( .A0(n921), .A1(n124), .B0(n919), .B1(n248), .Y(n273) );
  INVXL U735 ( .A(n273), .Y(n266) );
  OAI22XL U736 ( .A0(n855), .A1(n125), .B0(n9), .B1(n257), .Y(n271) );
  XNOR2X1 U737 ( .A(n1123), .B(A[15]), .Y(n259) );
  OAI22X1 U738 ( .A0(n1146), .A1(n126), .B0(n106), .B1(n259), .Y(n270) );
  XNOR2X1 U739 ( .A(n802), .B(A[19]), .Y(n263) );
  XNOR2X1 U740 ( .A(n802), .B(A[15]), .Y(n155) );
  XNOR2X1 U741 ( .A(B[3]), .B(A[23]), .Y(n156) );
  INVX1 U742 ( .A(B[0]), .Y(n559) );
  BUFX3 U743 ( .A(n559), .Y(n1073) );
  BUFX3 U744 ( .A(n714), .Y(n875) );
  CLKINVX3 U745 ( .A(n150), .Y(n926) );
  XNOR2X1 U746 ( .A(n926), .B(A[25]), .Y(n151) );
  CMPR32X1 U747 ( .A(n133), .B(n132), .C(n131), .CO(n142), .S(n362) );
  CMPR32X1 U748 ( .A(n136), .B(n135), .C(n134), .CO(n140), .S(n361) );
  CMPR32X1 U749 ( .A(n142), .B(n141), .C(n140), .CO(n338), .S(n179) );
  XNOR2XL U750 ( .A(n442), .B(A[21]), .Y(n157) );
  OAI22X1 U751 ( .A0(n921), .A1(n157), .B0(n919), .B1(n143), .Y(n175) );
  XNOR2X1 U752 ( .A(B[16]), .B(A[10]), .Y(n144) );
  NOR2XL U753 ( .A(n182), .B(n144), .Y(n174) );
  XNOR2X1 U754 ( .A(n1107), .B(A[13]), .Y(n172) );
  OAI22XL U755 ( .A0(n1121), .A1(n172), .B0(n5), .B1(n145), .Y(n173) );
  XNOR2X1 U756 ( .A(B[1]), .B(A[24]), .Y(n164) );
  OAI22X1 U757 ( .A0(n875), .A1(n164), .B0(n151), .B1(n1073), .Y(n163) );
  XNOR2XL U758 ( .A(B[16]), .B(A[9]), .Y(n152) );
  NOR2XL U759 ( .A(n182), .B(n152), .Y(n162) );
  XNOR2X1 U760 ( .A(n154), .B(n153), .Y(n176) );
  INVX8 U761 ( .A(n791), .Y(n802) );
  XNOR2X1 U762 ( .A(n802), .B(A[14]), .Y(n364) );
  XNOR2X1 U763 ( .A(B[3]), .B(A[22]), .Y(n365) );
  XNOR2XL U764 ( .A(n442), .B(A[20]), .Y(n366) );
  OAI22XL U765 ( .A0(n921), .A1(n366), .B0(n919), .B1(n157), .Y(n367) );
  OAI22XL U766 ( .A0(n932), .A1(n404), .B0(n930), .B1(n161), .Y(n372) );
  XNOR2X1 U767 ( .A(B[1]), .B(A[23]), .Y(n407) );
  XNOR2XL U768 ( .A(B[16]), .B(A[8]), .Y(n165) );
  NOR2XL U769 ( .A(n182), .B(n165), .Y(n405) );
  CMPR32X1 U770 ( .A(n168), .B(n167), .C(n166), .CO(n360), .S(n380) );
  XNOR2X1 U771 ( .A(n1123), .B(A[10]), .Y(n399) );
  XNOR2X1 U772 ( .A(n1107), .B(A[12]), .Y(n400) );
  CMPR32X1 U773 ( .A(n178), .B(n177), .C(n176), .CO(n166), .S(n376) );
  ADDFHX1 U774 ( .A(n181), .B(n180), .CI(n179), .CO(n336), .S(n358) );
  XNOR2X1 U775 ( .A(n1107), .B(A[20]), .Y(n195) );
  XNOR2X1 U776 ( .A(n1107), .B(A[21]), .Y(n191) );
  OAI22XL U777 ( .A0(n1121), .A1(n195), .B0(n5), .B1(n191), .Y(n201) );
  BUFX3 U778 ( .A(n182), .Y(n1143) );
  XNOR2X1 U779 ( .A(n1141), .B(A[17]), .Y(n183) );
  XNOR2XL U780 ( .A(n911), .B(A[24]), .Y(n256) );
  XNOR2X1 U781 ( .A(n1123), .B(A[18]), .Y(n194) );
  XNOR2X1 U782 ( .A(n1123), .B(A[19]), .Y(n190) );
  OAI22XL U783 ( .A0(n1146), .A1(n194), .B0(n106), .B1(n190), .Y(n198) );
  XNOR2XL U784 ( .A(n802), .B(A[23]), .Y(n192) );
  OAI22XL U785 ( .A0(n409), .A1(n223), .B0(n410), .B1(n192), .Y(n197) );
  XNOR2XL U786 ( .A(n928), .B(A[25]), .Y(n188) );
  XNOR2X1 U787 ( .A(n1141), .B(A[18]), .Y(n187) );
  OAI2BB1X1 U788 ( .A0N(n930), .A1N(n932), .B0(n189), .Y(n206) );
  XNOR2XL U789 ( .A(n1107), .B(A[22]), .Y(n205) );
  OAI22XL U790 ( .A0(n1121), .A1(n191), .B0(n5), .B1(n205), .Y(n210) );
  XNOR2X1 U791 ( .A(n802), .B(A[24]), .Y(n204) );
  XNOR2X1 U792 ( .A(n1123), .B(A[17]), .Y(n227) );
  XNOR2X1 U793 ( .A(n1107), .B(A[19]), .Y(n224) );
  CMPR32X1 U794 ( .A(n198), .B(n197), .C(n196), .CO(n214), .S(n239) );
  CMPR32X1 U795 ( .A(n201), .B(n200), .C(n199), .CO(n243), .S(n238) );
  XNOR2X1 U796 ( .A(n1123), .B(A[21]), .Y(n1090) );
  XNOR2X1 U797 ( .A(n802), .B(A[25]), .Y(n1087) );
  OAI22X1 U798 ( .A0(n409), .A1(n204), .B0(n410), .B1(n1087), .Y(n1103) );
  XNOR2X1 U799 ( .A(n1107), .B(A[23]), .Y(n1089) );
  CMPR32X1 U800 ( .A(n208), .B(n207), .C(n206), .CO(n1095), .S(n213) );
  CMPR32X1 U801 ( .A(n211), .B(n210), .C(n209), .CO(n1094), .S(n212) );
  CMPR32X1 U802 ( .A(n214), .B(n213), .C(n212), .CO(n1083), .S(n242) );
  NOR2XL U803 ( .A(n216), .B(n215), .Y(mult_x_1_n151) );
  NAND2XL U804 ( .A(n216), .B(n215), .Y(mult_x_1_n152) );
  INVXL U805 ( .A(n217), .Y(n220) );
  INVXL U806 ( .A(n218), .Y(n219) );
  XNOR2X1 U807 ( .A(n802), .B(A[21]), .Y(n228) );
  XNOR2X1 U808 ( .A(n1107), .B(A[18]), .Y(n264) );
  INVXL U809 ( .A(n233), .Y(n253) );
  XNOR2X1 U810 ( .A(n1141), .B(A[15]), .Y(n226) );
  XNOR2X1 U811 ( .A(n1123), .B(A[16]), .Y(n258) );
  CMPR32X1 U812 ( .A(n231), .B(n230), .C(n229), .CO(n240), .S(n280) );
  CMPR32X1 U813 ( .A(n234), .B(n233), .C(n232), .CO(n199), .S(n279) );
  ADDFHX1 U814 ( .A(n237), .B(n236), .CI(n235), .CO(n283), .S(n278) );
  CMPR32X1 U815 ( .A(n240), .B(n239), .C(n238), .CO(n241), .S(n281) );
  CMPR32X1 U816 ( .A(n243), .B(n242), .C(n241), .CO(n216), .S(n244) );
  NOR2XL U817 ( .A(n245), .B(n244), .Y(mult_x_1_n160) );
  NAND2XL U818 ( .A(n245), .B(n244), .Y(mult_x_1_n161) );
  CMPR32X1 U819 ( .A(n252), .B(n251), .C(n250), .CO(n235), .S(n293) );
  OAI22XL U820 ( .A0(n855), .A1(n257), .B0(n9), .B1(n256), .Y(n277) );
  OAI22X1 U821 ( .A0(n409), .A1(n263), .B0(n837), .B1(n262), .Y(n297) );
  CMPR32X1 U822 ( .A(n274), .B(n273), .C(n272), .CO(n294), .S(n323) );
  CMPR32X1 U823 ( .A(n277), .B(n276), .C(n275), .CO(n306), .S(n322) );
  CMPR32X1 U824 ( .A(n283), .B(n282), .C(n281), .CO(n245), .S(n284) );
  NOR2XL U825 ( .A(n285), .B(n284), .Y(mult_x_1_n169) );
  NAND2XL U826 ( .A(n285), .B(n284), .Y(mult_x_1_n170) );
  AOI21XL U827 ( .A0(n313), .A1(n316), .B0(n286), .Y(n287) );
  XNOR2X1 U828 ( .A(n291), .B(n290), .Y(PRODUCT[32]) );
  CMPR32X1 U829 ( .A(n294), .B(n293), .C(n292), .CO(n309), .S(n321) );
  CMPR32X1 U830 ( .A(n300), .B(n299), .C(n298), .CO(n326), .S(n330) );
  CMPR32X1 U831 ( .A(n306), .B(n305), .C(n304), .CO(n308), .S(n319) );
  ADDFHX1 U832 ( .A(n309), .B(n308), .CI(n307), .CO(n285), .S(n310) );
  NOR2XL U833 ( .A(n311), .B(n310), .Y(mult_x_1_n176) );
  NAND2XL U834 ( .A(n311), .B(n310), .Y(mult_x_1_n177) );
  ADDFHX1 U835 ( .A(n321), .B(n320), .CI(n319), .CO(n311), .S(n332) );
  ADDFHX1 U836 ( .A(n330), .B(n329), .CI(n328), .CO(n339), .S(n337) );
  NAND2XL U837 ( .A(n332), .B(n331), .Y(mult_x_1_n184) );
  NOR2XL U838 ( .A(n343), .B(n342), .Y(mult_x_1_n194) );
  NAND2XL U839 ( .A(n343), .B(n342), .Y(mult_x_1_n195) );
  INVXL U840 ( .A(n347), .Y(n384) );
  INVXL U841 ( .A(n348), .Y(n388) );
  NOR2XL U842 ( .A(n384), .B(n348), .Y(n352) );
  INVX1 U843 ( .A(n462), .Y(n389) );
  NAND2XL U844 ( .A(n352), .B(n389), .Y(n354) );
  INVXL U845 ( .A(n385), .Y(n350) );
  OAI21XL U846 ( .A0(n350), .A1(n348), .B0(n387), .Y(n351) );
  OAI21XL U847 ( .A0(n354), .A1(n551), .B0(n353), .Y(n357) );
  ADDFHX1 U848 ( .A(n363), .B(n362), .CI(n361), .CO(n181), .S(n1021) );
  XNOR2X1 U849 ( .A(n802), .B(A[13]), .Y(n411) );
  XNOR2X1 U850 ( .A(B[3]), .B(A[21]), .Y(n412) );
  XNOR2X1 U851 ( .A(n442), .B(A[19]), .Y(n413) );
  OAI22XL U852 ( .A0(n921), .A1(n413), .B0(n919), .B1(n366), .Y(n414) );
  CMPR32X1 U853 ( .A(n372), .B(n371), .C(n370), .CO(n373), .S(n423) );
  ADDFHX4 U854 ( .A(n381), .B(n380), .CI(n379), .CO(n359), .S(n1019) );
  NOR2X1 U855 ( .A(n383), .B(n382), .Y(mult_x_1_n206) );
  NAND2XL U856 ( .A(n383), .B(n382), .Y(mult_x_1_n207) );
  NAND2XL U857 ( .A(n389), .B(n347), .Y(n386) );
  INVXL U858 ( .A(n464), .Y(n390) );
  XNOR2X1 U859 ( .A(n1107), .B(A[11]), .Y(n431) );
  ADDHXL U860 ( .A(n406), .B(n405), .CO(n370), .S(n418) );
  OAI22X1 U861 ( .A0(n875), .A1(n438), .B0(n407), .B1(n1073), .Y(n437) );
  XNOR2XL U862 ( .A(B[16]), .B(n852), .Y(n408) );
  NOR2XL U863 ( .A(n182), .B(n408), .Y(n436) );
  XNOR2X1 U864 ( .A(B[3]), .B(A[20]), .Y(n441) );
  XNOR2X1 U865 ( .A(n442), .B(A[18]), .Y(n443) );
  CMPR32X1 U866 ( .A(n416), .B(n415), .C(n414), .CO(n425), .S(n454) );
  CMPR32X1 U867 ( .A(n419), .B(n417), .C(n418), .CO(n420), .S(n453) );
  CMPR32X1 U868 ( .A(n422), .B(n421), .C(n420), .CO(n1024), .S(n457) );
  CMPR32X1 U869 ( .A(n425), .B(n424), .C(n423), .CO(n428), .S(n456) );
  XNOR2X1 U870 ( .A(n1107), .B(A[10]), .Y(n476) );
  XNOR2X1 U871 ( .A(B[1]), .B(A[21]), .Y(n483) );
  XNOR2XL U872 ( .A(B[16]), .B(A[6]), .Y(n439) );
  NOR2XL U873 ( .A(n182), .B(n439), .Y(n481) );
  XNOR2X1 U874 ( .A(B[3]), .B(A[19]), .Y(n486) );
  XNOR2X1 U875 ( .A(n442), .B(A[17]), .Y(n487) );
  CMPR32X1 U876 ( .A(n449), .B(n448), .C(n447), .CO(n450), .S(n497) );
  ADDFX2 U877 ( .A(n452), .B(n451), .CI(n450), .CO(n1027), .S(n501) );
  NOR2X1 U878 ( .A(n460), .B(n459), .Y(mult_x_1_n226) );
  NAND2XL U879 ( .A(n460), .B(n459), .Y(mult_x_1_n227) );
  NAND2XL U880 ( .A(n534), .B(n539), .Y(n470) );
  INVXL U881 ( .A(n538), .Y(n468) );
  AOI21XL U882 ( .A0(n535), .A1(n539), .B0(n468), .Y(n469) );
  NAND2X1 U883 ( .A(n471), .B(n1272), .Y(n472) );
  XNOR2X1 U884 ( .A(n1123), .B(n852), .Y(n504) );
  ADDHXL U885 ( .A(n482), .B(n481), .CO(n447), .S(n492) );
  XNOR2X1 U886 ( .A(B[1]), .B(A[20]), .Y(n512) );
  OAI22X1 U887 ( .A0(n875), .A1(n512), .B0(n483), .B1(n1073), .Y(n511) );
  XNOR2X1 U888 ( .A(B[16]), .B(A[5]), .Y(n484) );
  NOR2XL U889 ( .A(n182), .B(n484), .Y(n510) );
  XNOR2X1 U890 ( .A(B[3]), .B(A[18]), .Y(n515) );
  XNOR2XL U891 ( .A(n442), .B(A[16]), .Y(n516) );
  CMPR32X1 U892 ( .A(n493), .B(n491), .C(n492), .CO(n494), .S(n526) );
  XNOR2XL U893 ( .A(B[16]), .B(A[4]), .Y(n513) );
  NOR2XL U894 ( .A(n182), .B(n513), .Y(n609) );
  XNOR2X1 U895 ( .A(n802), .B(A[9]), .Y(n577) );
  XNOR2X1 U896 ( .A(B[3]), .B(A[17]), .Y(n579) );
  XNOR2XL U897 ( .A(n442), .B(A[15]), .Y(n581) );
  OAI22XL U898 ( .A0(n921), .A1(n581), .B0(n919), .B1(n516), .Y(n604) );
  CMPR32X1 U899 ( .A(n522), .B(n521), .C(n520), .CO(n523), .S(n1049) );
  ADDFHX4 U900 ( .A(n531), .B(n530), .CI(n529), .CO(n1029), .S(n1031) );
  NOR2X1 U901 ( .A(n533), .B(n532), .Y(mult_x_1_n244) );
  NAND2XL U902 ( .A(n533), .B(n532), .Y(mult_x_1_n245) );
  INVXL U903 ( .A(n534), .Y(n537) );
  INVXL U904 ( .A(n535), .Y(n536) );
  OAI21XL U905 ( .A0(n551), .A1(n537), .B0(n536), .Y(n541) );
  XNOR2X1 U906 ( .A(n541), .B(n540), .Y(PRODUCT[23]) );
  OAI21XL U907 ( .A0(n551), .A1(n547), .B0(n548), .Y(n546) );
  INVXL U908 ( .A(n542), .Y(n544) );
  XNOR2X1 U909 ( .A(n546), .B(n545), .Y(PRODUCT[22]) );
  INVXL U910 ( .A(n547), .Y(n549) );
  NAND2X1 U911 ( .A(n549), .B(n548), .Y(n550) );
  XOR2X1 U912 ( .A(n551), .B(n550), .Y(PRODUCT[21]) );
  XNOR2XL U913 ( .A(n928), .B(A[9]), .Y(n617) );
  XNOR2XL U914 ( .A(n928), .B(A[10]), .Y(n583) );
  XNOR2X1 U915 ( .A(n442), .B(A[13]), .Y(n563) );
  XNOR2X1 U916 ( .A(n442), .B(A[14]), .Y(n582) );
  XNOR2X1 U917 ( .A(n1107), .B(A[6]), .Y(n557) );
  XNOR2XL U918 ( .A(n911), .B(A[12]), .Y(n558) );
  XNOR2X1 U919 ( .A(n1123), .B(A[5]), .Y(n596) );
  XNOR2X1 U920 ( .A(n1107), .B(n852), .Y(n598) );
  XNOR2X1 U921 ( .A(B[1]), .B(A[17]), .Y(n561) );
  XNOR2X1 U922 ( .A(n926), .B(A[18]), .Y(n585) );
  OAI22X1 U923 ( .A0(n875), .A1(n561), .B0(n585), .B1(n559), .Y(n588) );
  XNOR2XL U924 ( .A(B[16]), .B(A[2]), .Y(n560) );
  NOR2XL U925 ( .A(n182), .B(n560), .Y(n587) );
  XNOR2X1 U926 ( .A(B[1]), .B(A[16]), .Y(n623) );
  XNOR2X1 U927 ( .A(n802), .B(A[6]), .Y(n632) );
  XNOR2X1 U928 ( .A(n802), .B(n852), .Y(n573) );
  XNOR2X1 U929 ( .A(B[3]), .B(A[14]), .Y(n626) );
  XNOR2X1 U930 ( .A(B[3]), .B(A[15]), .Y(n576) );
  XNOR2X1 U931 ( .A(n442), .B(A[12]), .Y(n631) );
  CMPR32X1 U932 ( .A(n569), .B(n568), .C(n567), .CO(n570), .S(n640) );
  XNOR2X1 U933 ( .A(B[3]), .B(A[16]), .Y(n580) );
  OAI22X1 U934 ( .A0(n8), .A1(n580), .B0(n883), .B1(n579), .Y(n603) );
  OAI22XL U935 ( .A0(n921), .A1(n582), .B0(n919), .B1(n581), .Y(n602) );
  OAI22XL U936 ( .A0(n932), .A1(n583), .B0(n930), .B1(n608), .Y(n601) );
  OAI22X1 U937 ( .A0(n875), .A1(n585), .B0(n584), .B1(n1073), .Y(n612) );
  XNOR2XL U938 ( .A(B[16]), .B(A[3]), .Y(n586) );
  NOR2XL U939 ( .A(n182), .B(n586), .Y(n611) );
  CMPR32X1 U940 ( .A(n591), .B(n590), .C(n589), .CO(n1063), .S(n643) );
  OAI22X1 U941 ( .A0(n1121), .A1(n598), .B0(n5), .B1(n597), .Y(n1034) );
  CMPR32X1 U942 ( .A(n601), .B(n600), .C(n599), .CO(n1058), .S(n589) );
  ADDHXL U943 ( .A(n610), .B(n609), .CO(n520), .S(n1041) );
  XNOR2X1 U944 ( .A(n1123), .B(A[2]), .Y(n624) );
  OAI22X1 U945 ( .A0(n1146), .A1(n624), .B0(n698), .B1(n613), .Y(n636) );
  XNOR2X1 U946 ( .A(B[16]), .B(A[1]), .Y(n614) );
  NOR2X1 U947 ( .A(n1143), .B(n614), .Y(n635) );
  XNOR2X1 U948 ( .A(n1107), .B(A[4]), .Y(n627) );
  OAI22XL U949 ( .A0(n932), .A1(n625), .B0(n930), .B1(n617), .Y(n638) );
  ADDHXL U950 ( .A(n619), .B(n618), .CO(n567), .S(n637) );
  ADDFHX1 U951 ( .A(n622), .B(n621), .CI(n620), .CO(n591), .S(n654) );
  XNOR2X1 U952 ( .A(B[1]), .B(A[15]), .Y(n657) );
  XNOR2X1 U953 ( .A(B[3]), .B(A[13]), .Y(n672) );
  XNOR2X1 U954 ( .A(n442), .B(A[11]), .Y(n697) );
  XNOR2X1 U955 ( .A(n802), .B(A[5]), .Y(n673) );
  ADDFX2 U956 ( .A(n636), .B(n635), .CI(n634), .CO(n656), .S(n695) );
  CMPR32X1 U957 ( .A(n639), .B(n638), .C(n637), .CO(n655), .S(n694) );
  ADDFHX4 U958 ( .A(n645), .B(n644), .CI(n643), .CO(n1071), .S(n651) );
  NOR2X1 U959 ( .A(n647), .B(n646), .Y(mult_x_1_n273) );
  NAND2X1 U960 ( .A(n647), .B(n646), .Y(mult_x_1_n274) );
  INVXL U961 ( .A(n1275), .Y(n648) );
  CMPR32X1 U962 ( .A(n656), .B(n655), .C(n654), .CO(n653), .S(n693) );
  XNOR2X1 U963 ( .A(n926), .B(A[14]), .Y(n699) );
  OAI22X1 U964 ( .A0(n875), .A1(n699), .B0(n657), .B1(n1073), .Y(n702) );
  OAI22X1 U965 ( .A0(n1146), .A1(n659), .B0(n698), .B1(n658), .Y(n701) );
  OAI22XL U966 ( .A0(n932), .A1(n706), .B0(n930), .B1(n663), .Y(n711) );
  XNOR2X1 U967 ( .A(n1123), .B(A[0]), .Y(n665) );
  XNOR2X1 U968 ( .A(n1107), .B(A[2]), .Y(n700) );
  OAI22XL U969 ( .A0(n1121), .A1(n700), .B0(n5), .B1(n666), .Y(n709) );
  XNOR2X1 U970 ( .A(n802), .B(A[4]), .Y(n707) );
  OAI22XL U971 ( .A0(n409), .A1(n707), .B0(n837), .B1(n673), .Y(n731) );
  CMPR32X1 U972 ( .A(n680), .B(n679), .C(n678), .CO(n696), .S(n727) );
  NOR2XL U973 ( .A(n685), .B(n684), .Y(mult_x_1_n276) );
  INVXL U974 ( .A(n1277), .Y(n688) );
  NAND2X1 U975 ( .A(n688), .B(n1278), .Y(n689) );
  XOR2X1 U976 ( .A(n690), .B(n689), .Y(PRODUCT[18]) );
  XNOR2X1 U977 ( .A(n442), .B(A[10]), .Y(n712) );
  OAI22X2 U978 ( .A0(n875), .A1(n715), .B0(n699), .B1(n1073), .Y(n737) );
  XNOR2X1 U979 ( .A(n1107), .B(A[1]), .Y(n760) );
  OAI22X1 U980 ( .A0(n1121), .A1(n760), .B0(n5), .B1(n700), .Y(n736) );
  XNOR2X1 U981 ( .A(n802), .B(A[3]), .Y(n762) );
  XNOR2X1 U982 ( .A(B[3]), .B(A[11]), .Y(n740) );
  ADDFHX1 U983 ( .A(n711), .B(n710), .CI(n709), .CO(n703), .S(n757) );
  XNOR2X1 U984 ( .A(n442), .B(A[9]), .Y(n741) );
  XNOR2X1 U985 ( .A(n926), .B(A[12]), .Y(n768) );
  OAI22XL U986 ( .A0(n1121), .A1(n717), .B0(n5), .B1(n716), .Y(n766) );
  NOR2XL U987 ( .A(n722), .B(n721), .Y(mult_x_1_n281) );
  NAND2XL U988 ( .A(n722), .B(n721), .Y(mult_x_1_n282) );
  CMPR32X1 U989 ( .A(n729), .B(n728), .C(n727), .CO(n718), .S(n755) );
  CMPR32X1 U990 ( .A(n732), .B(n731), .C(n730), .CO(n729), .S(n775) );
  ADDFHX4 U991 ( .A(n738), .B(n737), .CI(n736), .CO(n734), .S(n781) );
  XNOR2X1 U992 ( .A(B[3]), .B(A[10]), .Y(n771) );
  XNOR2XL U993 ( .A(n442), .B(A[8]), .Y(n772) );
  ADDFHX1 U994 ( .A(n747), .B(n746), .CI(n745), .CO(n725), .S(n753) );
  NOR2XL U995 ( .A(n749), .B(n748), .Y(mult_x_1_n286) );
  OAI21XL U996 ( .A0(n829), .A1(n1283), .B0(n1287), .Y(n752) );
  INVXL U997 ( .A(n1281), .Y(n750) );
  NAND2XL U998 ( .A(n750), .B(n1282), .Y(n751) );
  CMPR32X1 U999 ( .A(n755), .B(n754), .C(n753), .CO(n748), .S(n777) );
  CMPR32X1 U1000 ( .A(n758), .B(n757), .C(n756), .CO(n745), .S(n818) );
  XNOR2X1 U1001 ( .A(n1107), .B(A[0]), .Y(n761) );
  OAI22X1 U1002 ( .A0(n1121), .A1(n761), .B0(n5), .B1(n760), .Y(n783) );
  XNOR2X1 U1003 ( .A(n802), .B(A[2]), .Y(n769) );
  ADDHXL U1004 ( .A(n767), .B(n766), .CO(n763), .S(n800) );
  NOR2BX1 U1005 ( .AN(A[0]), .B(n5), .Y(n794) );
  XNOR2X1 U1006 ( .A(n926), .B(A[11]), .Y(n789) );
  OAI22X1 U1007 ( .A0(n875), .A1(n789), .B0(n768), .B1(n1073), .Y(n793) );
  XNOR2X1 U1008 ( .A(n802), .B(A[1]), .Y(n803) );
  OAI22XL U1009 ( .A0(n409), .A1(n803), .B0(n837), .B1(n769), .Y(n792) );
  XNOR2XL U1010 ( .A(n911), .B(A[5]), .Y(n801) );
  XNOR2X1 U1011 ( .A(B[3]), .B(A[9]), .Y(n805) );
  XNOR2X1 U1012 ( .A(n442), .B(n852), .Y(n806) );
  OAI22XL U1013 ( .A0(n921), .A1(n806), .B0(n919), .B1(n772), .Y(n810) );
  CMPR32X1 U1014 ( .A(n775), .B(n774), .C(n773), .CO(n754), .S(n816) );
  NOR2XL U1015 ( .A(n777), .B(n776), .Y(mult_x_1_n292) );
  NAND2XL U1016 ( .A(n777), .B(n776), .Y(mult_x_1_n293) );
  CMPR32X1 U1017 ( .A(n784), .B(n783), .C(n782), .CO(n797), .S(n815) );
  CMPR32X1 U1018 ( .A(n787), .B(n786), .C(n785), .CO(n780), .S(n814) );
  OAI22X1 U1019 ( .A0(n875), .A1(n838), .B0(n789), .B1(n1073), .Y(n809) );
  CMPR32X1 U1020 ( .A(n794), .B(n793), .C(n792), .CO(n799), .S(n834) );
  ADDFHX1 U1021 ( .A(n800), .B(n799), .CI(n798), .CO(n795), .S(n833) );
  OAI22XL U1022 ( .A0(n938), .A1(n840), .B0(n9), .B1(n801), .Y(n845) );
  XNOR2X1 U1023 ( .A(n802), .B(A[0]), .Y(n804) );
  XNOR2X1 U1024 ( .A(B[3]), .B(A[8]), .Y(n842) );
  INVX1 U1025 ( .A(n1081), .Y(n828) );
  NAND2XL U1026 ( .A(n828), .B(n830), .Y(mult_x_1_n295) );
  NAND2X1 U1027 ( .A(n825), .B(n824), .Y(n1082) );
  NAND2XL U1028 ( .A(n830), .B(mult_x_1_n307), .Y(mult_x_1_n84) );
  CMPR32X1 U1029 ( .A(n836), .B(n835), .C(n834), .CO(n813), .S(n995) );
  XNOR2X1 U1030 ( .A(n926), .B(A[9]), .Y(n927) );
  OAI22X2 U1031 ( .A0(n875), .A1(n927), .B0(n838), .B1(n1073), .Y(n966) );
  OAI22X1 U1032 ( .A0(n932), .A1(n913), .B0(n930), .B1(n839), .Y(n965) );
  OAI22X1 U1033 ( .A0(n938), .A1(n912), .B0(n9), .B1(n840), .Y(n976) );
  XNOR2X1 U1034 ( .A(n442), .B(A[5]), .Y(n915) );
  OAI22X2 U1035 ( .A0(n921), .A1(n915), .B0(n919), .B1(n841), .Y(n975) );
  XNOR2X1 U1036 ( .A(B[3]), .B(n852), .Y(n924) );
  NOR2X1 U1037 ( .A(n851), .B(n850), .Y(n849) );
  INVX1 U1038 ( .A(n849), .Y(n1077) );
  NAND2XL U1039 ( .A(n1077), .B(n1074), .Y(mult_x_1_n85) );
  XNOR2X1 U1040 ( .A(n926), .B(A[6]), .Y(n856) );
  XNOR2XL U1041 ( .A(n926), .B(n852), .Y(n935) );
  OAI22X1 U1042 ( .A0(n714), .A1(n856), .B0(n935), .B1(n1073), .Y(n923) );
  NOR2BX1 U1043 ( .AN(A[0]), .B(n9), .Y(n865) );
  XNOR2X1 U1044 ( .A(n926), .B(A[5]), .Y(n860) );
  OAI22X1 U1045 ( .A0(n875), .A1(n860), .B0(n856), .B1(n1073), .Y(n864) );
  XNOR2X1 U1046 ( .A(n442), .B(A[1]), .Y(n870) );
  XNOR2X1 U1047 ( .A(n442), .B(A[2]), .Y(n858) );
  OAI22X1 U1048 ( .A0(n921), .A1(n870), .B0(n919), .B1(n858), .Y(n863) );
  XNOR2X1 U1049 ( .A(B[3]), .B(A[4]), .Y(n859) );
  XNOR2X1 U1050 ( .A(B[3]), .B(A[5]), .Y(n917) );
  XNOR2XL U1051 ( .A(n911), .B(A[0]), .Y(n857) );
  OAI22X2 U1052 ( .A0(n938), .A1(n857), .B0(n9), .B1(n937), .Y(n943) );
  XNOR2X1 U1053 ( .A(n926), .B(A[4]), .Y(n887) );
  OAI22X1 U1054 ( .A0(n875), .A1(n887), .B0(n860), .B1(n1073), .Y(n873) );
  OAI22X1 U1055 ( .A0(n921), .A1(n862), .B0(n919), .B1(n861), .Y(n872) );
  CMPR32X1 U1056 ( .A(n865), .B(n864), .C(n863), .CO(n952), .S(n866) );
  CMPR32X1 U1057 ( .A(n868), .B(n867), .C(n866), .CO(n907), .S(n906) );
  XNOR2X1 U1058 ( .A(B[3]), .B(A[2]), .Y(n889) );
  XNOR2XL U1059 ( .A(n442), .B(A[0]), .Y(n871) );
  OAI22XL U1060 ( .A0(n916), .A1(n871), .B0(n919), .B1(n870), .Y(n898) );
  NOR2XL U1061 ( .A(n1178), .B(n1187), .Y(n910) );
  XNOR2X1 U1062 ( .A(n926), .B(A[1]), .Y(n874) );
  XNOR2X1 U1063 ( .A(n926), .B(A[2]), .Y(n880) );
  OR2X2 U1064 ( .A(n878), .B(n877), .Y(n1216) );
  XNOR2X1 U1065 ( .A(n926), .B(A[3]), .Y(n888) );
  OAI22X1 U1066 ( .A0(n875), .A1(n880), .B0(n888), .B1(n1073), .Y(n892) );
  XNOR2X1 U1067 ( .A(B[3]), .B(A[1]), .Y(n890) );
  OAI22X1 U1068 ( .A0(n8), .A1(n881), .B0(n883), .B1(n890), .Y(n891) );
  OAI21XL U1069 ( .A0(n1213), .A1(n1210), .B0(n1211), .Y(n1240) );
  CMPR22X1 U1070 ( .A(n892), .B(n891), .CO(n894), .S(n886) );
  CMPR32X1 U1071 ( .A(n899), .B(n898), .C(n897), .CO(n905), .S(n904) );
  CMPR32X1 U1072 ( .A(n902), .B(n901), .C(n900), .CO(n903), .S(n895) );
  NOR2XL U1073 ( .A(n904), .B(n903), .Y(n1192) );
  NAND2XL U1074 ( .A(n904), .B(n903), .Y(n1193) );
  OAI21XL U1075 ( .A0(n1195), .A1(n1192), .B0(n1193), .Y(n1177) );
  NAND2XL U1076 ( .A(n908), .B(n907), .Y(n1179) );
  OAI21XL U1077 ( .A0(n1178), .A1(n1188), .B0(n1179), .Y(n909) );
  XNOR2XL U1078 ( .A(n928), .B(A[0]), .Y(n914) );
  XNOR2X1 U1079 ( .A(B[3]), .B(A[6]), .Y(n925) );
  OAI22X1 U1080 ( .A0(n8), .A1(n917), .B0(n671), .B1(n925), .Y(n947) );
  OAI22X1 U1081 ( .A0(n921), .A1(n920), .B0(n919), .B1(n918), .Y(n946) );
  OAI22X1 U1082 ( .A0(n8), .A1(n925), .B0(n883), .B1(n924), .Y(n979) );
  XNOR2XL U1083 ( .A(n926), .B(A[8]), .Y(n934) );
  OAI22XL U1084 ( .A0(n714), .A1(n935), .B0(n934), .B1(n1073), .Y(n940) );
  OAI22XL U1085 ( .A0(n938), .A1(n937), .B0(n9), .B1(n936), .Y(n939) );
  CMPR32X1 U1086 ( .A(n941), .B(n940), .C(n939), .CO(n977), .S(n950) );
  ADDFHX1 U1087 ( .A(n953), .B(n952), .CI(n951), .CO(n954), .S(n908) );
  NOR2XL U1088 ( .A(n955), .B(n954), .Y(n1173) );
  NAND2XL U1089 ( .A(n955), .B(n954), .Y(n1174) );
  INVXL U1090 ( .A(n1174), .Y(n1013) );
  NAND2XL U1091 ( .A(n957), .B(n956), .Y(n1015) );
  INVXL U1092 ( .A(n1015), .Y(n958) );
  CMPR22X1 U1093 ( .A(n964), .B(n963), .CO(n982), .S(n978) );
  ADDFHX4 U1094 ( .A(n967), .B(n966), .CI(n965), .CO(n973), .S(n981) );
  CMPR32X1 U1095 ( .A(n985), .B(n984), .C(n983), .CO(n991), .S(n990) );
  CMPR32X1 U1096 ( .A(n988), .B(n987), .C(n986), .CO(n989), .S(n956) );
  AOI21XL U1097 ( .A0(n1002), .A1(n55), .B0(n1076), .Y(mult_x_1_n316) );
  INVXL U1098 ( .A(n1004), .Y(n1006) );
  NAND2XL U1099 ( .A(n37), .B(n1009), .Y(n1010) );
  INVXL U1100 ( .A(n1012), .Y(n1176) );
  AOI21XL U1101 ( .A0(n1176), .A1(n1014), .B0(n1013), .Y(n1018) );
  ADDFHX1 U1102 ( .A(n1039), .B(n1038), .CI(n1037), .CO(n525), .S(n1047) );
  CMPR32X1 U1103 ( .A(n1042), .B(n1040), .C(n1041), .CO(n1046), .S(n1043) );
  CMPR32X1 U1104 ( .A(n1045), .B(n1044), .C(n1043), .CO(n1066), .S(n1061) );
  CMPR32X1 U1105 ( .A(n1048), .B(n1047), .C(n1046), .CO(n1057), .S(n1065) );
  ADDFHX1 U1106 ( .A(n1057), .B(n1056), .CI(n1055), .CO(mult_x_1_n601), .S(
        mult_x_1_n602) );
  CMPR32X1 U1107 ( .A(n1060), .B(n1059), .C(n1058), .CO(n1069), .S(n1062) );
  CMPR32X1 U1108 ( .A(n1063), .B(n1062), .C(n1061), .CO(n1068), .S(n1070) );
  ADDFHX1 U1109 ( .A(n1069), .B(n1068), .CI(n1067), .CO(mult_x_1_n617), .S(
        mult_x_1_n618) );
  NAND2XL U1110 ( .A(n1077), .B(n55), .Y(n1079) );
  INVXL U1111 ( .A(n1074), .Y(n1075) );
  AOI21XL U1112 ( .A0(n1077), .A1(n1076), .B0(n1075), .Y(n1078) );
  OAI21XL U1113 ( .A0(n1080), .A1(n1079), .B0(n1078), .Y(mult_x_1_n309) );
  CMPR32X1 U1114 ( .A(n1085), .B(n1084), .C(n1083), .CO(n1098), .S(n215) );
  OAI2BB1X1 U1115 ( .A0N(n410), .A1N(n409), .B0(n1088), .Y(n1102) );
  XNOR2X1 U1116 ( .A(n1107), .B(A[24]), .Y(n1108) );
  OAI22XL U1117 ( .A0(n1121), .A1(n1089), .B0(n5), .B1(n1108), .Y(n1111) );
  XNOR2X1 U1118 ( .A(n1123), .B(A[22]), .Y(n1105) );
  CMPR32X1 U1119 ( .A(n1093), .B(n1092), .C(n1091), .CO(n1109), .S(n1085) );
  CMPR32X1 U1120 ( .A(n1096), .B(n1095), .C(n1094), .CO(n1099), .S(n1084) );
  CMPR32X1 U1121 ( .A(n1101), .B(n1100), .C(n1099), .CO(n1113), .S(n1097) );
  CMPR32X1 U1122 ( .A(n1104), .B(n1103), .C(n1102), .CO(n1130), .S(n1101) );
  XNOR2X1 U1123 ( .A(n1123), .B(A[23]), .Y(n1114) );
  XNOR2X1 U1124 ( .A(n1107), .B(A[25]), .Y(n1119) );
  OAI22X1 U1125 ( .A0(n1121), .A1(n1108), .B0(n5), .B1(n1119), .Y(n1127) );
  CMPR32X1 U1126 ( .A(n1111), .B(n1110), .C(n1109), .CO(n1128), .S(n1100) );
  XNOR2X1 U1127 ( .A(n1123), .B(A[24]), .Y(n1124) );
  CMPR32X1 U1128 ( .A(n1117), .B(n1116), .C(n1115), .CO(n1132), .S(n1129) );
  XNOR2X1 U1129 ( .A(n1123), .B(A[25]), .Y(n1144) );
  CMPR32X1 U1130 ( .A(n1127), .B(n1126), .C(n1125), .CO(n1138), .S(n1131) );
  CMPR32X1 U1131 ( .A(n1130), .B(n1129), .C(n1128), .CO(n1137), .S(n1112) );
  CMPR32X1 U1132 ( .A(n1133), .B(n1132), .C(n1131), .CO(n1135), .S(n1136) );
  CMPR32X1 U1133 ( .A(n1140), .B(n1139), .C(n1138), .CO(n1151), .S(n1134) );
  OAI2BB1X1 U1134 ( .A0N(n106), .A1N(n1146), .B0(n1145), .Y(n1147) );
  XOR3X2 U1135 ( .A(n1149), .B(n1148), .C(n1147), .Y(n1150) );
  OAI21XL U1136 ( .A0(n1159), .A1(n1258), .B0(n1158), .Y(n1229) );
  OAI21XL U1137 ( .A0(n1236), .A1(n1163), .B0(n1162), .Y(n1165) );
  AOI21XL U1138 ( .A0(n1204), .A1(n1167), .B0(n1166), .Y(n1168) );
  OAI21XL U1139 ( .A0(n1236), .A1(n1169), .B0(n1168), .Y(n1172) );
  OAI21XL U1140 ( .A0(n1190), .A1(n1187), .B0(n1188), .Y(n1182) );
  OAI21XL U1141 ( .A0(n1249), .A1(n1252), .B0(n1250), .Y(n1201) );
  AOI21XL U1142 ( .A0(n1204), .A1(n1197), .B0(n1201), .Y(n1183) );
  OAI21XL U1143 ( .A0(n1236), .A1(n1184), .B0(n1183), .Y(n1186) );
  AOI21XL U1144 ( .A0(n1204), .A1(n1203), .B0(n1202), .Y(n1205) );
  OAI21XL U1145 ( .A0(n1236), .A1(n1206), .B0(n1205), .Y(n1209) );
  OAI21XL U1146 ( .A0(n1226), .A1(n1245), .B0(n1246), .Y(n1227) );
  OAI21XL U1147 ( .A0(n1232), .A1(n1231), .B0(n1230), .Y(n1233) );
  OAI21XL U1148 ( .A0(n1236), .A1(n1235), .B0(n1234), .Y(n1237) );
  XNOR2XL U1149 ( .A(n1237), .B(n1244), .Y(PRODUCT[40]) );
  XNOR2XL U1150 ( .A(n1241), .B(n1240), .Y(n1321) );
endmodule


module FFT2048_DW02_mult_2_stage_J1_7 ( A, B, TC, CLK, PRODUCT );
  input [25:0] A;
  input [16:0] B;
  output [42:0] PRODUCT;
  input TC, CLK;
  wire   n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, mult_x_1_n601, mult_x_1_n586, mult_x_1_n569,
         mult_x_1_n554, mult_x_1_n537, mult_x_1_n522, mult_x_1_n321,
         mult_x_1_n316, mult_x_1_n309, mult_x_1_n307, mult_x_1_n306,
         mult_x_1_n296, mult_x_1_n295, mult_x_1_n293, mult_x_1_n292,
         mult_x_1_n287, mult_x_1_n286, mult_x_1_n282, mult_x_1_n281,
         mult_x_1_n277, mult_x_1_n276, mult_x_1_n274, mult_x_1_n273,
         mult_x_1_n266, mult_x_1_n265, mult_x_1_n263, mult_x_1_n262,
         mult_x_1_n245, mult_x_1_n244, mult_x_1_n227, mult_x_1_n226,
         mult_x_1_n207, mult_x_1_n206, mult_x_1_n198, mult_x_1_n197,
         mult_x_1_n195, mult_x_1_n194, mult_x_1_n184, mult_x_1_n183,
         mult_x_1_n177, mult_x_1_n176, mult_x_1_n170, mult_x_1_n169,
         mult_x_1_n161, mult_x_1_n160, mult_x_1_n152, mult_x_1_n151,
         mult_x_1_n137, mult_x_1_n136, mult_x_1_n130, mult_x_1_n129,
         mult_x_1_n121, mult_x_1_n120, mult_x_1_n110, mult_x_1_n109,
         mult_x_1_n86, mult_x_1_n85, mult_x_1_n84, mult_x_1_n83, mult_x_1_n58,
         n5, n6, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415;

  DFFHQXL mult_x_1_clk_r_REG16_S1 ( .D(mult_x_1_n169), .CK(CLK), .Q(n1372) );
  DFFHQXL mult_x_1_clk_r_REG18_S1 ( .D(mult_x_1_n160), .CK(CLK), .Q(n1370) );
  DFFHQX4 mult_x_1_clk_r_REG4_S1 ( .D(mult_x_1_n522), .CK(CLK), .Q(n1410) );
  DFFHQX4 mult_x_1_clk_r_REG50_S1 ( .D(mult_x_1_n296), .CK(CLK), .Q(n1407) );
  DFFHQX4 mult_x_1_clk_r_REG51_S1 ( .D(mult_x_1_n295), .CK(CLK), .Q(n1402) );
  DFFHQX2 mult_x_1_clk_r_REG47_S1 ( .D(mult_x_1_n293), .CK(CLK), .Q(n1401) );
  DFFHQX4 mult_x_1_clk_r_REG48_S1 ( .D(mult_x_1_n292), .CK(CLK), .Q(n1400) );
  DFFHQX4 mult_x_1_clk_r_REG45_S1 ( .D(mult_x_1_n287), .CK(CLK), .Q(n1399) );
  DFFHQX4 mult_x_1_clk_r_REG46_S1 ( .D(mult_x_1_n286), .CK(CLK), .Q(n1398) );
  DFFHQX4 mult_x_1_clk_r_REG44_S1 ( .D(mult_x_1_n281), .CK(CLK), .Q(n1396) );
  DFFHQX4 mult_x_1_clk_r_REG41_S1 ( .D(mult_x_1_n277), .CK(CLK), .Q(n1395) );
  DFFHQX4 mult_x_1_clk_r_REG42_S1 ( .D(mult_x_1_n276), .CK(CLK), .Q(n1394) );
  DFFHQX4 mult_x_1_clk_r_REG40_S1 ( .D(mult_x_1_n273), .CK(CLK), .Q(n1392) );
  DFFHQXL mult_x_1_clk_r_REG49_S1 ( .D(mult_x_1_n83), .CK(CLK), .Q(n1403) );
  DFFHQXL mult_x_1_clk_r_REG19_S1 ( .D(mult_x_1_n152), .CK(CLK), .Q(n1369) );
  DFFHQXL mult_x_1_clk_r_REG20_S1 ( .D(mult_x_1_n151), .CK(CLK), .Q(n1368) );
  DFFHQXL mult_x_1_clk_r_REG60_S1 ( .D(mult_x_1_n321), .CK(CLK), .Q(n1358) );
  DFFHQXL mult_x_1_clk_r_REG17_S1 ( .D(mult_x_1_n161), .CK(CLK), .Q(n1371) );
  DFFHQXL clk_r_REG59_S1 ( .D(n1428), .CK(CLK), .Q(PRODUCT[11]) );
  DFFHQXL mult_x_1_clk_r_REG15_S1 ( .D(mult_x_1_n170), .CK(CLK), .Q(n1373) );
  DFFHQXL mult_x_1_clk_r_REG31_S1 ( .D(mult_x_1_n245), .CK(CLK), .Q(n1387) );
  DFFHQXL mult_x_1_clk_r_REG1_S1 ( .D(mult_x_1_n227), .CK(CLK), .Q(n1385) );
  DFFHQXL mult_x_1_clk_r_REG5_S1 ( .D(mult_x_1_n207), .CK(CLK), .Q(n1383) );
  DFFHQXL clk_r_REG62_S1 ( .D(n1430), .CK(CLK), .Q(PRODUCT[9]) );
  DFFHQXL mult_x_1_clk_r_REG22_S1 ( .D(mult_x_1_n136), .CK(CLK), .Q(n1366) );
  DFFHQX4 mult_x_1_clk_r_REG6_S1 ( .D(mult_x_1_n206), .CK(CLK), .Q(n1382) );
  DFFHQX4 mult_x_1_clk_r_REG43_S1 ( .D(mult_x_1_n282), .CK(CLK), .Q(n1397) );
  DFFHQXL mult_x_1_clk_r_REG8_S1 ( .D(mult_x_1_n197), .CK(CLK), .Q(n1380) );
  DFFHQXL clk_r_REG63_S1 ( .D(n1431), .CK(CLK), .Q(PRODUCT[8]) );
  DFFHQXL clk_r_REG64_S1 ( .D(n1432), .CK(CLK), .Q(PRODUCT[7]) );
  DFFHQXL clk_r_REG65_S1 ( .D(n1433), .CK(CLK), .Q(PRODUCT[6]) );
  DFFHQXL clk_r_REG66_S1 ( .D(n1434), .CK(CLK), .Q(PRODUCT[5]) );
  DFFHQXL clk_r_REG67_S1 ( .D(n1435), .CK(CLK), .Q(PRODUCT[4]) );
  DFFHQXL clk_r_REG68_S1 ( .D(n1436), .CK(CLK), .Q(PRODUCT[3]) );
  DFFHQXL clk_r_REG69_S1 ( .D(n1437), .CK(CLK), .Q(PRODUCT[2]) );
  DFFHQXL clk_r_REG70_S1 ( .D(n1438), .CK(CLK), .Q(PRODUCT[1]) );
  DFFHQXL clk_r_REG71_S1 ( .D(n1439), .CK(CLK), .Q(PRODUCT[0]) );
  DFFHQXL mult_x_1_clk_r_REG58_S1 ( .D(mult_x_1_n316), .CK(CLK), .Q(n1409) );
  DFFHQXL mult_x_1_clk_r_REG57_S1 ( .D(mult_x_1_n86), .CK(CLK), .Q(n1406) );
  DFFHQXL mult_x_1_clk_r_REG52_S1 ( .D(mult_x_1_n84), .CK(CLK), .Q(n1404) );
  DFFHQXL mult_x_1_clk_r_REG7_S1 ( .D(mult_x_1_n198), .CK(CLK), .Q(n1381) );
  DFFHQXL mult_x_1_clk_r_REG10_S1 ( .D(mult_x_1_n194), .CK(CLK), .Q(n1378) );
  DFFHQXL mult_x_1_clk_r_REG11_S1 ( .D(mult_x_1_n184), .CK(CLK), .Q(n1377) );
  DFFHQXL mult_x_1_clk_r_REG12_S1 ( .D(mult_x_1_n183), .CK(CLK), .Q(n1376) );
  DFFHQXL mult_x_1_clk_r_REG13_S1 ( .D(mult_x_1_n177), .CK(CLK), .Q(n1375) );
  DFFHQXL mult_x_1_clk_r_REG14_S1 ( .D(mult_x_1_n176), .CK(CLK), .Q(n1374) );
  DFFHQXL mult_x_1_clk_r_REG21_S1 ( .D(mult_x_1_n137), .CK(CLK), .Q(n1367) );
  DFFHQXL mult_x_1_clk_r_REG23_S1 ( .D(mult_x_1_n130), .CK(CLK), .Q(n1365) );
  DFFHQXL mult_x_1_clk_r_REG24_S1 ( .D(mult_x_1_n129), .CK(CLK), .Q(n1364) );
  DFFHQXL mult_x_1_clk_r_REG25_S1 ( .D(mult_x_1_n121), .CK(CLK), .Q(n1363) );
  DFFHQXL mult_x_1_clk_r_REG26_S1 ( .D(mult_x_1_n120), .CK(CLK), .Q(n1362) );
  DFFHQXL mult_x_1_clk_r_REG27_S1 ( .D(mult_x_1_n110), .CK(CLK), .Q(n1361) );
  DFFHQXL mult_x_1_clk_r_REG28_S1 ( .D(mult_x_1_n109), .CK(CLK), .Q(n1360) );
  DFFHQXL mult_x_1_clk_r_REG29_S1 ( .D(mult_x_1_n58), .CK(CLK), .Q(n1359) );
  DFFHQXL mult_x_1_clk_r_REG53_S1 ( .D(mult_x_1_n307), .CK(CLK), .Q(n1357) );
  DFFHQXL mult_x_1_clk_r_REG54_S1 ( .D(mult_x_1_n306), .CK(CLK), .Q(n1356) );
  DFFHQXL clk_r_REG61_S1 ( .D(n1429), .CK(CLK), .Q(PRODUCT[10]) );
  DFFHQXL mult_x_1_clk_r_REG9_S1 ( .D(mult_x_1_n195), .CK(CLK), .Q(n1379) );
  DFFHQX4 mult_x_1_clk_r_REG56_S1 ( .D(mult_x_1_n309), .CK(CLK), .Q(n1408) );
  DFFHQXL mult_x_1_clk_r_REG32_S1 ( .D(mult_x_1_n244), .CK(CLK), .Q(n1386) );
  DFFHQXL mult_x_1_clk_r_REG2_S1 ( .D(mult_x_1_n226), .CK(CLK), .Q(n1384) );
  DFFHQX1 mult_x_1_clk_r_REG36_S1 ( .D(mult_x_1_n262), .CK(CLK), .Q(n1388) );
  DFFHQX1 mult_x_1_clk_r_REG38_S1 ( .D(mult_x_1_n265), .CK(CLK), .Q(n1390) );
  DFFHQXL mult_x_1_clk_r_REG35_S1 ( .D(mult_x_1_n263), .CK(CLK), .Q(n1389) );
  DFFHQXL mult_x_1_clk_r_REG55_S1 ( .D(mult_x_1_n85), .CK(CLK), .Q(n1405) );
  DFFHQX1 mult_x_1_clk_r_REG30_S1 ( .D(mult_x_1_n569), .CK(CLK), .Q(n1413) );
  DFFHQX2 mult_x_1_clk_r_REG0_S1 ( .D(mult_x_1_n554), .CK(CLK), .Q(n1412) );
  DFFHQX1 mult_x_1_clk_r_REG33_S1 ( .D(mult_x_1_n586), .CK(CLK), .Q(n1414) );
  DFFHQX1 mult_x_1_clk_r_REG3_S1 ( .D(mult_x_1_n537), .CK(CLK), .Q(n1411) );
  DFFHQX1 mult_x_1_clk_r_REG34_S1 ( .D(mult_x_1_n601), .CK(CLK), .Q(n1415) );
  DFFHQX1 mult_x_1_clk_r_REG37_S1 ( .D(mult_x_1_n266), .CK(CLK), .Q(n1391) );
  DFFHQX2 mult_x_1_clk_r_REG39_S1 ( .D(mult_x_1_n274), .CK(CLK), .Q(n1393) );
  CMPR32X1 U1 ( .A(n430), .B(n429), .C(n428), .CO(n403), .S(n431) );
  CMPR32X1 U2 ( .A(n1198), .B(n1197), .C(n1196), .CO(n1230), .S(n402) );
  OAI21XL U3 ( .A0(n42), .A1(n41), .B0(n40), .Y(n874) );
  ADDFHX1 U4 ( .A(n1174), .B(n1173), .CI(n1172), .CO(mult_x_1_n601), .S(n842)
         );
  ADDFHX1 U5 ( .A(n1162), .B(n1161), .CI(n1160), .CO(mult_x_1_n537), .S(n715)
         );
  ADDFHX1 U6 ( .A(n609), .B(n608), .CI(n607), .CO(n567), .S(n610) );
  ADDFHX1 U7 ( .A(n1159), .B(n1158), .CI(n1157), .CO(n646), .S(mult_x_1_n522)
         );
  ADDFHX2 U8 ( .A(n840), .B(n839), .CI(n838), .CO(n1173), .S(n844) );
  OAI21X2 U9 ( .A0(n171), .A1(n172), .B0(n170), .Y(n845) );
  ADDFHX1 U10 ( .A(n811), .B(n810), .CI(n809), .CO(n1170), .S(n1172) );
  ADDFHX1 U11 ( .A(n686), .B(n685), .CI(n684), .CO(n1158), .S(n1160) );
  ADDFHX1 U12 ( .A(n713), .B(n712), .CI(n711), .CO(n1161), .S(n1163) );
  ADDFHX1 U13 ( .A(n808), .B(n807), .CI(n806), .CO(n811), .S(n838) );
  ADDFHX1 U14 ( .A(n805), .B(n804), .CI(n803), .CO(n1174), .S(n839) );
  CMPR32X1 U15 ( .A(n1035), .B(n1034), .C(n1033), .CO(n1022), .S(n1105) );
  CMPR32X1 U16 ( .A(n529), .B(n528), .C(n527), .CO(n532), .S(n557) );
  ADDFX2 U17 ( .A(n496), .B(n495), .CI(n494), .CO(n514), .S(n530) );
  ADDFHX1 U18 ( .A(n1087), .B(n1086), .CI(n1085), .CO(n1104), .S(n1106) );
  ADDFHX1 U19 ( .A(n747), .B(n746), .CI(n745), .CO(n749), .S(n772) );
  ADDFHX1 U20 ( .A(n788), .B(n787), .CI(n786), .CO(n768), .S(n804) );
  ADDFHX2 U21 ( .A(n871), .B(n870), .CI(n869), .CO(n873), .S(n914) );
  ADDFHX2 U22 ( .A(n913), .B(n912), .CI(n911), .CO(n916), .S(n950) );
  ADDFHX1 U23 ( .A(n1071), .B(n1070), .CI(n1069), .CO(n1064), .S(n1108) );
  ADDFHX1 U24 ( .A(n934), .B(n933), .CI(n932), .CO(n941), .S(n973) );
  CMPR32X1 U25 ( .A(n727), .B(n726), .C(n725), .CO(n707), .S(n743) );
  ADDFHX1 U26 ( .A(n526), .B(n525), .CI(n524), .CO(n518), .S(n558) );
  ADDFHX2 U27 ( .A(n828), .B(n827), .CI(n826), .CO(n837), .S(n870) );
  CMPR32X1 U28 ( .A(n1074), .B(n1073), .C(n1072), .CO(n1087), .S(n1102) );
  OAI21XL U29 ( .A0(n126), .A1(n125), .B0(n124), .Y(n710) );
  ADDFHX1 U30 ( .A(n1137), .B(n1136), .CI(n1135), .CO(n1128), .S(n1143) );
  ADDFHX1 U31 ( .A(n901), .B(n900), .CI(n899), .CO(n913), .S(n939) );
  ADDFHX1 U32 ( .A(n893), .B(n892), .CI(n891), .CO(n871), .S(n924) );
  CMPR32X1 U33 ( .A(n1124), .B(n1123), .C(n1122), .CO(n1136), .S(n1138) );
  OAI22X1 U34 ( .A0(n1203), .A1(n823), .B0(n1052), .B1(n794), .Y(n828) );
  OAI22X1 U35 ( .A0(n1203), .A1(n903), .B0(n1052), .B1(n857), .Y(n901) );
  OAI21X1 U36 ( .A0(n697), .A1(n1052), .B0(n64), .Y(n63) );
  ADDFHX1 U37 ( .A(n1127), .B(n1126), .CI(n1125), .CO(n1117), .S(n1135) );
  ADDFHX1 U38 ( .A(n340), .B(n339), .CI(n338), .CO(n1139), .S(n348) );
  ADDFHX1 U39 ( .A(n306), .B(n305), .CI(n304), .CO(n328), .S(n307) );
  BUFX8 U40 ( .A(n931), .Y(n1262) );
  CLKBUFX8 U41 ( .A(n372), .Y(n1263) );
  BUFX4 U42 ( .A(n581), .Y(n11) );
  BUFX4 U43 ( .A(n450), .Y(n1259) );
  CLKBUFX8 U44 ( .A(B[13]), .Y(n1205) );
  CLKBUFX8 U45 ( .A(n365), .Y(n1243) );
  OAI22X2 U46 ( .A0(n729), .A1(n293), .B0(n1078), .B1(n292), .Y(n102) );
  XOR2X1 U47 ( .A(B[6]), .B(B[7]), .Y(n142) );
  OAI21X1 U48 ( .A0(n285), .A1(n1080), .B0(n79), .Y(n113) );
  XNOR2X2 U49 ( .A(B[6]), .B(B[5]), .Y(n227) );
  INVX4 U50 ( .A(n483), .Y(n12) );
  XNOR2X2 U51 ( .A(B[10]), .B(B[9]), .Y(n336) );
  XOR2XL U52 ( .A(n32), .B(n508), .Y(PRODUCT[31]) );
  XOR2X1 U53 ( .A(n20), .B(n536), .Y(PRODUCT[30]) );
  XOR2X1 U54 ( .A(n620), .B(n619), .Y(PRODUCT[28]) );
  XOR2X1 U55 ( .A(n29), .B(n782), .Y(PRODUCT[23]) );
  XNOR2X1 U56 ( .A(n653), .B(n652), .Y(PRODUCT[27]) );
  XOR2X1 U57 ( .A(n19), .B(n880), .Y(PRODUCT[20]) );
  AOI2BB1X2 U58 ( .A0N(n876), .A1N(n191), .B0(n877), .Y(n220) );
  OAI21X2 U59 ( .A0(n876), .A1(n190), .B0(n167), .Y(n613) );
  INVXL U60 ( .A(n1120), .Y(n5) );
  INVXL U61 ( .A(n5), .Y(n6) );
  OAI22X1 U62 ( .A0(n1050), .A1(n1049), .B0(n1048), .B1(n1175), .Y(n1084) );
  OAI22X1 U63 ( .A0(n965), .A1(n287), .B0(n194), .B1(n318), .Y(n325) );
  OAI22X1 U64 ( .A0(n174), .A1(n592), .B0(n1058), .B1(n549), .Y(n595) );
  OAI22X1 U65 ( .A0(n1050), .A1(n323), .B0(n334), .B1(n1175), .Y(n341) );
  OAI22X1 U66 ( .A0(n729), .A1(n488), .B0(n1078), .B1(n481), .Y(n520) );
  XOR2X1 U67 ( .A(n1182), .B(n843), .Y(PRODUCT[21]) );
  XNOR2XL U68 ( .A(n1295), .B(n1294), .Y(PRODUCT[38]) );
  XNOR2XL U69 ( .A(n1037), .B(n1176), .Y(n232) );
  XNOR2XL U70 ( .A(n1013), .B(n1176), .Y(n285) );
  XNOR2XL U71 ( .A(n1205), .B(A[17]), .Y(n449) );
  XNOR2XL U72 ( .A(n1013), .B(A[3]), .Y(n1079) );
  XNOR2XL U73 ( .A(n1205), .B(n1036), .Y(n848) );
  XOR2XL U74 ( .A(n238), .B(n982), .Y(n1018) );
  XOR2XL U75 ( .A(n238), .B(n1199), .Y(n629) );
  XNOR2XL U76 ( .A(n884), .B(A[18]), .Y(n374) );
  XNOR2XL U77 ( .A(n884), .B(A[16]), .Y(n367) );
  BUFX3 U78 ( .A(n965), .Y(n1063) );
  BUFX1 U79 ( .A(A[1]), .Y(n970) );
  XNOR2XL U80 ( .A(n578), .B(n577), .Y(n586) );
  XNOR2XL U81 ( .A(n1250), .B(A[11]), .Y(n580) );
  XNOR2XL U82 ( .A(n1250), .B(n984), .Y(n750) );
  XNOR2XL U83 ( .A(n945), .B(n90), .Y(n1002) );
  OAI21X2 U84 ( .A0(n145), .A1(n144), .B0(n143), .Y(n922) );
  ADDFX2 U85 ( .A(n424), .B(n423), .CI(n422), .CO(n466), .S(n461) );
  XOR2XL U86 ( .A(n1306), .B(n1305), .Y(n1433) );
  INVX1 U87 ( .A(n1060), .Y(n8) );
  BUFX1 U88 ( .A(n1060), .Y(n173) );
  INVX4 U89 ( .A(B[5]), .Y(n238) );
  ADDFX2 U90 ( .A(n941), .B(n940), .CI(n939), .CO(n952), .S(n992) );
  XNOR2XL U91 ( .A(n31), .B(n178), .Y(PRODUCT[29]) );
  NAND2X1 U92 ( .A(n1187), .B(n14), .Y(n95) );
  INVX1 U93 ( .A(n1188), .Y(n14) );
  NAND2XL U94 ( .A(n1189), .B(n1195), .Y(n1191) );
  INVX1 U95 ( .A(n331), .Y(n46) );
  NOR2X1 U96 ( .A(n610), .B(n611), .Y(mult_x_1_n197) );
  NOR2XL U97 ( .A(n875), .B(n874), .Y(mult_x_1_n265) );
  NAND2BX1 U98 ( .AN(n1129), .B(n153), .Y(n1189) );
  OAI21XL U99 ( .A0(n1065), .A1(n1066), .B0(n1064), .Y(n148) );
  NAND2X1 U100 ( .A(n1129), .B(n1128), .Y(n1187) );
  INVX1 U101 ( .A(n1128), .Y(n153) );
  INVX1 U102 ( .A(n1143), .Y(n84) );
  INVX1 U103 ( .A(n681), .Y(n132) );
  INVXL U104 ( .A(n837), .Y(n188) );
  INVXL U105 ( .A(n499), .Y(n82) );
  NAND2BX1 U106 ( .AN(n324), .B(n10), .Y(n79) );
  OR2X2 U107 ( .A(n333), .B(n1078), .Y(n108) );
  INVXL U108 ( .A(n11), .Y(n184) );
  OAI22X1 U109 ( .A0(n1063), .A1(n1061), .B0(n194), .B1(n1018), .Y(n1075) );
  OAI22X1 U110 ( .A0(n11), .A1(n990), .B0(n1243), .B1(n989), .Y(n1046) );
  NOR2X1 U111 ( .A(n1259), .B(n600), .Y(n665) );
  INVXL U112 ( .A(n701), .Y(n125) );
  NOR2X1 U113 ( .A(n1259), .B(n451), .Y(n492) );
  OAI22X1 U114 ( .A0(n176), .A1(n1057), .B0(n1058), .B1(n1016), .Y(n1076) );
  NOR2X1 U115 ( .A(n1259), .B(n696), .Y(n730) );
  NAND2BXL U116 ( .AN(n177), .B(n51), .Y(n50) );
  NAND2X1 U117 ( .A(B[5]), .B(n13), .Y(n237) );
  INVX1 U118 ( .A(n123), .Y(n122) );
  XOR2X1 U119 ( .A(n238), .B(n970), .Y(n246) );
  XOR2X1 U120 ( .A(n238), .B(A[2]), .Y(n233) );
  XOR2X1 U121 ( .A(n238), .B(A[3]), .Y(n288) );
  NAND2XL U122 ( .A(n48), .B(n51), .Y(n47) );
  XOR2X1 U123 ( .A(n238), .B(n1221), .Y(n593) );
  XOR2X1 U124 ( .A(n238), .B(n967), .Y(n859) );
  XOR2X1 U125 ( .A(n238), .B(n927), .Y(n204) );
  XNOR2XL U126 ( .A(n884), .B(A[17]), .Y(n366) );
  XOR2X1 U127 ( .A(n12), .B(n984), .Y(n51) );
  NAND2X1 U128 ( .A(n39), .B(n470), .Y(n474) );
  AOI21X1 U129 ( .A0(n31), .A1(n505), .B0(n506), .Y(n32) );
  OAI21XL U130 ( .A0(n1181), .A1(n1182), .B0(n1180), .Y(n1186) );
  NAND2XL U131 ( .A(n30), .B(n778), .Y(n29) );
  INVX1 U132 ( .A(n405), .Y(n406) );
  NAND2BXL U133 ( .AN(n779), .B(n613), .Y(n30) );
  INVX1 U134 ( .A(n1183), .Y(n17) );
  INVX1 U135 ( .A(n650), .Y(n18) );
  NAND2X1 U136 ( .A(n507), .B(n1377), .Y(n508) );
  NAND2X1 U137 ( .A(n568), .B(n1381), .Y(n178) );
  NAND2X1 U138 ( .A(n721), .B(n1387), .Y(n722) );
  NAND2XL U139 ( .A(n996), .B(n1399), .Y(n997) );
  INVX1 U140 ( .A(n1176), .Y(n13) );
  INVXL U141 ( .A(n1017), .Y(n121) );
  NAND2BXL U142 ( .AN(n1356), .B(n1408), .Y(n213) );
  NAND2X1 U143 ( .A(n1410), .B(n1411), .Y(n651) );
  BUFX2 U144 ( .A(A[21]), .Y(n1221) );
  NAND2X1 U145 ( .A(n1134), .B(n15), .Y(n54) );
  NOR2X1 U146 ( .A(n84), .B(n96), .Y(n1188) );
  NAND2X1 U147 ( .A(n331), .B(n330), .Y(n1145) );
  INVX1 U148 ( .A(n1147), .Y(n1156) );
  OAI21XL U149 ( .A0(n748), .A1(n749), .B0(n68), .Y(n67) );
  INVXL U150 ( .A(n330), .Y(n45) );
  OAI2BB1X1 U151 ( .A0N(n81), .A1N(n497), .B0(n80), .Y(n501) );
  NAND2BXL U152 ( .AN(n710), .B(n136), .Y(n135) );
  OAI21XL U153 ( .A0(n682), .A1(n683), .B0(n681), .Y(n131) );
  INVX1 U154 ( .A(n709), .Y(n136) );
  OAI2BB1X1 U155 ( .A0N(n188), .A1N(n73), .B0(n835), .Y(n72) );
  NAND2X1 U156 ( .A(n280), .B(n279), .Y(n1303) );
  OR2X2 U157 ( .A(n320), .B(n321), .Y(n141) );
  NAND2X1 U158 ( .A(n320), .B(n321), .Y(n140) );
  ADDFHX1 U159 ( .A(n1088), .B(n1089), .CI(n1090), .CO(n1085), .S(n1118) );
  NAND2XL U160 ( .A(n130), .B(n341), .Y(n159) );
  NAND2XL U161 ( .A(n573), .B(n118), .Y(n114) );
  ADDFHX1 U162 ( .A(n851), .B(n850), .CI(n849), .CO(n834), .S(n867) );
  ADDFHX1 U163 ( .A(n691), .B(n690), .CI(n689), .CO(n680), .S(n706) );
  ADDFHX1 U164 ( .A(n663), .B(n662), .CI(n661), .CO(n641), .S(n679) );
  NAND2BXL U165 ( .AN(n569), .B(n193), .Y(n195) );
  ADDFHX1 U166 ( .A(n817), .B(n816), .CI(n815), .CO(n805), .S(n833) );
  NAND2XL U167 ( .A(n184), .B(n183), .Y(n182) );
  OAI22X1 U168 ( .A0(n1262), .A1(n1251), .B0(n1263), .B1(n1260), .Y(n1266) );
  OAI21XL U169 ( .A0(n1058), .A1(n347), .B0(n50), .Y(n342) );
  OR2X2 U170 ( .A(n548), .B(n1204), .Y(n60) );
  NAND2XL U171 ( .A(n106), .B(n105), .Y(n104) );
  OAI22X1 U172 ( .A0(n231), .A1(n812), .B0(n1055), .B1(n783), .Y(n817) );
  NOR2X1 U173 ( .A(n1259), .B(n374), .Y(n395) );
  NOR2X1 U174 ( .A(n1259), .B(n435), .Y(n457) );
  NOR2BX1 U175 ( .AN(n1176), .B(n1263), .Y(n1012) );
  NAND2BXL U176 ( .AN(n760), .B(n16), .Y(n198) );
  NOR2X1 U177 ( .A(n1259), .B(n793), .Y(n819) );
  NOR2X1 U178 ( .A(n1259), .B(n668), .Y(n693) );
  INVXL U179 ( .A(n183), .Y(n181) );
  NOR2X1 U180 ( .A(n1259), .B(n367), .Y(n421) );
  NOR2X1 U181 ( .A(n1259), .B(n366), .Y(n387) );
  NOR2X1 U182 ( .A(n1259), .B(n1200), .Y(n1219) );
  NOR2X1 U183 ( .A(n1259), .B(n1222), .Y(n1237) );
  NOR2X1 U184 ( .A(n1259), .B(n1249), .Y(n1257) );
  NOR2X1 U185 ( .A(n1259), .B(n1240), .Y(n1253) );
  NOR2X1 U186 ( .A(n1259), .B(n885), .Y(n906) );
  NOR2X1 U187 ( .A(n1259), .B(n856), .Y(n889) );
  NOR2X1 U188 ( .A(n1259), .B(n413), .Y(n440) );
  NAND2X1 U189 ( .A(n49), .B(n47), .Y(n321) );
  NOR2X1 U190 ( .A(n1259), .B(n390), .Y(n1209) );
  NOR2X1 U191 ( .A(n1259), .B(n822), .Y(n853) );
  XOR2X1 U192 ( .A(n238), .B(A[11]), .Y(n964) );
  INVX1 U193 ( .A(n1052), .Y(n9) );
  XOR2X1 U194 ( .A(n238), .B(A[18]), .Y(n699) );
  XOR2X1 U195 ( .A(n238), .B(A[17]), .Y(n736) );
  XOR2X1 U196 ( .A(n238), .B(n1015), .Y(n983) );
  XOR2X1 U197 ( .A(n238), .B(n894), .Y(n796) );
  XOR2X1 U198 ( .A(n238), .B(A[16]), .Y(n760) );
  XNOR2X1 U199 ( .A(n1286), .B(n1285), .Y(PRODUCT[37]) );
  OR2X2 U200 ( .A(n173), .B(n291), .Y(n49) );
  XOR2X1 U201 ( .A(n238), .B(n1176), .Y(n247) );
  XOR2X1 U202 ( .A(n238), .B(A[19]), .Y(n671) );
  XOR2X1 U203 ( .A(n238), .B(n1017), .Y(n1061) );
  XNOR2X1 U204 ( .A(n1291), .B(n1290), .Y(PRODUCT[36]) );
  XOR2X1 U205 ( .A(n238), .B(n986), .Y(n902) );
  INVX1 U206 ( .A(n1078), .Y(n10) );
  XNOR2X1 U207 ( .A(n474), .B(n473), .Y(PRODUCT[32]) );
  XNOR2X1 U208 ( .A(n363), .B(n362), .Y(PRODUCT[35]) );
  XNOR2X1 U209 ( .A(n1319), .B(n1318), .Y(PRODUCT[39]) );
  XOR2X1 U210 ( .A(n33), .B(n434), .Y(PRODUCT[33]) );
  INVX1 U211 ( .A(n1058), .Y(n48) );
  NAND2X1 U212 ( .A(n230), .B(n257), .Y(n1060) );
  OAI22X1 U213 ( .A0(n988), .A1(n235), .B0(n228), .B1(n1175), .Y(n240) );
  AOI21XL U214 ( .A0(n1179), .A1(n615), .B0(n26), .Y(n616) );
  OAI21XL U215 ( .A0(n1182), .A1(n649), .B0(n648), .Y(n653) );
  NAND2XL U216 ( .A(n27), .B(n651), .Y(n26) );
  NOR2X1 U217 ( .A(n1340), .B(n1280), .Y(n1308) );
  NAND2X1 U218 ( .A(n614), .B(n18), .Y(n27) );
  NAND2X1 U219 ( .A(n28), .B(n1385), .Y(n614) );
  AND2X2 U220 ( .A(n18), .B(n612), .Y(n615) );
  NAND2BX1 U221 ( .AN(n1384), .B(n17), .Y(n28) );
  INVX1 U222 ( .A(n654), .Y(n1184) );
  INVX1 U223 ( .A(n894), .Y(n56) );
  INVX1 U224 ( .A(A[16]), .Y(n139) );
  NAND2X1 U225 ( .A(n1273), .B(n1371), .Y(n408) );
  OAI21XL U226 ( .A0(n1378), .A1(n1381), .B0(n1379), .Y(n506) );
  INVX1 U227 ( .A(n1370), .Y(n1273) );
  INVX1 U228 ( .A(n1380), .Y(n568) );
  BUFX2 U229 ( .A(A[15]), .Y(n894) );
  BUFX2 U230 ( .A(A[14]), .Y(n927) );
  BUFX2 U231 ( .A(A[22]), .Y(n1239) );
  XOR2X1 U232 ( .A(n1409), .B(n1405), .Y(PRODUCT[13]) );
  INVX1 U233 ( .A(n1144), .Y(n15) );
  NOR2X1 U234 ( .A(n995), .B(n994), .Y(mult_x_1_n281) );
  ADDFHX2 U235 ( .A(n960), .B(n959), .CI(n958), .CO(n953), .S(n995) );
  NAND2X1 U236 ( .A(n351), .B(n352), .Y(n1130) );
  OAI2BB1X1 U237 ( .A0N(n1066), .A1N(n1065), .B0(n148), .Y(n1031) );
  NAND2X1 U238 ( .A(n1110), .B(n1109), .Y(mult_x_1_n307) );
  NAND2X1 U239 ( .A(n67), .B(n66), .Y(n1164) );
  NOR2X1 U240 ( .A(n647), .B(n646), .Y(mult_x_1_n206) );
  ADDFHX2 U241 ( .A(n1168), .B(n1167), .CI(n1166), .CO(mult_x_1_n569), .S(n776) );
  XNOR2X1 U242 ( .A(n1301), .B(n1300), .Y(n1432) );
  NAND2XL U243 ( .A(n534), .B(n533), .Y(mult_x_1_n184) );
  ADDFHX2 U244 ( .A(n623), .B(n622), .CI(n621), .CO(n611), .S(n647) );
  ADDFHX1 U245 ( .A(n1108), .B(n1107), .CI(n1106), .CO(n1111), .S(n1110) );
  XOR2X1 U246 ( .A(n86), .B(n1064), .Y(n1103) );
  XOR2X1 U247 ( .A(n69), .B(n68), .Y(n1166) );
  XOR2X1 U248 ( .A(n748), .B(n749), .Y(n69) );
  OAI2BB1X1 U249 ( .A0N(n135), .A1N(n708), .B0(n134), .Y(n713) );
  NAND2X1 U250 ( .A(n748), .B(n749), .Y(n66) );
  ADDFHX2 U251 ( .A(n846), .B(n845), .CI(n844), .CO(n841), .S(n875) );
  NAND2X1 U252 ( .A(n498), .B(n499), .Y(n80) );
  INVX1 U253 ( .A(n710), .Y(n137) );
  OAI2BB1X1 U254 ( .A0N(n683), .A1N(n682), .B0(n131), .Y(n686) );
  ADDFHX2 U255 ( .A(n547), .B(n546), .CI(n545), .CO(n563), .S(n608) );
  NAND2X1 U256 ( .A(n72), .B(n187), .Y(n840) );
  OAI2BB1X1 U257 ( .A0N(n738), .A1N(n63), .B0(n62), .Y(n747) );
  NAND2XL U258 ( .A(n207), .B(n206), .Y(n766) );
  NOR2X1 U259 ( .A(n1297), .B(n1302), .Y(n283) );
  OAI2BB1X1 U260 ( .A0N(n141), .A1N(n319), .B0(n140), .Y(n349) );
  NAND2BX1 U261 ( .AN(n498), .B(n82), .Y(n81) );
  INVX1 U262 ( .A(n882), .Y(n44) );
  XOR2X1 U263 ( .A(n166), .B(n519), .Y(n547) );
  OR2XL U264 ( .A(n1268), .B(n1267), .Y(n1270) );
  NAND2BXL U265 ( .AN(n91), .B(n946), .Y(n88) );
  XOR2X1 U266 ( .A(n1065), .B(n1066), .Y(n86) );
  XOR3X2 U267 ( .A(n701), .B(n127), .C(n700), .Y(n746) );
  OAI2BB1XL U268 ( .A0N(n150), .A1N(n752), .B0(n149), .Y(n744) );
  XOR3X2 U269 ( .A(n1076), .B(n100), .C(n1075), .Y(n1101) );
  NAND2X1 U270 ( .A(n58), .B(n57), .Y(n626) );
  INVX1 U271 ( .A(n113), .Y(n112) );
  NOR2X1 U272 ( .A(n282), .B(n281), .Y(n1297) );
  XOR3X2 U273 ( .A(n325), .B(n113), .C(n326), .Y(n329) );
  OAI2BB1X1 U274 ( .A0N(n160), .A1N(n107), .B0(n159), .Y(n1124) );
  NAND2BXL U275 ( .AN(n573), .B(n116), .Y(n115) );
  INVX1 U276 ( .A(n836), .Y(n73) );
  NAND2BXL U277 ( .AN(n753), .B(n151), .Y(n150) );
  XOR2X1 U278 ( .A(n572), .B(n117), .Y(n590) );
  INVX1 U279 ( .A(n127), .Y(n126) );
  XOR2X1 U280 ( .A(n61), .B(n59), .Y(n637) );
  OAI21XL U281 ( .A0(n1080), .A1(n120), .B0(n119), .Y(n909) );
  ADDFHX1 U282 ( .A(n1021), .B(n1020), .CI(n1019), .CO(n1035), .S(n1069) );
  NAND2BXL U283 ( .AN(n671), .B(n193), .Y(n202) );
  NAND2BXL U284 ( .AN(n629), .B(n193), .Y(n197) );
  ADDFHX1 U285 ( .A(n241), .B(n240), .CI(n239), .CO(n311), .S(n242) );
  NAND2BXL U286 ( .AN(n699), .B(n193), .Y(n201) );
  NAND2BX1 U287 ( .AN(n1014), .B(n10), .Y(n101) );
  AND2X2 U288 ( .A(n85), .B(n966), .Y(n974) );
  NAND2BX1 U289 ( .AN(n734), .B(n65), .Y(n64) );
  NAND2BXL U290 ( .AN(n736), .B(n193), .Y(n200) );
  INVXL U291 ( .A(n420), .Y(n441) );
  OAI21XL U292 ( .A0(n783), .A1(n231), .B0(n104), .Y(n788) );
  NAND2BXL U293 ( .AN(n760), .B(n193), .Y(n199) );
  INVXL U294 ( .A(n519), .Y(n165) );
  INVXL U295 ( .A(n539), .Y(n551) );
  OAI2BB1XL U296 ( .A0N(n194), .A1N(n1063), .B0(n437), .Y(n455) );
  INVXL U297 ( .A(n158), .Y(n156) );
  XOR2X1 U298 ( .A(n595), .B(n594), .Y(n61) );
  INVX1 U299 ( .A(n105), .Y(n103) );
  NAND2X1 U300 ( .A(n1176), .B(n9), .Y(n161) );
  NOR2XL U301 ( .A(n1259), .B(n1258), .Y(n1265) );
  AND2XL U302 ( .A(n1323), .B(n1322), .Y(n1438) );
  XNOR2XL U303 ( .A(n884), .B(n1239), .Y(n1240) );
  OR2XL U304 ( .A(n1321), .B(n1320), .Y(n1323) );
  XNOR2XL U305 ( .A(n884), .B(A[23]), .Y(n1249) );
  XNOR2XL U306 ( .A(n884), .B(n1199), .Y(n1200) );
  CLKINVX3 U307 ( .A(n930), .Y(n1234) );
  NAND2X1 U308 ( .A(n31), .B(n471), .Y(n39) );
  AOI2BB1X1 U309 ( .A0N(n655), .A1N(n1182), .B0(n37), .Y(n36) );
  INVX1 U310 ( .A(n194), .Y(n16) );
  NAND2X1 U311 ( .A(B[1]), .B(n968), .Y(n1050) );
  INVXL U312 ( .A(n179), .Y(n1181) );
  AND2X2 U313 ( .A(n781), .B(n780), .Y(n782) );
  INVX1 U314 ( .A(n35), .Y(n21) );
  AND2XL U315 ( .A(n505), .B(n507), .Y(n471) );
  INVX1 U316 ( .A(n1015), .Y(n71) );
  AND2X2 U317 ( .A(n618), .B(n1383), .Y(n619) );
  AND2X2 U318 ( .A(n879), .B(n1393), .Y(n880) );
  NOR2X1 U319 ( .A(n1398), .B(n1396), .Y(n878) );
  INVXL U320 ( .A(n1381), .Y(n215) );
  BUFX2 U321 ( .A(A[10]), .Y(n1015) );
  BUFX2 U322 ( .A(A[9]), .Y(n982) );
  INVXL U323 ( .A(A[11]), .Y(n210) );
  BUFX2 U324 ( .A(A[20]), .Y(n1199) );
  INVXL U325 ( .A(n1398), .Y(n996) );
  BUFX2 U326 ( .A(A[6]), .Y(n1036) );
  BUFX2 U327 ( .A(A[5]), .Y(n975) );
  BUFX2 U328 ( .A(A[12]), .Y(n986) );
  BUFX2 U329 ( .A(A[13]), .Y(n967) );
  INVXL U330 ( .A(n1391), .Y(n218) );
  OAI21XL U331 ( .A0(n220), .A1(n1394), .B0(n1395), .Y(n19) );
  AOI21X4 U332 ( .A0(n1408), .A1(n169), .B0(n168), .Y(n876) );
  AOI21X1 U333 ( .A0(n31), .A1(n568), .B0(n215), .Y(n20) );
  NAND4X2 U334 ( .A(n25), .B(n23), .C(n22), .D(n21), .Y(n31) );
  NAND2X1 U335 ( .A(n614), .B(n357), .Y(n22) );
  NAND3X1 U336 ( .A(n214), .B(n179), .C(n613), .Y(n23) );
  NOR2BX1 U337 ( .AN(n612), .B(n24), .Y(n214) );
  INVX1 U338 ( .A(n357), .Y(n24) );
  NAND2X1 U339 ( .A(n214), .B(n1179), .Y(n25) );
  NOR2X1 U340 ( .A(n1411), .B(n1410), .Y(n650) );
  NOR2X2 U341 ( .A(n1384), .B(n654), .Y(n612) );
  CLKINVX3 U342 ( .A(n613), .Y(n1182) );
  INVX1 U343 ( .A(n31), .Y(n1350) );
  AOI21X1 U344 ( .A0(n31), .A1(n189), .B0(n34), .Y(n33) );
  INVX1 U345 ( .A(n1347), .Y(n34) );
  OAI21XL U346 ( .A0(n1382), .A1(n651), .B0(n1383), .Y(n35) );
  NAND2BX2 U347 ( .AN(n222), .B(n221), .Y(n1179) );
  XOR2X2 U348 ( .A(n36), .B(n657), .Y(PRODUCT[26]) );
  NAND2X1 U349 ( .A(n38), .B(n1183), .Y(n37) );
  NAND2X1 U350 ( .A(n1179), .B(n1184), .Y(n38) );
  NOR2X1 U351 ( .A(n1386), .B(n716), .Y(n356) );
  OAI21XL U352 ( .A0(n1350), .A1(n407), .B0(n406), .Y(n409) );
  XNOR2X1 U353 ( .A(n409), .B(n408), .Y(PRODUCT[34]) );
  AND2X2 U354 ( .A(n356), .B(n777), .Y(n179) );
  OAI22X1 U355 ( .A0(n1203), .A1(n857), .B0(n1052), .B1(n823), .Y(n893) );
  XOR2X1 U356 ( .A(n643), .B(n642), .Y(n644) );
  XOR2X1 U357 ( .A(n645), .B(n644), .Y(n1157) );
  XOR2X1 U358 ( .A(n573), .B(n118), .Y(n117) );
  NAND2X1 U359 ( .A(n1026), .B(n1025), .Y(mult_x_1_n287) );
  NOR2BX1 U360 ( .AN(n1176), .B(n1259), .Y(n934) );
  XOR3X2 U361 ( .A(n993), .B(n992), .C(n991), .Y(n998) );
  XNOR2X2 U362 ( .A(n1041), .B(n1017), .Y(n823) );
  NAND2BX1 U363 ( .AN(n669), .B(n9), .Y(n128) );
  NOR2X1 U364 ( .A(n1259), .B(n758), .Y(n790) );
  INVX4 U365 ( .A(B[7]), .Y(n368) );
  INVX1 U366 ( .A(n43), .Y(n41) );
  NAND2X1 U367 ( .A(n954), .B(n953), .Y(mult_x_1_n277) );
  BUFX12 U368 ( .A(n335), .Y(n1203) );
  OAI22X1 U369 ( .A0(n1203), .A1(n669), .B0(n1204), .B1(n627), .Y(n674) );
  XNOR2X1 U370 ( .A(n497), .B(n83), .Y(n509) );
  AOI21X1 U371 ( .A0(n1194), .A1(n1114), .B0(n1113), .Y(mult_x_1_n296) );
  XNOR2X1 U372 ( .A(n1234), .B(A[16]), .Y(n445) );
  AOI21X1 U373 ( .A0(n1134), .A1(n1133), .B0(n1132), .Y(n1192) );
  NAND2X1 U374 ( .A(n918), .B(n917), .Y(mult_x_1_n274) );
  INVX8 U375 ( .A(n293), .Y(n1013) );
  NAND2X1 U376 ( .A(n881), .B(n882), .Y(n40) );
  NOR2X1 U377 ( .A(n881), .B(n882), .Y(n42) );
  XNOR3X2 U378 ( .A(n44), .B(n43), .C(n881), .Y(n918) );
  XNOR3X4 U379 ( .A(n873), .B(n172), .C(n872), .Y(n43) );
  NOR2X1 U380 ( .A(n1131), .B(n1144), .Y(n1133) );
  AND2X2 U381 ( .A(n46), .B(n45), .Y(n1144) );
  NOR2X1 U382 ( .A(n351), .B(n352), .Y(n1131) );
  CLKINVX3 U383 ( .A(B[3]), .Y(n483) );
  XOR2X1 U384 ( .A(n319), .B(n52), .Y(n327) );
  XOR2X1 U385 ( .A(n320), .B(n321), .Y(n52) );
  XOR2X2 U386 ( .A(n322), .B(n102), .Y(n320) );
  AOI21X1 U387 ( .A0(n1148), .A1(n1150), .B0(n53), .Y(n74) );
  INVX1 U388 ( .A(n1149), .Y(n53) );
  NAND2X1 U389 ( .A(n316), .B(n315), .Y(n1149) );
  OR2X2 U390 ( .A(n316), .B(n315), .Y(n1150) );
  NOR2BX1 U391 ( .AN(n314), .B(n75), .Y(n1148) );
  XOR2X2 U392 ( .A(B[8]), .B(B[9]), .Y(n87) );
  NAND2X1 U393 ( .A(n54), .B(n1145), .Y(n355) );
  XNOR2X1 U394 ( .A(n1146), .B(n1134), .Y(n1429) );
  OAI22X1 U395 ( .A0(n627), .A1(n1203), .B0(n1204), .B1(n55), .Y(n632) );
  OAI21X1 U396 ( .A0(n1203), .A1(n55), .B0(n60), .Y(n59) );
  XOR2X1 U397 ( .A(n1041), .B(n56), .Y(n55) );
  NAND2X1 U398 ( .A(n59), .B(n595), .Y(n57) );
  OAI21XL U399 ( .A0(n59), .A1(n595), .B0(n594), .Y(n58) );
  OAI21XL U400 ( .A0(n738), .A1(n63), .B0(n737), .Y(n62) );
  XOR3X2 U401 ( .A(n738), .B(n63), .C(n737), .Y(n770) );
  INVX1 U402 ( .A(n1203), .Y(n65) );
  XNOR3X2 U403 ( .A(n709), .B(n137), .C(n708), .Y(n68) );
  OAI22X1 U404 ( .A0(n794), .A1(n1203), .B0(n1052), .B1(n70), .Y(n799) );
  OAI22X1 U405 ( .A0(n734), .A1(n1052), .B0(n1203), .B1(n70), .Y(n763) );
  XOR2X1 U406 ( .A(n1041), .B(n71), .Y(n70) );
  XNOR3X4 U407 ( .A(n837), .B(n836), .C(n835), .Y(n172) );
  INVX1 U408 ( .A(n1148), .Y(n1153) );
  OAI21X2 U409 ( .A0(n78), .A1(n1147), .B0(n74), .Y(n1134) );
  INVXL U410 ( .A(n313), .Y(n75) );
  NOR2X1 U411 ( .A(n77), .B(n76), .Y(n1147) );
  OAI21XL U412 ( .A0(n1297), .A1(n1303), .B0(n1298), .Y(n76) );
  NAND2X1 U413 ( .A(n282), .B(n281), .Y(n1298) );
  AND2X2 U414 ( .A(n283), .B(n1296), .Y(n77) );
  NAND2X1 U415 ( .A(n1150), .B(n1154), .Y(n78) );
  XOR2X2 U416 ( .A(B[11]), .B(B[10]), .Y(n133) );
  XNOR2X1 U417 ( .A(n498), .B(n499), .Y(n83) );
  XOR2X1 U418 ( .A(n238), .B(n192), .Y(n123) );
  XOR2X1 U419 ( .A(n238), .B(A[24]), .Y(n211) );
  XOR2X1 U420 ( .A(n238), .B(n1036), .Y(n332) );
  XOR2X1 U421 ( .A(n238), .B(n975), .Y(n318) );
  XOR2X1 U422 ( .A(n238), .B(A[4]), .Y(n287) );
  XOR2X1 U423 ( .A(n238), .B(n1239), .Y(n569) );
  XOR2X1 U424 ( .A(n238), .B(A[25]), .Y(n436) );
  XOR2X1 U425 ( .A(n238), .B(n984), .Y(n1062) );
  XOR2X1 U426 ( .A(n85), .B(n966), .Y(n1008) );
  OAI22X1 U427 ( .A0(n1263), .A1(n929), .B0(n931), .B1(n930), .Y(n85) );
  XNOR2X2 U428 ( .A(B[14]), .B(B[13]), .Y(n372) );
  NAND2X4 U429 ( .A(n87), .B(n284), .Y(n1080) );
  XNOR2X4 U430 ( .A(B[8]), .B(B[7]), .Y(n284) );
  OAI2BB1X1 U431 ( .A0N(n89), .A1N(n945), .B0(n88), .Y(n940) );
  NAND2BXL U432 ( .AN(n946), .B(n91), .Y(n89) );
  XOR2X1 U433 ( .A(n946), .B(n91), .Y(n90) );
  AOI2BB1X2 U434 ( .A0N(n935), .A1N(n1080), .B0(n92), .Y(n91) );
  NOR2X1 U435 ( .A(n120), .B(n1078), .Y(n92) );
  OAI2BB1X2 U436 ( .A0N(n94), .A1N(n991), .B0(n93), .Y(n959) );
  NAND2X1 U437 ( .A(n993), .B(n992), .Y(n93) );
  OR2X2 U438 ( .A(n992), .B(n993), .Y(n94) );
  NAND2X1 U439 ( .A(n95), .B(n1189), .Y(n1190) );
  INVX1 U440 ( .A(n1142), .Y(n96) );
  OAI2BB2X2 U441 ( .B0(n99), .B1(n98), .A0N(n1075), .A1N(n97), .Y(n1070) );
  NAND2BX1 U442 ( .AN(n1076), .B(n99), .Y(n97) );
  INVX1 U443 ( .A(n1076), .Y(n98) );
  INVX1 U444 ( .A(n100), .Y(n99) );
  OAI21X1 U445 ( .A0(n1080), .A1(n1077), .B0(n101), .Y(n100) );
  AND2X2 U446 ( .A(n322), .B(n102), .Y(n340) );
  OAI22X1 U447 ( .A0(n231), .A1(n103), .B0(n1055), .B1(n138), .Y(n753) );
  XOR2X1 U448 ( .A(n1037), .B(n894), .Y(n105) );
  INVX1 U449 ( .A(n1055), .Y(n106) );
  XOR2X2 U450 ( .A(n162), .B(n107), .Y(n339) );
  NAND2X1 U451 ( .A(n109), .B(n108), .Y(n107) );
  OR2X2 U452 ( .A(n1080), .B(n324), .Y(n109) );
  OAI2BB1X1 U453 ( .A0N(n113), .A1N(n325), .B0(n110), .Y(n338) );
  NAND2X1 U454 ( .A(n111), .B(n326), .Y(n110) );
  NAND2BX1 U455 ( .AN(n325), .B(n112), .Y(n111) );
  OAI2BB1X1 U456 ( .A0N(n115), .A1N(n572), .B0(n114), .Y(n559) );
  INVX1 U457 ( .A(n118), .Y(n116) );
  OAI22X1 U458 ( .A0(n231), .A1(n543), .B0(n1055), .B1(n521), .Y(n118) );
  NAND2BX1 U459 ( .AN(n888), .B(n10), .Y(n119) );
  XOR2X1 U460 ( .A(n1013), .B(n121), .Y(n120) );
  OAI22X1 U461 ( .A0(n211), .A1(n236), .B0(n122), .B1(n1063), .Y(n526) );
  OAI2BB1X1 U462 ( .A0N(n123), .A1N(n16), .B0(n195), .Y(n552) );
  NAND2X1 U463 ( .A(n995), .B(n994), .Y(mult_x_1_n282) );
  OAI21XL U464 ( .A0(n701), .A1(n127), .B0(n700), .Y(n124) );
  OAI21X2 U465 ( .A0(n1203), .A1(n697), .B0(n128), .Y(n127) );
  OAI21XL U466 ( .A0(n341), .A1(n161), .B0(n129), .Y(n162) );
  OAI21XL U467 ( .A0(n1052), .A1(n13), .B0(n341), .Y(n129) );
  INVXL U468 ( .A(n161), .Y(n130) );
  XNOR3X2 U469 ( .A(n683), .B(n682), .C(n132), .Y(n711) );
  NAND2X2 U470 ( .A(n336), .B(n133), .Y(n335) );
  NAND2X1 U471 ( .A(n710), .B(n709), .Y(n134) );
  OAI22X1 U472 ( .A0(n231), .A1(n138), .B0(n1055), .B1(n687), .Y(n727) );
  XOR2X1 U473 ( .A(n1037), .B(n139), .Y(n138) );
  NAND2X4 U474 ( .A(n142), .B(n227), .Y(n231) );
  OAI21X4 U475 ( .A0(n951), .A1(n952), .B0(n950), .Y(n143) );
  INVX1 U476 ( .A(n952), .Y(n144) );
  INVX1 U477 ( .A(n951), .Y(n145) );
  XOR3X2 U478 ( .A(n952), .B(n950), .C(n951), .Y(n958) );
  NAND2X1 U479 ( .A(n147), .B(n146), .Y(n1167) );
  NAND2X1 U480 ( .A(n772), .B(n774), .Y(n146) );
  OAI21XL U481 ( .A0(n774), .A1(n772), .B0(n773), .Y(n147) );
  XOR3X2 U482 ( .A(n774), .B(n772), .C(n773), .Y(n1169) );
  CLKINVX3 U483 ( .A(B[15]), .Y(n930) );
  XOR3X2 U484 ( .A(n753), .B(n152), .C(n752), .Y(n767) );
  OAI22X2 U485 ( .A0(n750), .A1(n1262), .B0(n724), .B1(n1263), .Y(n152) );
  NAND2XL U486 ( .A(n753), .B(n152), .Y(n149) );
  INVXL U487 ( .A(n152), .Y(n151) );
  OAI2BB1X1 U488 ( .A0N(n155), .A1N(n1083), .B0(n154), .Y(n1089) );
  NAND2XL U489 ( .A(n1084), .B(n158), .Y(n154) );
  NAND2BX1 U490 ( .AN(n1084), .B(n156), .Y(n155) );
  XOR2X1 U491 ( .A(n1083), .B(n157), .Y(n1119) );
  XOR2X1 U492 ( .A(n1084), .B(n158), .Y(n157) );
  NOR2X1 U493 ( .A(n1243), .B(n13), .Y(n158) );
  NAND2BX1 U494 ( .AN(n341), .B(n161), .Y(n160) );
  OAI21XL U495 ( .A0(n165), .A1(n164), .B0(n163), .Y(n516) );
  OAI21XL U496 ( .A0(n519), .A1(n520), .B0(n518), .Y(n163) );
  INVXL U497 ( .A(n520), .Y(n164) );
  XOR2X1 U498 ( .A(n518), .B(n520), .Y(n166) );
  NAND2BX1 U499 ( .AN(n593), .B(n193), .Y(n196) );
  CLKINVX3 U500 ( .A(n1063), .Y(n193) );
  AOI21X1 U501 ( .A0(n613), .A1(n219), .B0(n218), .Y(n217) );
  AOI21X1 U502 ( .A0(n877), .A1(n224), .B0(n223), .Y(n167) );
  NOR2X1 U503 ( .A(n1394), .B(n1392), .Y(n224) );
  OAI21X4 U504 ( .A0(n1399), .A1(n1396), .B0(n1397), .Y(n877) );
  OAI21X2 U505 ( .A0(n1400), .A1(n1407), .B0(n1401), .Y(n168) );
  NOR2X2 U506 ( .A(n1400), .B(n1402), .Y(n169) );
  NAND2X1 U507 ( .A(n872), .B(n873), .Y(n170) );
  NOR2X1 U508 ( .A(n872), .B(n873), .Y(n171) );
  INVX4 U509 ( .A(B[11]), .Y(n373) );
  NOR2X1 U510 ( .A(n650), .B(n1382), .Y(n357) );
  NOR2X1 U511 ( .A(n1413), .B(n1412), .Y(n654) );
  NOR2X1 U512 ( .A(n1259), .B(n733), .Y(n755) );
  XNOR2X1 U513 ( .A(n884), .B(n975), .Y(n733) );
  INVXL U514 ( .A(n8), .Y(n174) );
  INVXL U515 ( .A(n8), .Y(n175) );
  INVXL U516 ( .A(n8), .Y(n176) );
  INVXL U517 ( .A(n8), .Y(n177) );
  XNOR2X2 U518 ( .A(B[12]), .B(B[11]), .Y(n365) );
  BUFX3 U519 ( .A(n336), .Y(n1052) );
  XOR2XL U520 ( .A(B[2]), .B(B[3]), .Y(n230) );
  INVXL U521 ( .A(n1344), .Y(n1279) );
  INVXL U522 ( .A(n1339), .Y(n1280) );
  NAND2XL U523 ( .A(n1273), .B(n1275), .Y(n1278) );
  INVXL U524 ( .A(n1366), .Y(n1289) );
  XNOR2XL U525 ( .A(B[1]), .B(A[11]), .Y(n1049) );
  XNOR2XL U526 ( .A(B[1]), .B(n986), .Y(n1048) );
  XNOR2XL U527 ( .A(n1250), .B(A[4]), .Y(n824) );
  XNOR2XL U528 ( .A(n1250), .B(A[3]), .Y(n883) );
  XNOR2X1 U529 ( .A(n1037), .B(A[11]), .Y(n887) );
  XNOR2XL U530 ( .A(n1013), .B(n982), .Y(n888) );
  OAI22XL U531 ( .A0(n988), .A1(n895), .B0(n855), .B1(n968), .Y(n890) );
  NAND2BXL U532 ( .AN(n1176), .B(n884), .Y(n856) );
  XNOR2XL U533 ( .A(n1205), .B(n970), .Y(n1039) );
  XOR2XL U534 ( .A(n1205), .B(n1015), .Y(n183) );
  BUFX3 U535 ( .A(A[7]), .Y(n984) );
  BUFX3 U536 ( .A(A[8]), .Y(n1017) );
  INVXL U537 ( .A(n1338), .Y(n1313) );
  NOR2XL U538 ( .A(n1278), .B(n1372), .Y(n1339) );
  AOI21X1 U539 ( .A0(n506), .A1(n359), .B0(n358), .Y(n1347) );
  NOR2XL U540 ( .A(n1338), .B(n1360), .Y(n1343) );
  INVXL U541 ( .A(n1362), .Y(n1310) );
  INVX4 U542 ( .A(n930), .Y(n1250) );
  XNOR2XL U543 ( .A(n1234), .B(n1239), .Y(n1220) );
  XOR2XL U544 ( .A(n293), .B(n967), .Y(n754) );
  BUFX4 U545 ( .A(n227), .Y(n1055) );
  BUFX4 U546 ( .A(n284), .Y(n1078) );
  XNOR2XL U547 ( .A(B[1]), .B(A[4]), .Y(n261) );
  BUFX3 U548 ( .A(n236), .Y(n194) );
  XNOR2XL U549 ( .A(n12), .B(A[4]), .Y(n234) );
  NAND2XL U550 ( .A(n1339), .B(n1343), .Y(n1346) );
  ADDFX2 U551 ( .A(n329), .B(n328), .CI(n327), .CO(n330), .S(n316) );
  OAI2BB1XL U552 ( .A0N(n1243), .A1N(n11), .B0(n1242), .Y(n1252) );
  XNOR2XL U553 ( .A(n1234), .B(A[23]), .Y(n1235) );
  OAI22XL U554 ( .A0(n789), .A1(n1080), .B0(n1078), .B1(n754), .Y(n205) );
  OAI21XL U555 ( .A0(n796), .A1(n1063), .B0(n198), .Y(n797) );
  AOI21XL U556 ( .A0(n1353), .A1(n1354), .B0(n254), .Y(n1327) );
  INVXL U557 ( .A(n1352), .Y(n254) );
  NAND2XL U558 ( .A(n260), .B(n259), .Y(n1325) );
  NAND2XL U559 ( .A(n269), .B(n268), .Y(n1329) );
  INVXL U560 ( .A(n1371), .Y(n1276) );
  NAND2X1 U561 ( .A(n356), .B(n717), .Y(n221) );
  NOR2XL U562 ( .A(n1366), .B(n1364), .Y(n1307) );
  INVXL U563 ( .A(n1376), .Y(n507) );
  INVXL U564 ( .A(n1308), .Y(n1288) );
  INVXL U565 ( .A(n1314), .Y(n1287) );
  INVXL U566 ( .A(n1368), .Y(n1275) );
  INVXL U567 ( .A(n1390), .Y(n219) );
  OAI21XL U568 ( .A0(n1392), .A1(n1395), .B0(n1393), .Y(n223) );
  NAND2XL U569 ( .A(n615), .B(n179), .Y(n617) );
  INVXL U570 ( .A(n1382), .Y(n618) );
  INVXL U571 ( .A(n1340), .Y(n189) );
  INVXL U572 ( .A(n1372), .Y(n433) );
  XNOR2X1 U573 ( .A(n1037), .B(A[4]), .Y(n345) );
  XNOR2X1 U574 ( .A(n1041), .B(n970), .Y(n1053) );
  XNOR2X1 U575 ( .A(n1250), .B(n927), .Y(n486) );
  XNOR2XL U576 ( .A(n1041), .B(A[18]), .Y(n490) );
  XNOR2XL U577 ( .A(n1205), .B(A[4]), .Y(n898) );
  XNOR2XL U578 ( .A(n1205), .B(A[3]), .Y(n938) );
  XNOR2XL U579 ( .A(n1013), .B(n975), .Y(n1014) );
  XNOR2XL U580 ( .A(n1013), .B(n1036), .Y(n976) );
  XNOR2XL U581 ( .A(n1205), .B(n1176), .Y(n1040) );
  XNOR2XL U582 ( .A(n1041), .B(A[2]), .Y(n1051) );
  NAND2BXL U583 ( .AN(n1176), .B(n1250), .Y(n929) );
  XNOR2X1 U584 ( .A(n1013), .B(A[4]), .Y(n1077) );
  OAI22X1 U585 ( .A0(n1203), .A1(n373), .B0(n1204), .B1(n337), .Y(n1081) );
  NAND2BXL U586 ( .AN(n1176), .B(n1041), .Y(n337) );
  NAND2BX1 U587 ( .AN(n1176), .B(n1013), .Y(n292) );
  XNOR2X1 U588 ( .A(n1041), .B(A[11]), .Y(n734) );
  XNOR2X1 U589 ( .A(n1041), .B(n986), .Y(n697) );
  XNOR2XL U590 ( .A(n12), .B(A[19]), .Y(n735) );
  XNOR2XL U591 ( .A(n12), .B(n1199), .Y(n698) );
  XNOR2XL U592 ( .A(n1234), .B(n894), .Y(n453) );
  XNOR2XL U593 ( .A(n1041), .B(A[19]), .Y(n454) );
  ADDFX2 U594 ( .A(n493), .B(n492), .CI(n491), .CO(n478), .S(n531) );
  INVXL U595 ( .A(n456), .Y(n491) );
  OAI22X1 U596 ( .A0(n11), .A1(n489), .B0(n1243), .B1(n449), .Y(n493) );
  OAI22X1 U597 ( .A0(n436), .A1(n194), .B0(n1063), .B1(n211), .Y(n456) );
  XNOR2X1 U598 ( .A(n1205), .B(A[18]), .Y(n448) );
  XNOR2XL U599 ( .A(n1041), .B(n1199), .Y(n447) );
  NOR2XL U600 ( .A(n1380), .B(n1378), .Y(n505) );
  NAND2XL U601 ( .A(n1308), .B(n1307), .Y(n1293) );
  NAND2XL U602 ( .A(n1284), .B(n1365), .Y(n1285) );
  NAND2XL U603 ( .A(n956), .B(n1397), .Y(n957) );
  XOR2X1 U604 ( .A(n220), .B(n920), .Y(PRODUCT[19]) );
  NAND2XL U605 ( .A(n919), .B(n1395), .Y(n920) );
  OAI22XL U606 ( .A0(n988), .A1(n987), .B0(n969), .B1(n968), .Y(n1011) );
  OAI22XL U607 ( .A0(n11), .A1(n1039), .B0(n1243), .B1(n971), .Y(n1010) );
  OAI22XL U608 ( .A0(n988), .A1(n1048), .B0(n987), .B1(n1175), .Y(n1047) );
  INVXL U609 ( .A(n1205), .Y(n990) );
  XNOR2XL U610 ( .A(n1205), .B(A[23]), .Y(n1206) );
  OAI22XL U611 ( .A0(n231), .A1(n887), .B0(n1055), .B1(n852), .Y(n865) );
  OAI22X1 U612 ( .A0(n859), .A1(n1063), .B0(n194), .B1(n204), .Y(n861) );
  OAI22XL U613 ( .A0(n1063), .A1(n902), .B0(n194), .B1(n859), .Y(n899) );
  OAI22XL U614 ( .A0(n173), .A1(n858), .B0(n257), .B1(n825), .Y(n891) );
  XNOR2XL U615 ( .A(n12), .B(n1239), .Y(n628) );
  XNOR2XL U616 ( .A(n12), .B(A[24]), .Y(n549) );
  INVXL U617 ( .A(n575), .Y(n550) );
  XNOR2XL U618 ( .A(n12), .B(A[23]), .Y(n592) );
  XNOR2X1 U619 ( .A(n1041), .B(A[16]), .Y(n548) );
  XNOR2XL U620 ( .A(n1041), .B(A[17]), .Y(n542) );
  XNOR2X1 U621 ( .A(B[9]), .B(A[18]), .Y(n574) );
  XNOR2X1 U622 ( .A(n1205), .B(n927), .Y(n571) );
  XNOR2X1 U623 ( .A(n1250), .B(n986), .Y(n544) );
  XNOR2XL U624 ( .A(n1037), .B(A[19]), .Y(n579) );
  XNOR2XL U625 ( .A(n1205), .B(n967), .Y(n582) );
  XNOR2XL U626 ( .A(n1205), .B(n986), .Y(n660) );
  XNOR2X1 U627 ( .A(n1037), .B(A[18]), .Y(n658) );
  XNOR2XL U628 ( .A(n1037), .B(A[17]), .Y(n687) );
  XOR2XL U629 ( .A(n1205), .B(n210), .Y(n209) );
  XNOR2XL U630 ( .A(n12), .B(A[18]), .Y(n759) );
  XNOR2XL U631 ( .A(n1205), .B(n1199), .Y(n382) );
  OAI2BB1XL U632 ( .A0N(n1078), .A1N(n729), .B0(n376), .Y(n393) );
  INVXL U633 ( .A(n375), .Y(n376) );
  OAI22XL U634 ( .A0(n1262), .A1(n377), .B0(n1263), .B1(n389), .Y(n398) );
  OAI22XL U635 ( .A0(n11), .A1(n378), .B0(n1243), .B1(n392), .Y(n397) );
  XNOR2XL U636 ( .A(n1041), .B(n1221), .Y(n415) );
  OAI2BB1XL U637 ( .A0N(n227), .A1N(n231), .B0(n370), .Y(n419) );
  INVXL U638 ( .A(n1341), .Y(n1312) );
  NAND2XL U639 ( .A(n1308), .B(n1313), .Y(n1316) );
  INVXL U640 ( .A(n1360), .Y(n1317) );
  AOI21XL U641 ( .A0(n1344), .A1(n1343), .B0(n1342), .Y(n1345) );
  OAI22XL U642 ( .A0(n1262), .A1(n1220), .B0(n1263), .B1(n1235), .Y(n1238) );
  INVXL U643 ( .A(n1254), .Y(n1236) );
  OAI22XL U644 ( .A0(n1262), .A1(n389), .B0(n1263), .B1(n1207), .Y(n1210) );
  INVXL U645 ( .A(n1218), .Y(n1208) );
  OAI22X1 U646 ( .A0(n751), .A1(n11), .B0(n1243), .B1(n181), .Y(n752) );
  OAI22X2 U647 ( .A0(n1262), .A1(n784), .B0(n1263), .B1(n750), .Y(n787) );
  OAI22X1 U648 ( .A0(n1262), .A1(n813), .B0(n1263), .B1(n784), .Y(n816) );
  OAI22XL U649 ( .A0(n11), .A1(n814), .B0(n1243), .B1(n785), .Y(n815) );
  OAI22X1 U650 ( .A0(n796), .A1(n194), .B0(n1063), .B1(n204), .Y(n826) );
  XOR2XL U651 ( .A(n185), .B(n764), .Y(n806) );
  XOR2XL U652 ( .A(n765), .B(n205), .Y(n185) );
  BUFX3 U653 ( .A(n1050), .Y(n988) );
  OAI22XL U654 ( .A0(n173), .A1(n483), .B0(n257), .B1(n258), .Y(n259) );
  NAND2BXL U655 ( .AN(n1176), .B(n12), .Y(n258) );
  OAI22XL U656 ( .A0(n175), .A1(n264), .B0(n1058), .B1(n263), .Y(n274) );
  OAI22XL U657 ( .A0(n1050), .A1(n262), .B0(n261), .B1(n1175), .Y(n275) );
  NOR2BXL U658 ( .AN(n1176), .B(n194), .Y(n276) );
  OAI22XL U659 ( .A0(n177), .A1(n263), .B0(n1058), .B1(n245), .Y(n273) );
  OAI22XL U660 ( .A0(n965), .A1(n247), .B0(n194), .B1(n246), .Y(n272) );
  OAI22XL U661 ( .A0(n176), .A1(n245), .B0(n1058), .B1(n234), .Y(n244) );
  OAI2BB1XL U662 ( .A0N(n1263), .A1N(n1262), .B0(n1261), .Y(n1264) );
  INVXL U663 ( .A(n1260), .Y(n1261) );
  INVXL U664 ( .A(n1266), .Y(n1256) );
  OAI22XL U665 ( .A0(n988), .A1(n1176), .B0(n250), .B1(n1175), .Y(n1321) );
  NAND2XL U666 ( .A(n251), .B(n988), .Y(n1320) );
  NAND2BXL U667 ( .AN(n1176), .B(B[1]), .Y(n251) );
  NAND2XL U668 ( .A(n1321), .B(n1320), .Y(n1322) );
  INVXL U669 ( .A(n1322), .Y(n1354) );
  INVXL U670 ( .A(n1329), .Y(n270) );
  NOR2XL U671 ( .A(n278), .B(n277), .Y(n1333) );
  NAND2XL U672 ( .A(n278), .B(n277), .Y(n1334) );
  NOR2X1 U673 ( .A(n280), .B(n279), .Y(n1302) );
  INVXL U674 ( .A(n1296), .Y(n1305) );
  OAI21XL U675 ( .A0(n1388), .A1(n1391), .B0(n1389), .Y(n717) );
  NOR2X1 U676 ( .A(n1388), .B(n1390), .Y(n777) );
  XNOR2X1 U677 ( .A(n1205), .B(A[16]), .Y(n489) );
  XNOR2XL U678 ( .A(n1037), .B(A[25]), .Y(n369) );
  NAND2XL U679 ( .A(n1307), .B(n1310), .Y(n1338) );
  INVXL U680 ( .A(n1367), .Y(n1281) );
  NAND2XL U681 ( .A(n1308), .B(n1289), .Y(n1283) );
  INVXL U682 ( .A(n1364), .Y(n1284) );
  INVXL U683 ( .A(n1378), .Y(n535) );
  XNOR2X1 U684 ( .A(n1403), .B(n212), .Y(PRODUCT[15]) );
  NAND2X1 U685 ( .A(n213), .B(n1357), .Y(n212) );
  INVX1 U686 ( .A(n1408), .Y(n216) );
  INVXL U687 ( .A(n1399), .Y(n955) );
  INVX1 U688 ( .A(n878), .Y(n191) );
  INVXL U689 ( .A(n716), .Y(n781) );
  NAND2XL U690 ( .A(n179), .B(n612), .Y(n649) );
  NAND2XL U691 ( .A(n179), .B(n1184), .Y(n655) );
  INVXL U692 ( .A(n1384), .Y(n656) );
  INVXL U693 ( .A(n1377), .Y(n469) );
  INVXL U694 ( .A(n1374), .Y(n472) );
  XNOR2XL U695 ( .A(B[1]), .B(n927), .Y(n969) );
  NAND2BXL U696 ( .AN(n1176), .B(n1205), .Y(n989) );
  XNOR2XL U697 ( .A(B[1]), .B(n967), .Y(n987) );
  XNOR2XL U698 ( .A(n1013), .B(n1199), .Y(n488) );
  XNOR2XL U699 ( .A(n1013), .B(n1015), .Y(n847) );
  XNOR2XL U700 ( .A(n12), .B(n894), .Y(n858) );
  XNOR2X1 U701 ( .A(n1041), .B(n1036), .Y(n903) );
  XNOR2XL U702 ( .A(n1041), .B(n967), .Y(n669) );
  XNOR2XL U703 ( .A(n12), .B(n1221), .Y(n670) );
  XNOR2XL U704 ( .A(n1013), .B(A[25]), .Y(n375) );
  INVXL U705 ( .A(n369), .Y(n370) );
  XNOR2XL U706 ( .A(n1234), .B(A[19]), .Y(n377) );
  XNOR2XL U707 ( .A(n1041), .B(A[23]), .Y(n379) );
  XNOR2XL U708 ( .A(n1234), .B(A[18]), .Y(n381) );
  XNOR2XL U709 ( .A(B[1]), .B(n1017), .Y(n294) );
  AOI21XL U710 ( .A0(n1276), .A1(n1275), .B0(n1274), .Y(n1277) );
  INVXL U711 ( .A(n1369), .Y(n1274) );
  AOI21XL U712 ( .A0(n1311), .A1(n1310), .B0(n1309), .Y(n1341) );
  INVXL U713 ( .A(n1363), .Y(n1309) );
  NAND2XL U714 ( .A(n1289), .B(n1367), .Y(n1290) );
  NAND2XL U715 ( .A(n1275), .B(n1369), .Y(n362) );
  NAND2XL U716 ( .A(n1177), .B(n1389), .Y(n1178) );
  NAND2XL U717 ( .A(n433), .B(n1373), .Y(n434) );
  ADDFX2 U718 ( .A(n344), .B(n343), .CI(n342), .CO(n1123), .S(n350) );
  OAI22XL U719 ( .A0(n965), .A1(n318), .B0(n194), .B1(n332), .Y(n343) );
  OAI22XL U720 ( .A0(n231), .A1(n317), .B0(n1055), .B1(n345), .Y(n344) );
  OAI22X1 U721 ( .A0(n231), .A1(n296), .B0(n1055), .B1(n317), .Y(n326) );
  ADDFX2 U722 ( .A(n1093), .B(n1092), .CI(n1091), .CO(n1127), .S(n1122) );
  OAI22XL U723 ( .A0(n174), .A1(n347), .B0(n1058), .B1(n1059), .Y(n1091) );
  OAI22XL U724 ( .A0(n231), .A1(n345), .B0(n1055), .B1(n1056), .Y(n1093) );
  OAI22XL U725 ( .A0(n1203), .A1(n1053), .B0(n1052), .B1(n1051), .Y(n1083) );
  OAI22XL U726 ( .A0(n1063), .A1(n1062), .B0(n194), .B1(n1061), .Y(n1097) );
  OAI22XL U727 ( .A0(n1060), .A1(n1059), .B0(n1058), .B1(n1057), .Y(n1098) );
  OAI22XL U728 ( .A0(n231), .A1(n1056), .B0(n1055), .B1(n1054), .Y(n1099) );
  INVXL U729 ( .A(n1241), .Y(n1242) );
  XNOR2XL U730 ( .A(n1234), .B(n1199), .Y(n389) );
  OAI22XL U731 ( .A0(n1203), .A1(n490), .B0(n1204), .B1(n454), .Y(n494) );
  OAI22XL U732 ( .A0(n231), .A1(n487), .B0(n227), .B1(n452), .Y(n496) );
  ADDFX2 U733 ( .A(n540), .B(n539), .CI(n538), .CO(n519), .S(n561) );
  OAI2BB1XL U734 ( .A0N(n1058), .A1N(n173), .B0(n485), .Y(n538) );
  INVXL U735 ( .A(n484), .Y(n485) );
  OAI22X1 U736 ( .A0(n231), .A1(n852), .B0(n1055), .B1(n812), .Y(n851) );
  OAI22XL U737 ( .A0(n11), .A1(n848), .B0(n1243), .B1(n814), .Y(n849) );
  OAI22XL U738 ( .A0(n1262), .A1(n896), .B0(n1263), .B1(n883), .Y(n907) );
  OAI22XL U739 ( .A0(n231), .A1(n904), .B0(n1055), .B1(n887), .Y(n910) );
  CMPR32X1 U740 ( .A(n949), .B(n948), .C(n947), .CO(n963), .S(n1001) );
  OAI22XL U741 ( .A0(n231), .A1(n944), .B0(n1055), .B1(n904), .Y(n947) );
  OAI22XL U742 ( .A0(n1063), .A1(n964), .B0(n194), .B1(n902), .Y(n949) );
  OAI22XL U743 ( .A0(n1203), .A1(n943), .B0(n1052), .B1(n903), .Y(n948) );
  OAI22X1 U744 ( .A0(n175), .A1(n942), .B0(n1058), .B1(n897), .Y(n946) );
  OAI22X1 U745 ( .A0(n1262), .A1(n937), .B0(n1263), .B1(n936), .Y(n980) );
  OAI22XL U746 ( .A0(n174), .A1(n1016), .B0(n1058), .B1(n978), .Y(n1019) );
  OAI22XL U747 ( .A0(n231), .A1(n1038), .B0(n1055), .B1(n985), .Y(n1044) );
  OAI22XL U748 ( .A0(n1063), .A1(n1018), .B0(n194), .B1(n983), .Y(n1045) );
  OAI22XL U749 ( .A0(n1203), .A1(n1051), .B0(n1052), .B1(n1042), .Y(n1072) );
  OAI22XL U750 ( .A0(n231), .A1(n985), .B0(n1055), .B1(n944), .Y(n1004) );
  OAI22XL U751 ( .A0(n174), .A1(n978), .B0(n1058), .B1(n942), .Y(n1006) );
  OAI22XL U752 ( .A0(n1203), .A1(n977), .B0(n1052), .B1(n943), .Y(n1005) );
  OAI22XL U753 ( .A0(n965), .A1(n983), .B0(n194), .B1(n964), .Y(n1009) );
  CMPR32X1 U754 ( .A(n1121), .B(n6), .C(n1119), .CO(n1100), .S(n1137) );
  OAI22XL U755 ( .A0(n1080), .A1(n1079), .B0(n1078), .B1(n1077), .Y(n1121) );
  OAI22XL U756 ( .A0(n1063), .A1(n332), .B0(n194), .B1(n1062), .Y(n1096) );
  OAI22XL U757 ( .A0(n1080), .A1(n333), .B0(n1078), .B1(n1079), .Y(n1095) );
  XNOR2X1 U758 ( .A(n1205), .B(n894), .Y(n537) );
  INVX1 U759 ( .A(A[23]), .Y(n192) );
  XNOR2XL U760 ( .A(n1013), .B(A[16]), .Y(n664) );
  OAI22XL U761 ( .A0(n988), .A1(n667), .B0(n599), .B1(n1175), .Y(n666) );
  XNOR2XL U762 ( .A(n1013), .B(n894), .Y(n692) );
  XNOR2XL U763 ( .A(n1013), .B(n927), .Y(n728) );
  OAI22XL U764 ( .A0(n988), .A1(n732), .B0(n695), .B1(n968), .Y(n731) );
  ADDFX2 U765 ( .A(n674), .B(n673), .CI(n672), .CO(n683), .S(n709) );
  OAI22X1 U766 ( .A0(n177), .A1(n670), .B0(n257), .B1(n628), .Y(n673) );
  OAI21XL U767 ( .A0(n629), .A1(n194), .B0(n202), .Y(n672) );
  XNOR2XL U768 ( .A(B[1]), .B(A[19]), .Y(n792) );
  XNOR2XL U769 ( .A(B[1]), .B(n1221), .Y(n732) );
  OAI22X1 U770 ( .A0(n173), .A1(n698), .B0(n1058), .B1(n670), .Y(n701) );
  OAI21XL U771 ( .A0(n671), .A1(n194), .B0(n201), .Y(n700) );
  XNOR2X1 U772 ( .A(n1205), .B(n982), .Y(n751) );
  XNOR2XL U773 ( .A(n1037), .B(n927), .Y(n783) );
  XNOR2X1 U774 ( .A(n1250), .B(n1036), .Y(n784) );
  XNOR2X1 U775 ( .A(n1250), .B(n975), .Y(n813) );
  XNOR2XL U776 ( .A(n1037), .B(n967), .Y(n812) );
  XNOR2XL U777 ( .A(n12), .B(A[16]), .Y(n825) );
  XNOR2X1 U778 ( .A(n1041), .B(n982), .Y(n794) );
  XNOR2XL U779 ( .A(n12), .B(A[17]), .Y(n795) );
  ADDFX2 U780 ( .A(n763), .B(n762), .CI(n761), .CO(n771), .S(n807) );
  OAI22X1 U781 ( .A0(n173), .A1(n759), .B0(n1058), .B1(n735), .Y(n762) );
  OAI21XL U782 ( .A0(n736), .A1(n194), .B0(n199), .Y(n761) );
  OAI22X1 U783 ( .A0(n177), .A1(n735), .B0(n257), .B1(n698), .Y(n738) );
  OAI21XL U784 ( .A0(n699), .A1(n194), .B0(n200), .Y(n737) );
  OAI22XL U785 ( .A0(n729), .A1(n481), .B0(n1078), .B1(n446), .Y(n458) );
  OAI22XL U786 ( .A0(n1203), .A1(n454), .B0(n1204), .B1(n447), .Y(n480) );
  OAI22XL U787 ( .A0(n11), .A1(n449), .B0(n1243), .B1(n448), .Y(n479) );
  ADDFX2 U788 ( .A(n457), .B(n456), .CI(n455), .CO(n477), .S(n513) );
  INVXL U789 ( .A(n436), .Y(n437) );
  XNOR2XL U790 ( .A(n1041), .B(n1239), .Y(n410) );
  ADDFX2 U791 ( .A(n385), .B(n384), .CI(n383), .CO(n401), .S(n426) );
  OAI22XL U792 ( .A0(n1203), .A1(n410), .B0(n1204), .B1(n379), .Y(n384) );
  INVXL U793 ( .A(n394), .Y(n383) );
  OAI22XL U794 ( .A0(n1262), .A1(n381), .B0(n1263), .B1(n377), .Y(n385) );
  ADDFX2 U795 ( .A(n418), .B(n417), .CI(n416), .CO(n427), .S(n463) );
  OAI22XL U796 ( .A0(n11), .A1(n411), .B0(n1243), .B1(n382), .Y(n416) );
  OAI22XL U797 ( .A0(n1262), .A1(n414), .B0(n1263), .B1(n381), .Y(n417) );
  OAI22XL U798 ( .A0(n729), .A1(n412), .B0(n1078), .B1(n380), .Y(n418) );
  XNOR2XL U799 ( .A(B[1]), .B(A[2]), .Y(n255) );
  XNOR2XL U800 ( .A(B[1]), .B(A[3]), .Y(n262) );
  XNOR2XL U801 ( .A(n12), .B(A[2]), .Y(n263) );
  XNOR2XL U802 ( .A(n12), .B(A[3]), .Y(n245) );
  NAND2BXL U803 ( .AN(n1176), .B(n1037), .Y(n226) );
  ADDFX2 U804 ( .A(n303), .B(n302), .CI(n301), .CO(n308), .S(n310) );
  OAI22X1 U805 ( .A0(n231), .A1(n232), .B0(n1055), .B1(n297), .Y(n302) );
  OAI22XL U806 ( .A0(n174), .A1(n234), .B0(n1058), .B1(n286), .Y(n303) );
  ADDFX2 U807 ( .A(n300), .B(n299), .CI(n298), .CO(n319), .S(n309) );
  OAI22XL U808 ( .A0(n988), .A1(n295), .B0(n294), .B1(n1175), .Y(n299) );
  NOR2BXL U809 ( .AN(n1176), .B(n1078), .Y(n300) );
  OAI22XL U810 ( .A0(n231), .A1(n297), .B0(n1055), .B1(n296), .Y(n298) );
  NAND2XL U811 ( .A(n1310), .B(n1363), .Y(n1294) );
  OAI22XL U812 ( .A0(n11), .A1(n392), .B0(n1243), .B1(n1206), .Y(n1213) );
  OAI22XL U813 ( .A0(n1262), .A1(n1207), .B0(n1263), .B1(n1220), .Y(n1225) );
  OAI22XL U814 ( .A0(n11), .A1(n1206), .B0(n1243), .B1(n1223), .Y(n1226) );
  OAI2BB1XL U815 ( .A0N(n1204), .A1N(n1203), .B0(n1202), .Y(n1217) );
  INVXL U816 ( .A(n1201), .Y(n1202) );
  ADDFX2 U817 ( .A(n517), .B(n516), .CI(n515), .CO(n510), .S(n564) );
  OAI22XL U818 ( .A0(n177), .A1(n628), .B0(n1058), .B1(n592), .Y(n631) );
  OAI21XL U819 ( .A0(n593), .A1(n194), .B0(n197), .Y(n630) );
  OAI2BB1XL U820 ( .A0N(n1175), .A1N(n988), .B0(n550), .Y(n594) );
  OR2XL U821 ( .A(n578), .B(n577), .Y(n554) );
  OAI22XL U822 ( .A0(n729), .A1(n596), .B0(n1078), .B1(n574), .Y(n588) );
  OAI22XL U823 ( .A0(n11), .A1(n582), .B0(n1243), .B1(n571), .Y(n583) );
  OAI21XL U824 ( .A0(n569), .A1(n194), .B0(n196), .Y(n585) );
  OAI22X1 U825 ( .A0(n1262), .A1(n659), .B0(n1263), .B1(n580), .Y(n662) );
  OAI22X1 U826 ( .A0(n1262), .A1(n688), .B0(n1263), .B1(n659), .Y(n690) );
  OAI22X1 U827 ( .A0(n231), .A1(n687), .B0(n1055), .B1(n658), .Y(n691) );
  OAI22X1 U828 ( .A0(n660), .A1(n1243), .B0(n11), .B1(n209), .Y(n689) );
  OAI22X2 U829 ( .A0(n1262), .A1(n724), .B0(n1263), .B1(n688), .Y(n726) );
  OAI21XL U830 ( .A0(n209), .A1(n1243), .B0(n182), .Y(n725) );
  OAI22XL U831 ( .A0(n11), .A1(n382), .B0(n1243), .B1(n378), .Y(n388) );
  CMPR32X1 U832 ( .A(n427), .B(n426), .C(n425), .CO(n428), .S(n464) );
  NOR2BXL U833 ( .AN(n1176), .B(n1058), .Y(n252) );
  OAI22XL U834 ( .A0(n988), .A1(n250), .B0(n255), .B1(n1175), .Y(n253) );
  NAND2XL U835 ( .A(n1317), .B(n1361), .Y(n1318) );
  INVXL U836 ( .A(n1348), .Y(n1349) );
  OR2XL U837 ( .A(n1340), .B(n1346), .Y(n225) );
  OAI22XL U838 ( .A0(n1262), .A1(n1235), .B0(n1263), .B1(n1251), .Y(n1248) );
  ADDFX2 U839 ( .A(n1216), .B(n1215), .CI(n1214), .CO(n1228), .S(n1229) );
  OAI2BB1X1 U840 ( .A0N(n916), .A1N(n915), .B0(n203), .Y(n881) );
  OAI21XL U841 ( .A0(n915), .A1(n916), .B0(n914), .Y(n203) );
  INVXL U842 ( .A(mult_x_1_n306), .Y(n1115) );
  ADDFX2 U843 ( .A(n641), .B(n640), .CI(n639), .CO(n642), .S(n684) );
  ADDFX2 U844 ( .A(n638), .B(n637), .CI(n636), .CO(n645), .S(n685) );
  NAND2XL U845 ( .A(n765), .B(n205), .Y(n206) );
  NAND2XL U846 ( .A(n764), .B(n208), .Y(n207) );
  NAND2X1 U847 ( .A(n836), .B(n837), .Y(n187) );
  NAND2XL U848 ( .A(n253), .B(n252), .Y(n1352) );
  OAI21XL U849 ( .A0(n1192), .A1(n1191), .B0(n1190), .Y(mult_x_1_n309) );
  NOR2XL U850 ( .A(n1230), .B(n1229), .Y(mult_x_1_n136) );
  NAND2XL U851 ( .A(n1150), .B(n1149), .Y(n1151) );
  NAND2XL U852 ( .A(n1270), .B(n1269), .Y(mult_x_1_n58) );
  NAND2XL U853 ( .A(n1268), .B(n1267), .Y(n1269) );
  NOR2XL U854 ( .A(n1272), .B(n1271), .Y(mult_x_1_n109) );
  NAND2XL U855 ( .A(n1272), .B(n1271), .Y(mult_x_1_n110) );
  NOR2XL U856 ( .A(n1245), .B(n1244), .Y(mult_x_1_n120) );
  NAND2XL U857 ( .A(n1245), .B(n1244), .Y(mult_x_1_n121) );
  NOR2XL U858 ( .A(n1228), .B(n1227), .Y(mult_x_1_n129) );
  NAND2XL U859 ( .A(n1228), .B(n1227), .Y(mult_x_1_n130) );
  NAND2XL U860 ( .A(n1230), .B(n1229), .Y(mult_x_1_n137) );
  NOR2XL U861 ( .A(n842), .B(n841), .Y(mult_x_1_n262) );
  NOR2BXL U862 ( .AN(n1176), .B(n1175), .Y(n1439) );
  XNOR2XL U863 ( .A(n1355), .B(n1354), .Y(n1437) );
  NAND2XL U864 ( .A(n1353), .B(n1352), .Y(n1355) );
  NAND2XL U865 ( .A(n1326), .B(n1325), .Y(n1328) );
  INVXL U866 ( .A(n1324), .Y(n1326) );
  NAND2XL U867 ( .A(n1330), .B(n1329), .Y(n1332) );
  NAND2XL U868 ( .A(n1335), .B(n1334), .Y(n1337) );
  INVXL U869 ( .A(n1333), .Y(n1335) );
  NAND2XL U870 ( .A(n1304), .B(n1303), .Y(n1306) );
  INVXL U871 ( .A(n1302), .Y(n1304) );
  NAND2XL U872 ( .A(n1299), .B(n1298), .Y(n1300) );
  BUFX4 U873 ( .A(B[16]), .Y(n884) );
  INVX8 U874 ( .A(n368), .Y(n1037) );
  XOR2X1 U875 ( .A(n186), .B(n957), .Y(PRODUCT[18]) );
  AOI2BB1X2 U876 ( .A0N(n876), .A1N(n1398), .B0(n955), .Y(n186) );
  CMPR22X1 U877 ( .A(n694), .B(n693), .CO(n675), .S(n703) );
  CMPR22X1 U878 ( .A(n854), .B(n853), .CO(n829), .S(n864) );
  OAI22X1 U879 ( .A0(n1050), .A1(n294), .B0(n323), .B1(n1175), .Y(n322) );
  CMPR22X1 U880 ( .A(n756), .B(n755), .CO(n739), .S(n765) );
  CMPR22X1 U881 ( .A(n249), .B(n248), .CO(n243), .S(n271) );
  OAI22X1 U882 ( .A0(n1063), .A1(n238), .B0(n194), .B1(n237), .Y(n248) );
  CMPR22X1 U883 ( .A(n598), .B(n597), .CO(n587), .S(n634) );
  CMPR22X1 U884 ( .A(n290), .B(n289), .CO(n304), .S(n312) );
  OAI22X1 U885 ( .A0(n231), .A1(n368), .B0(n1055), .B1(n226), .Y(n289) );
  OAI22X1 U886 ( .A0(n729), .A1(n380), .B0(n1078), .B1(n375), .Y(n394) );
  CMPR22X1 U887 ( .A(n266), .B(n265), .CO(n268), .S(n260) );
  OAI22X1 U888 ( .A0(n176), .A1(n256), .B0(n1058), .B1(n264), .Y(n265) );
  OR2X2 U889 ( .A(n765), .B(n205), .Y(n208) );
  OAI21XL U890 ( .A0(n1347), .A1(n1280), .B0(n1279), .Y(n180) );
  AOI21XL U891 ( .A0(n180), .A1(n1289), .B0(n1281), .Y(n1282) );
  XOR2X1 U892 ( .A(n217), .B(n1178), .Y(PRODUCT[22]) );
  XNOR2XL U893 ( .A(n884), .B(n1221), .Y(n1222) );
  XNOR2XL U894 ( .A(n1234), .B(n1221), .Y(n1207) );
  XNOR2X1 U895 ( .A(n1037), .B(n1221), .Y(n521) );
  CMPR22X1 U896 ( .A(n791), .B(n790), .CO(n764), .S(n801) );
  NOR2XL U897 ( .A(n776), .B(n775), .Y(mult_x_1_n244) );
  NAND2X1 U898 ( .A(n224), .B(n878), .Y(n190) );
  XOR2X1 U899 ( .A(n876), .B(n997), .Y(PRODUCT[17]) );
  XOR3X2 U900 ( .A(n916), .B(n914), .C(n915), .Y(n921) );
  XOR2X1 U901 ( .A(n216), .B(n1404), .Y(PRODUCT[14]) );
  XNOR2X1 U902 ( .A(n884), .B(n986), .Y(n482) );
  OAI22X1 U903 ( .A0(n1203), .A1(n1042), .B0(n1052), .B1(n977), .Y(n1020) );
  NOR2X1 U904 ( .A(n1259), .B(n522), .Y(n573) );
  OAI21XL U905 ( .A0(n1182), .A1(n720), .B0(n719), .Y(n723) );
  OAI21XL U906 ( .A0(n1386), .A1(n780), .B0(n1387), .Y(n222) );
  CMPR22X1 U907 ( .A(n820), .B(n819), .CO(n800), .S(n830) );
  ADDFHX4 U908 ( .A(n963), .B(n962), .CI(n961), .CO(n951), .S(n1000) );
  NAND2X1 U909 ( .A(n1412), .B(n1413), .Y(n1183) );
  ADDFHX1 U910 ( .A(n1024), .B(n1023), .CI(n1022), .CO(n999), .S(n1030) );
  NAND2X1 U911 ( .A(n364), .B(n365), .Y(n581) );
  XNOR2X2 U912 ( .A(B[2]), .B(B[1]), .Y(n257) );
  XNOR2X1 U913 ( .A(n1250), .B(n970), .Y(n936) );
  XNOR2X1 U914 ( .A(n1013), .B(A[2]), .Y(n333) );
  XNOR2XL U915 ( .A(B[1]), .B(A[23]), .Y(n667) );
  XNOR2XL U916 ( .A(n1234), .B(A[17]), .Y(n414) );
  OAI22X1 U917 ( .A0(n1063), .A1(n246), .B0(n194), .B1(n233), .Y(n239) );
  OAI22X1 U918 ( .A0(n231), .A1(n1054), .B0(n1055), .B1(n1038), .Y(n1074) );
  INVX1 U919 ( .A(B[0]), .Y(n968) );
  XNOR2X1 U920 ( .A(B[1]), .B(n1036), .Y(n228) );
  XNOR2X1 U921 ( .A(B[1]), .B(n984), .Y(n295) );
  BUFX3 U922 ( .A(n968), .Y(n1175) );
  OAI22X1 U923 ( .A0(n988), .A1(n228), .B0(n295), .B1(n1175), .Y(n290) );
  BUFX3 U924 ( .A(A[0]), .Y(n1176) );
  NOR2BX1 U925 ( .AN(n1176), .B(n1055), .Y(n241) );
  XNOR2X1 U926 ( .A(B[1]), .B(n975), .Y(n235) );
  XOR2X1 U927 ( .A(B[4]), .B(B[5]), .Y(n229) );
  XNOR2X1 U928 ( .A(B[4]), .B(B[3]), .Y(n236) );
  NAND2X2 U929 ( .A(n229), .B(n236), .Y(n965) );
  BUFX3 U930 ( .A(n257), .Y(n1058) );
  XNOR2X1 U931 ( .A(n12), .B(n975), .Y(n286) );
  XNOR2X1 U932 ( .A(n1037), .B(n970), .Y(n297) );
  OAI22XL U933 ( .A0(n1063), .A1(n233), .B0(n194), .B1(n288), .Y(n301) );
  OAI22X1 U934 ( .A0(n988), .A1(n261), .B0(n235), .B1(n1175), .Y(n249) );
  CMPR32X1 U935 ( .A(n244), .B(n243), .C(n242), .CO(n281), .S(n280) );
  XNOR2X1 U936 ( .A(B[1]), .B(n970), .Y(n250) );
  OR2X2 U937 ( .A(n253), .B(n252), .Y(n1353) );
  OAI22X1 U938 ( .A0(n988), .A1(n255), .B0(n262), .B1(n1175), .Y(n266) );
  XNOR2X1 U939 ( .A(n12), .B(n1176), .Y(n256) );
  XNOR2XL U940 ( .A(n12), .B(n970), .Y(n264) );
  NOR2XL U941 ( .A(n260), .B(n259), .Y(n1324) );
  OAI21XL U942 ( .A0(n1327), .A1(n1324), .B0(n1325), .Y(n1331) );
  NOR2XL U943 ( .A(n269), .B(n268), .Y(n267) );
  INVXL U944 ( .A(n267), .Y(n1330) );
  AOI21XL U945 ( .A0(n1331), .A1(n1330), .B0(n270), .Y(n1336) );
  CMPR32X1 U946 ( .A(n273), .B(n272), .C(n271), .CO(n279), .S(n278) );
  CMPR32X1 U947 ( .A(n276), .B(n275), .C(n274), .CO(n277), .S(n269) );
  OAI21XL U948 ( .A0(n1336), .A1(n1333), .B0(n1334), .Y(n1296) );
  XNOR2X1 U949 ( .A(n1037), .B(A[2]), .Y(n296) );
  XNOR2X1 U950 ( .A(n1037), .B(A[3]), .Y(n317) );
  INVX4 U951 ( .A(B[9]), .Y(n293) );
  XNOR2X1 U952 ( .A(n1013), .B(n970), .Y(n324) );
  XNOR2X1 U953 ( .A(n12), .B(n1036), .Y(n291) );
  OAI22X1 U954 ( .A0(n176), .A1(n286), .B0(n1058), .B1(n291), .Y(n306) );
  OAI22X2 U955 ( .A0(n1063), .A1(n288), .B0(n194), .B1(n287), .Y(n305) );
  XNOR2X1 U956 ( .A(B[1]), .B(n982), .Y(n323) );
  BUFX4 U957 ( .A(n1080), .Y(n729) );
  CMPR32X1 U958 ( .A(n309), .B(n308), .C(n307), .CO(n315), .S(n314) );
  CMPR32X1 U959 ( .A(n312), .B(n311), .C(n310), .CO(n313), .S(n282) );
  OR2X2 U960 ( .A(n314), .B(n313), .Y(n1154) );
  XNOR2X1 U961 ( .A(n12), .B(n1017), .Y(n347) );
  XNOR2X1 U962 ( .A(B[1]), .B(n1015), .Y(n334) );
  OAI22XL U963 ( .A0(n988), .A1(n334), .B0(n1049), .B1(n1175), .Y(n1082) );
  BUFX3 U964 ( .A(n336), .Y(n1204) );
  INVX8 U965 ( .A(n373), .Y(n1041) );
  XNOR2X1 U966 ( .A(n1037), .B(n975), .Y(n1056) );
  XNOR2X1 U967 ( .A(n1041), .B(n1176), .Y(n346) );
  OAI22X1 U968 ( .A0(n1203), .A1(n346), .B0(n1052), .B1(n1053), .Y(n1092) );
  XNOR2X1 U969 ( .A(n12), .B(n982), .Y(n1059) );
  CMPR32X1 U970 ( .A(n350), .B(n349), .C(n348), .CO(n352), .S(n331) );
  INVXL U971 ( .A(n1131), .Y(n353) );
  NAND2XL U972 ( .A(n353), .B(n1130), .Y(n354) );
  XNOR2X1 U973 ( .A(n355), .B(n354), .Y(n1428) );
  NOR2X1 U974 ( .A(n1414), .B(n1415), .Y(n716) );
  NAND2X1 U975 ( .A(n1414), .B(n1415), .Y(n780) );
  NOR2XL U976 ( .A(n1376), .B(n1374), .Y(n359) );
  NAND2XL U977 ( .A(n505), .B(n359), .Y(n1340) );
  NOR2XL U978 ( .A(n1340), .B(n1372), .Y(n404) );
  NAND2XL U979 ( .A(n404), .B(n1273), .Y(n361) );
  OAI21XL U980 ( .A0(n1374), .A1(n1377), .B0(n1375), .Y(n358) );
  OAI21XL U981 ( .A0(n1347), .A1(n1372), .B0(n1373), .Y(n405) );
  AOI21XL U982 ( .A0(n405), .A1(n1273), .B0(n1276), .Y(n360) );
  OAI21XL U983 ( .A0(n1350), .A1(n361), .B0(n360), .Y(n363) );
  XOR2X1 U984 ( .A(B[12]), .B(B[13]), .Y(n364) );
  XNOR2X1 U985 ( .A(n1205), .B(n1221), .Y(n378) );
  XNOR2X1 U986 ( .A(B[16]), .B(B[15]), .Y(n450) );
  XNOR2XL U987 ( .A(n1037), .B(A[24]), .Y(n444) );
  OAI22X1 U988 ( .A0(n231), .A1(n444), .B0(n1055), .B1(n369), .Y(n420) );
  XOR2X1 U989 ( .A(B[14]), .B(B[15]), .Y(n371) );
  NAND2X2 U990 ( .A(n372), .B(n371), .Y(n931) );
  XNOR2XL U991 ( .A(n1013), .B(A[24]), .Y(n380) );
  XNOR2X1 U992 ( .A(n1205), .B(n1239), .Y(n392) );
  XNOR2XL U993 ( .A(n1041), .B(A[24]), .Y(n391) );
  OAI22XL U994 ( .A0(n1203), .A1(n379), .B0(n1204), .B1(n391), .Y(n396) );
  XNOR2XL U995 ( .A(n1013), .B(A[23]), .Y(n412) );
  XNOR2X1 U996 ( .A(n1205), .B(A[19]), .Y(n411) );
  CMPR32X1 U997 ( .A(n388), .B(n387), .C(n386), .CO(n430), .S(n425) );
  XNOR2X1 U998 ( .A(n884), .B(A[19]), .Y(n390) );
  XNOR2XL U999 ( .A(n1041), .B(A[25]), .Y(n1201) );
  OAI22X1 U1000 ( .A0(n1203), .A1(n391), .B0(n1204), .B1(n1201), .Y(n1218) );
  CMPR32X1 U1001 ( .A(n395), .B(n394), .C(n393), .CO(n1212), .S(n400) );
  CMPR32X1 U1002 ( .A(n398), .B(n397), .C(n396), .CO(n1211), .S(n399) );
  CMPR32X1 U1003 ( .A(n401), .B(n400), .C(n399), .CO(n1196), .S(n429) );
  NOR2XL U1004 ( .A(n403), .B(n402), .Y(mult_x_1_n151) );
  NAND2XL U1005 ( .A(n403), .B(n402), .Y(mult_x_1_n152) );
  INVXL U1006 ( .A(n404), .Y(n407) );
  OAI22XL U1007 ( .A0(n1203), .A1(n415), .B0(n1204), .B1(n410), .Y(n424) );
  OAI22X1 U1008 ( .A0(n11), .A1(n448), .B0(n1243), .B1(n411), .Y(n443) );
  XNOR2X1 U1009 ( .A(B[9]), .B(n1239), .Y(n446) );
  OAI22X1 U1010 ( .A0(n729), .A1(n446), .B0(n1078), .B1(n412), .Y(n442) );
  XNOR2X1 U1011 ( .A(n884), .B(n894), .Y(n413) );
  OAI22XL U1012 ( .A0(n1262), .A1(n445), .B0(n1263), .B1(n414), .Y(n439) );
  OAI22XL U1013 ( .A0(n1203), .A1(n447), .B0(n1204), .B1(n415), .Y(n438) );
  CMPR32X1 U1014 ( .A(n421), .B(n420), .C(n419), .CO(n386), .S(n462) );
  NOR2XL U1015 ( .A(n432), .B(n431), .Y(mult_x_1_n160) );
  NAND2XL U1016 ( .A(n432), .B(n431), .Y(mult_x_1_n161) );
  XNOR2XL U1017 ( .A(n884), .B(n927), .Y(n435) );
  CMPR32X1 U1018 ( .A(n440), .B(n439), .C(n438), .CO(n422), .S(n476) );
  ADDFHX1 U1019 ( .A(n443), .B(n442), .CI(n441), .CO(n423), .S(n475) );
  XNOR2X1 U1020 ( .A(n1037), .B(A[23]), .Y(n452) );
  OAI22XL U1021 ( .A0(n231), .A1(n452), .B0(n227), .B1(n444), .Y(n460) );
  OAI22XL U1022 ( .A0(n1262), .A1(n453), .B0(n1263), .B1(n445), .Y(n459) );
  XNOR2X1 U1023 ( .A(B[9]), .B(n1221), .Y(n481) );
  XNOR2XL U1024 ( .A(n884), .B(n967), .Y(n451) );
  XNOR2X1 U1025 ( .A(n1037), .B(n1239), .Y(n487) );
  OAI22X1 U1026 ( .A0(n1262), .A1(n486), .B0(n1263), .B1(n453), .Y(n495) );
  CMPR32X1 U1027 ( .A(n460), .B(n459), .C(n458), .CO(n499), .S(n512) );
  ADDFHX1 U1028 ( .A(n463), .B(n462), .CI(n461), .CO(n465), .S(n500) );
  CMPR32X1 U1029 ( .A(n466), .B(n465), .C(n464), .CO(n432), .S(n467) );
  NOR2XL U1030 ( .A(n468), .B(n467), .Y(mult_x_1_n169) );
  NAND2XL U1031 ( .A(n468), .B(n467), .Y(mult_x_1_n170) );
  AOI21XL U1032 ( .A0(n506), .A1(n507), .B0(n469), .Y(n470) );
  NAND2X1 U1033 ( .A(n472), .B(n1375), .Y(n473) );
  CMPR32X1 U1034 ( .A(n477), .B(n476), .C(n475), .CO(n502), .S(n511) );
  CMPR32X1 U1035 ( .A(n480), .B(n479), .C(n478), .CO(n498), .S(n517) );
  NOR2X1 U1036 ( .A(n1259), .B(n482), .Y(n540) );
  XNOR2X1 U1037 ( .A(n12), .B(A[25]), .Y(n484) );
  OAI22X1 U1038 ( .A0(n173), .A1(n549), .B0(n1058), .B1(n484), .Y(n539) );
  XNOR2X1 U1039 ( .A(n1250), .B(n967), .Y(n523) );
  OAI22X2 U1040 ( .A0(n1262), .A1(n523), .B0(n1263), .B1(n486), .Y(n525) );
  OAI22XL U1041 ( .A0(n231), .A1(n521), .B0(n1055), .B1(n487), .Y(n524) );
  XNOR2X1 U1042 ( .A(n1013), .B(A[19]), .Y(n541) );
  OAI22X1 U1043 ( .A0(n729), .A1(n541), .B0(n1078), .B1(n488), .Y(n529) );
  OAI22X1 U1044 ( .A0(n11), .A1(n537), .B0(n1243), .B1(n489), .Y(n528) );
  OAI22XL U1045 ( .A0(n1203), .A1(n542), .B0(n1204), .B1(n490), .Y(n527) );
  CMPR32X1 U1046 ( .A(n502), .B(n501), .C(n500), .CO(n468), .S(n503) );
  NOR2XL U1047 ( .A(n504), .B(n503), .Y(mult_x_1_n176) );
  NAND2XL U1048 ( .A(n504), .B(n503), .Y(mult_x_1_n177) );
  ADDFHX1 U1049 ( .A(n511), .B(n510), .CI(n509), .CO(n504), .S(n534) );
  CMPR32X1 U1050 ( .A(n514), .B(n513), .C(n512), .CO(n497), .S(n565) );
  XNOR2X1 U1051 ( .A(n1037), .B(n1199), .Y(n543) );
  XNOR2XL U1052 ( .A(n884), .B(A[11]), .Y(n522) );
  OAI22XL U1053 ( .A0(n1262), .A1(n544), .B0(n1263), .B1(n523), .Y(n572) );
  CMPR32X1 U1054 ( .A(n532), .B(n531), .C(n530), .CO(n515), .S(n545) );
  NOR2XL U1055 ( .A(n534), .B(n533), .Y(mult_x_1_n183) );
  NAND2X1 U1056 ( .A(n535), .B(n1379), .Y(n536) );
  OAI22X1 U1057 ( .A0(n11), .A1(n571), .B0(n1243), .B1(n537), .Y(n553) );
  OAI22XL U1058 ( .A0(n729), .A1(n574), .B0(n1078), .B1(n541), .Y(n556) );
  OAI22XL U1059 ( .A0(n1203), .A1(n548), .B0(n1204), .B1(n542), .Y(n555) );
  OAI22XL U1060 ( .A0(n231), .A1(n579), .B0(n1055), .B1(n543), .Y(n578) );
  OAI22X1 U1061 ( .A0(n1262), .A1(n580), .B0(n1263), .B1(n544), .Y(n577) );
  XNOR2XL U1062 ( .A(B[1]), .B(A[25]), .Y(n575) );
  ADDFX2 U1063 ( .A(n553), .B(n552), .CI(n551), .CO(n562), .S(n625) );
  CMPR32X1 U1064 ( .A(n556), .B(n555), .C(n554), .CO(n560), .S(n624) );
  CMPR32X1 U1065 ( .A(n559), .B(n558), .C(n557), .CO(n546), .S(n605) );
  CMPR32X1 U1066 ( .A(n562), .B(n561), .C(n560), .CO(n609), .S(n604) );
  ADDFHX1 U1067 ( .A(n565), .B(n564), .CI(n563), .CO(n533), .S(n566) );
  NOR2XL U1068 ( .A(n567), .B(n566), .Y(mult_x_1_n194) );
  NAND2XL U1069 ( .A(n567), .B(n566), .Y(mult_x_1_n195) );
  XNOR2X1 U1070 ( .A(n884), .B(n1015), .Y(n570) );
  NOR2XL U1071 ( .A(n1259), .B(n570), .Y(n584) );
  XNOR2X1 U1072 ( .A(n1013), .B(A[17]), .Y(n596) );
  XNOR2XL U1073 ( .A(B[1]), .B(A[24]), .Y(n599) );
  OAI22X1 U1074 ( .A0(n988), .A1(n599), .B0(n575), .B1(n1175), .Y(n598) );
  XNOR2X1 U1075 ( .A(n884), .B(n982), .Y(n576) );
  NOR2X1 U1076 ( .A(n1259), .B(n576), .Y(n597) );
  OAI22X1 U1077 ( .A0(n231), .A1(n658), .B0(n1055), .B1(n579), .Y(n663) );
  XNOR2X1 U1078 ( .A(n1250), .B(n1015), .Y(n659) );
  OAI22X1 U1079 ( .A0(n11), .A1(n660), .B0(n1243), .B1(n582), .Y(n661) );
  CMPR32X1 U1080 ( .A(n585), .B(n584), .C(n583), .CO(n591), .S(n640) );
  CMPR32X1 U1081 ( .A(n588), .B(n587), .C(n586), .CO(n589), .S(n639) );
  CMPR32X1 U1082 ( .A(n591), .B(n590), .C(n589), .CO(n623), .S(n643) );
  NAND2XL U1083 ( .A(n642), .B(n643), .Y(n603) );
  XNOR2X1 U1084 ( .A(n1041), .B(n927), .Y(n627) );
  OAI22XL U1085 ( .A0(n729), .A1(n664), .B0(n1078), .B1(n596), .Y(n635) );
  XNOR2XL U1086 ( .A(n884), .B(n1017), .Y(n600) );
  NAND2XL U1087 ( .A(n643), .B(n645), .Y(n602) );
  NAND2XL U1088 ( .A(n642), .B(n645), .Y(n601) );
  NAND3X1 U1089 ( .A(n603), .B(n602), .C(n601), .Y(n622) );
  CMPR32X1 U1090 ( .A(n606), .B(n605), .C(n604), .CO(n607), .S(n621) );
  NAND2XL U1091 ( .A(n611), .B(n610), .Y(mult_x_1_n198) );
  OAI21XL U1092 ( .A0(n617), .A1(n1182), .B0(n616), .Y(n620) );
  ADDFHX1 U1093 ( .A(n626), .B(n625), .CI(n624), .CO(n606), .S(n1159) );
  CMPR32X1 U1094 ( .A(n632), .B(n631), .C(n630), .CO(n638), .S(n682) );
  CMPR32X1 U1095 ( .A(n635), .B(n634), .C(n633), .CO(n636), .S(n681) );
  NAND2XL U1096 ( .A(n647), .B(n646), .Y(mult_x_1_n207) );
  AOI21XL U1097 ( .A0(n1179), .A1(n612), .B0(n614), .Y(n648) );
  NAND2X1 U1098 ( .A(n18), .B(n651), .Y(n652) );
  NAND2X1 U1099 ( .A(n656), .B(n1385), .Y(n657) );
  XNOR2X1 U1100 ( .A(n1250), .B(n982), .Y(n688) );
  OAI22XL U1101 ( .A0(n729), .A1(n692), .B0(n1078), .B1(n664), .Y(n677) );
  ADDHXL U1102 ( .A(n666), .B(n665), .CO(n633), .S(n676) );
  XNOR2X1 U1103 ( .A(B[1]), .B(n1239), .Y(n695) );
  OAI22X1 U1104 ( .A0(n988), .A1(n695), .B0(n667), .B1(n1175), .Y(n694) );
  XNOR2XL U1105 ( .A(n884), .B(n984), .Y(n668) );
  CMPR32X1 U1106 ( .A(n677), .B(n675), .C(n676), .CO(n678), .S(n708) );
  CMPR32X1 U1107 ( .A(n680), .B(n679), .C(n678), .CO(n1162), .S(n712) );
  XNOR2X1 U1108 ( .A(n1250), .B(n1017), .Y(n724) );
  OAI22XL U1109 ( .A0(n729), .A1(n728), .B0(n1078), .B1(n692), .Y(n704) );
  XNOR2XL U1110 ( .A(n884), .B(n1036), .Y(n696) );
  CMPR32X1 U1111 ( .A(n704), .B(n703), .C(n702), .CO(n705), .S(n745) );
  CMPR32X1 U1112 ( .A(n707), .B(n706), .C(n705), .CO(n1165), .S(n748) );
  NOR2X1 U1113 ( .A(n715), .B(n714), .Y(mult_x_1_n226) );
  NAND2XL U1114 ( .A(n715), .B(n714), .Y(mult_x_1_n227) );
  NAND2XL U1115 ( .A(n777), .B(n781), .Y(n720) );
  INVXL U1116 ( .A(n780), .Y(n718) );
  AOI21XL U1117 ( .A0(n717), .A1(n781), .B0(n718), .Y(n719) );
  INVXL U1118 ( .A(n1386), .Y(n721) );
  XNOR2X1 U1119 ( .A(n723), .B(n722), .Y(PRODUCT[24]) );
  OAI22XL U1120 ( .A0(n729), .A1(n754), .B0(n1078), .B1(n728), .Y(n741) );
  ADDHXL U1121 ( .A(n731), .B(n730), .CO(n702), .S(n740) );
  XNOR2X1 U1122 ( .A(B[1]), .B(n1199), .Y(n757) );
  OAI22X1 U1123 ( .A0(n988), .A1(n757), .B0(n732), .B1(n1175), .Y(n756) );
  CMPR32X1 U1124 ( .A(n741), .B(n739), .C(n740), .CO(n742), .S(n769) );
  CMPR32X1 U1125 ( .A(n744), .B(n743), .C(n742), .CO(n1168), .S(n773) );
  XNOR2X1 U1126 ( .A(n1205), .B(n1017), .Y(n785) );
  OAI22XL U1127 ( .A0(n11), .A1(n785), .B0(n1243), .B1(n751), .Y(n786) );
  XNOR2X1 U1128 ( .A(n1013), .B(n986), .Y(n789) );
  OAI22X1 U1129 ( .A0(n988), .A1(n792), .B0(n757), .B1(n968), .Y(n791) );
  XNOR2XL U1130 ( .A(n884), .B(A[4]), .Y(n758) );
  OAI22X2 U1131 ( .A0(n175), .A1(n795), .B0(n1058), .B1(n759), .Y(n798) );
  CMPR32X1 U1132 ( .A(n768), .B(n767), .C(n766), .CO(n1171), .S(n810) );
  ADDFHX1 U1133 ( .A(n771), .B(n770), .CI(n769), .CO(n774), .S(n809) );
  NAND2XL U1134 ( .A(n776), .B(n775), .Y(mult_x_1_n245) );
  INVXL U1135 ( .A(n777), .Y(n779) );
  INVXL U1136 ( .A(n717), .Y(n778) );
  XNOR2X1 U1137 ( .A(n1205), .B(n984), .Y(n814) );
  XNOR2X1 U1138 ( .A(n1013), .B(A[11]), .Y(n818) );
  OAI22XL U1139 ( .A0(n1080), .A1(n818), .B0(n1078), .B1(n789), .Y(n802) );
  XNOR2X1 U1140 ( .A(B[1]), .B(A[18]), .Y(n821) );
  OAI22X1 U1141 ( .A0(n988), .A1(n821), .B0(n792), .B1(n1175), .Y(n820) );
  XNOR2XL U1142 ( .A(n884), .B(A[3]), .Y(n793) );
  OAI22X2 U1143 ( .A0(n173), .A1(n825), .B0(n1058), .B1(n795), .Y(n827) );
  ADDFHX4 U1144 ( .A(n799), .B(n798), .CI(n797), .CO(n808), .S(n836) );
  CMPR32X1 U1145 ( .A(n802), .B(n801), .C(n800), .CO(n803), .S(n835) );
  XNOR2X1 U1146 ( .A(n1037), .B(n986), .Y(n852) );
  OAI22X1 U1147 ( .A0(n1262), .A1(n824), .B0(n1263), .B1(n813), .Y(n850) );
  OAI22XL U1148 ( .A0(n1080), .A1(n847), .B0(n1078), .B1(n818), .Y(n831) );
  XNOR2X1 U1149 ( .A(B[1]), .B(A[17]), .Y(n855) );
  OAI22X1 U1150 ( .A0(n988), .A1(n855), .B0(n821), .B1(n1175), .Y(n854) );
  XNOR2XL U1151 ( .A(n884), .B(A[2]), .Y(n822) );
  XNOR2X1 U1152 ( .A(n1041), .B(n984), .Y(n857) );
  OAI22X2 U1153 ( .A0(n1262), .A1(n883), .B0(n1263), .B1(n824), .Y(n892) );
  CMPR32X1 U1154 ( .A(n831), .B(n830), .C(n829), .CO(n832), .S(n869) );
  ADDFX2 U1155 ( .A(n834), .B(n833), .CI(n832), .CO(n846), .S(n872) );
  NAND2XL U1156 ( .A(n842), .B(n841), .Y(mult_x_1_n263) );
  NAND2X1 U1157 ( .A(n219), .B(n1391), .Y(n843) );
  OAI22X1 U1158 ( .A0(n1080), .A1(n888), .B0(n1078), .B1(n847), .Y(n862) );
  XNOR2XL U1159 ( .A(n1205), .B(n975), .Y(n886) );
  OAI22XL U1160 ( .A0(n11), .A1(n886), .B0(n1243), .B1(n848), .Y(n860) );
  XNOR2X1 U1161 ( .A(B[1]), .B(A[16]), .Y(n895) );
  XNOR2X1 U1162 ( .A(n12), .B(n927), .Y(n897) );
  OAI22X2 U1163 ( .A0(n173), .A1(n897), .B0(n1058), .B1(n858), .Y(n900) );
  CMPR32X1 U1164 ( .A(n862), .B(n861), .C(n860), .CO(n868), .S(n912) );
  CMPR32X1 U1165 ( .A(n865), .B(n864), .C(n863), .CO(n866), .S(n911) );
  ADDFX2 U1166 ( .A(n868), .B(n867), .CI(n866), .CO(n882), .S(n915) );
  NAND2XL U1167 ( .A(n875), .B(n874), .Y(mult_x_1_n266) );
  INVXL U1168 ( .A(n1392), .Y(n879) );
  XNOR2X1 U1169 ( .A(n1250), .B(A[2]), .Y(n896) );
  XNOR2X1 U1170 ( .A(n884), .B(n970), .Y(n885) );
  OAI22XL U1171 ( .A0(n11), .A1(n898), .B0(n1243), .B1(n886), .Y(n905) );
  XNOR2X1 U1172 ( .A(n1037), .B(n1015), .Y(n904) );
  ADDHXL U1173 ( .A(n890), .B(n889), .CO(n863), .S(n908) );
  XNOR2X1 U1174 ( .A(B[1]), .B(n894), .Y(n928) );
  OAI22X2 U1175 ( .A0(n988), .A1(n928), .B0(n895), .B1(n1175), .Y(n933) );
  OAI22X1 U1176 ( .A0(n931), .A1(n936), .B0(n1263), .B1(n896), .Y(n932) );
  XNOR2X1 U1177 ( .A(n1013), .B(n984), .Y(n935) );
  XNOR2X1 U1178 ( .A(n12), .B(n967), .Y(n942) );
  OAI22XL U1179 ( .A0(n11), .A1(n938), .B0(n1243), .B1(n898), .Y(n945) );
  XNOR2X1 U1180 ( .A(n1041), .B(n975), .Y(n943) );
  XNOR2X1 U1181 ( .A(n1037), .B(n982), .Y(n944) );
  CMPR32X1 U1182 ( .A(n907), .B(n906), .C(n905), .CO(n926), .S(n962) );
  CMPR32X1 U1183 ( .A(n910), .B(n909), .C(n908), .CO(n925), .S(n961) );
  NOR2XL U1184 ( .A(n918), .B(n917), .Y(mult_x_1_n273) );
  INVXL U1185 ( .A(n1394), .Y(n919) );
  ADDFHX1 U1186 ( .A(n923), .B(n922), .CI(n921), .CO(n917), .S(n954) );
  CMPR32X1 U1187 ( .A(n926), .B(n925), .C(n924), .CO(n923), .S(n960) );
  OAI22X1 U1188 ( .A0(n988), .A1(n969), .B0(n928), .B1(n1175), .Y(n966) );
  OAI22XL U1189 ( .A0(n1080), .A1(n976), .B0(n1078), .B1(n935), .Y(n981) );
  XNOR2XL U1190 ( .A(n1250), .B(n1176), .Y(n937) );
  XNOR2X1 U1191 ( .A(n1205), .B(A[2]), .Y(n971) );
  OAI22XL U1192 ( .A0(n11), .A1(n971), .B0(n1243), .B1(n938), .Y(n979) );
  XNOR2X1 U1193 ( .A(n12), .B(n986), .Y(n978) );
  XNOR2X1 U1194 ( .A(n1041), .B(A[4]), .Y(n977) );
  XNOR2X1 U1195 ( .A(n1037), .B(n1017), .Y(n985) );
  NOR2XL U1196 ( .A(n954), .B(n953), .Y(mult_x_1_n276) );
  INVXL U1197 ( .A(n1396), .Y(n956) );
  CMPR32X1 U1198 ( .A(n974), .B(n973), .C(n972), .CO(n993), .S(n1023) );
  OAI22X1 U1199 ( .A0(n1080), .A1(n1014), .B0(n1078), .B1(n976), .Y(n1021) );
  XNOR2X1 U1200 ( .A(n1041), .B(A[3]), .Y(n1042) );
  XNOR2XL U1201 ( .A(n12), .B(A[11]), .Y(n1016) );
  CMPR32X1 U1202 ( .A(n981), .B(n980), .C(n979), .CO(n972), .S(n1034) );
  XNOR2X1 U1203 ( .A(n1037), .B(n984), .Y(n1038) );
  CMPR32X1 U1204 ( .A(n1000), .B(n999), .C(n998), .CO(n994), .S(n1026) );
  CMPR32X1 U1205 ( .A(n1003), .B(n1002), .C(n1001), .CO(n991), .S(n1032) );
  CMPR32X1 U1206 ( .A(n1006), .B(n1005), .C(n1004), .CO(n1003), .S(n1066) );
  CMPR32X1 U1207 ( .A(n1009), .B(n1008), .C(n1007), .CO(n1024), .S(n1065) );
  CMPR32X1 U1208 ( .A(n1012), .B(n1011), .C(n1010), .CO(n1007), .S(n1071) );
  XNOR2X1 U1209 ( .A(n12), .B(n1015), .Y(n1057) );
  NOR2XL U1210 ( .A(n1026), .B(n1025), .Y(mult_x_1_n286) );
  OAI21XL U1211 ( .A0(n216), .A1(n1402), .B0(n1407), .Y(n1029) );
  INVXL U1212 ( .A(n1400), .Y(n1027) );
  NAND2XL U1213 ( .A(n1027), .B(n1401), .Y(n1028) );
  XNOR2X1 U1214 ( .A(n1029), .B(n1028), .Y(PRODUCT[16]) );
  CMPR32X1 U1215 ( .A(n1032), .B(n1031), .C(n1030), .CO(n1025), .S(n1068) );
  XNOR2X1 U1216 ( .A(n1037), .B(n1036), .Y(n1054) );
  OAI22X1 U1217 ( .A0(n11), .A1(n1040), .B0(n1243), .B1(n1039), .Y(n1073) );
  CMPR32X1 U1218 ( .A(n1045), .B(n1044), .C(n1043), .CO(n1033), .S(n1086) );
  ADDHXL U1219 ( .A(n1047), .B(n1046), .CO(n1043), .S(n1090) );
  NOR2XL U1220 ( .A(n1068), .B(n1067), .Y(mult_x_1_n292) );
  NAND2XL U1221 ( .A(n1068), .B(n1067), .Y(mult_x_1_n293) );
  ADDHXL U1222 ( .A(n1082), .B(n1081), .CO(n1120), .S(n1094) );
  CMPR32X1 U1223 ( .A(n1096), .B(n1095), .C(n1094), .CO(n1126), .S(n1140) );
  CMPR32X1 U1224 ( .A(n1099), .B(n1098), .C(n1097), .CO(n1088), .S(n1125) );
  CMPR32X1 U1225 ( .A(n1102), .B(n1101), .C(n1100), .CO(n1107), .S(n1116) );
  NOR2XL U1226 ( .A(n1110), .B(n1109), .Y(mult_x_1_n306) );
  CMPR32X1 U1227 ( .A(n1105), .B(n1104), .C(n1103), .CO(n1067), .S(n1112) );
  OR2X2 U1228 ( .A(n1112), .B(n1111), .Y(n1194) );
  NAND2XL U1229 ( .A(n1194), .B(n1115), .Y(mult_x_1_n295) );
  INVXL U1230 ( .A(mult_x_1_n307), .Y(n1114) );
  NAND2XL U1231 ( .A(n1112), .B(n1111), .Y(n1193) );
  INVXL U1232 ( .A(n1193), .Y(n1113) );
  NAND2XL U1233 ( .A(n1115), .B(mult_x_1_n307), .Y(mult_x_1_n84) );
  ADDFHX1 U1234 ( .A(n1118), .B(n1117), .CI(n1116), .CO(n1109), .S(n1129) );
  NAND2XL U1235 ( .A(n1189), .B(n1187), .Y(mult_x_1_n85) );
  XNOR2X1 U1236 ( .A(n1358), .B(n1406), .Y(PRODUCT[12]) );
  OAI21XL U1237 ( .A0(n1131), .A1(n1145), .B0(n1130), .Y(n1132) );
  INVXL U1238 ( .A(n1192), .Y(mult_x_1_n321) );
  CMPR32X1 U1239 ( .A(n1140), .B(n1139), .C(n1138), .CO(n1142), .S(n351) );
  NOR2XL U1240 ( .A(n1143), .B(n1142), .Y(n1141) );
  INVXL U1241 ( .A(n1141), .Y(n1195) );
  AOI21XL U1242 ( .A0(mult_x_1_n321), .A1(n1195), .B0(n1188), .Y(mult_x_1_n316) );
  NAND2XL U1243 ( .A(n15), .B(n1145), .Y(n1146) );
  AOI21XL U1244 ( .A0(n1156), .A1(n1154), .B0(n1148), .Y(n1152) );
  XOR2X1 U1245 ( .A(n1152), .B(n1151), .Y(n1430) );
  NAND2XL U1246 ( .A(n1154), .B(n1153), .Y(n1155) );
  XNOR2X1 U1247 ( .A(n1156), .B(n1155), .Y(n1431) );
  ADDFHX1 U1248 ( .A(n1165), .B(n1164), .CI(n1163), .CO(n714), .S(
        mult_x_1_n554) );
  ADDFHX1 U1249 ( .A(n1171), .B(n1170), .CI(n1169), .CO(n775), .S(
        mult_x_1_n586) );
  INVXL U1250 ( .A(n1388), .Y(n1177) );
  INVXL U1251 ( .A(n1179), .Y(n1180) );
  NAND2XL U1252 ( .A(n1184), .B(n1183), .Y(n1185) );
  XNOR2X1 U1253 ( .A(n1186), .B(n1185), .Y(PRODUCT[25]) );
  NAND2XL U1254 ( .A(n1194), .B(n1193), .Y(mult_x_1_n83) );
  NAND2XL U1255 ( .A(n1195), .B(n14), .Y(mult_x_1_n86) );
  XNOR2XL U1256 ( .A(n1205), .B(A[24]), .Y(n1223) );
  CMPR32X1 U1257 ( .A(n1210), .B(n1209), .C(n1208), .CO(n1224), .S(n1198) );
  CMPR32X1 U1258 ( .A(n1213), .B(n1212), .C(n1211), .CO(n1214), .S(n1197) );
  CMPR32X1 U1259 ( .A(n1219), .B(n1218), .C(n1217), .CO(n1233), .S(n1216) );
  XNOR2XL U1260 ( .A(n1205), .B(A[25]), .Y(n1241) );
  OAI22X1 U1261 ( .A0(n11), .A1(n1223), .B0(n1243), .B1(n1241), .Y(n1254) );
  CMPR32X1 U1262 ( .A(n1226), .B(n1225), .C(n1224), .CO(n1231), .S(n1215) );
  CMPR32X1 U1263 ( .A(n1233), .B(n1232), .C(n1231), .CO(n1245), .S(n1227) );
  XNOR2XL U1264 ( .A(n1234), .B(A[24]), .Y(n1251) );
  CMPR32X1 U1265 ( .A(n1238), .B(n1237), .C(n1236), .CO(n1247), .S(n1232) );
  CMPR32X1 U1266 ( .A(n1248), .B(n1247), .C(n1246), .CO(n1272), .S(n1244) );
  XNOR2XL U1267 ( .A(n1250), .B(A[25]), .Y(n1260) );
  CMPR32X1 U1268 ( .A(n1254), .B(n1253), .C(n1252), .CO(n1255), .S(n1246) );
  CMPR32X1 U1269 ( .A(n1257), .B(n1256), .C(n1255), .CO(n1268), .S(n1271) );
  XNOR2XL U1270 ( .A(n884), .B(A[24]), .Y(n1258) );
  XOR3X2 U1271 ( .A(n1266), .B(n1265), .C(n1264), .Y(n1267) );
  OAI21XL U1272 ( .A0(n1278), .A1(n1373), .B0(n1277), .Y(n1344) );
  OAI21XL U1273 ( .A0(n1347), .A1(n1280), .B0(n1279), .Y(n1314) );
  OAI21XL U1274 ( .A0(n1350), .A1(n1283), .B0(n1282), .Y(n1286) );
  OAI21XL U1275 ( .A0(n1350), .A1(n1288), .B0(n1287), .Y(n1291) );
  OAI21XL U1276 ( .A0(n1364), .A1(n1367), .B0(n1365), .Y(n1311) );
  AOI21XL U1277 ( .A0(n180), .A1(n1307), .B0(n1311), .Y(n1292) );
  OAI21XL U1278 ( .A0(n1350), .A1(n1293), .B0(n1292), .Y(n1295) );
  OAI21XL U1279 ( .A0(n1305), .A1(n1302), .B0(n1303), .Y(n1301) );
  INVXL U1280 ( .A(n1297), .Y(n1299) );
  AOI21XL U1281 ( .A0(n180), .A1(n1313), .B0(n1312), .Y(n1315) );
  OAI21XL U1282 ( .A0(n1350), .A1(n1316), .B0(n1315), .Y(n1319) );
  XOR2XL U1283 ( .A(n1328), .B(n1327), .Y(n1436) );
  XNOR2XL U1284 ( .A(n1332), .B(n1331), .Y(n1435) );
  XOR2XL U1285 ( .A(n1337), .B(n1336), .Y(n1434) );
  OAI21XL U1286 ( .A0(n1341), .A1(n1360), .B0(n1361), .Y(n1342) );
  OAI21XL U1287 ( .A0(n1347), .A1(n1346), .B0(n1345), .Y(n1348) );
  OAI21XL U1288 ( .A0(n1350), .A1(n225), .B0(n1349), .Y(n1351) );
  XNOR2XL U1289 ( .A(n1351), .B(n1359), .Y(PRODUCT[40]) );
endmodule


module FFT2048_DW02_mult_2_stage_J1_6 ( A, B, TC, CLK, PRODUCT );
  input [25:0] A;
  input [16:0] B;
  output [42:0] PRODUCT;
  input TC, CLK;
  wire   n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, mult_x_1_n569, mult_x_1_n554, mult_x_1_n537,
         mult_x_1_n522, mult_x_1_n316, mult_x_1_n309, mult_x_1_n308,
         mult_x_1_n301, mult_x_1_n294, mult_x_1_n291, mult_x_1_n290,
         mult_x_1_n287, mult_x_1_n286, mult_x_1_n282, mult_x_1_n281,
         mult_x_1_n277, mult_x_1_n276, mult_x_1_n274, mult_x_1_n273,
         mult_x_1_n266, mult_x_1_n265, mult_x_1_n263, mult_x_1_n262,
         mult_x_1_n252, mult_x_1_n251, mult_x_1_n245, mult_x_1_n244,
         mult_x_1_n227, mult_x_1_n226, mult_x_1_n207, mult_x_1_n206,
         mult_x_1_n198, mult_x_1_n197, mult_x_1_n195, mult_x_1_n194,
         mult_x_1_n184, mult_x_1_n183, mult_x_1_n177, mult_x_1_n176,
         mult_x_1_n170, mult_x_1_n169, mult_x_1_n161, mult_x_1_n160,
         mult_x_1_n152, mult_x_1_n151, mult_x_1_n137, mult_x_1_n136,
         mult_x_1_n130, mult_x_1_n129, mult_x_1_n121, mult_x_1_n120,
         mult_x_1_n110, mult_x_1_n109, mult_x_1_n85, mult_x_1_n84,
         mult_x_1_n83, mult_x_1_n82, mult_x_1_n58, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295;

  DFFHQXL mult_x_1_clk_r_REG18_S1 ( .D(mult_x_1_n160), .CK(CLK), .Q(n1250) );
  DFFHQXL mult_x_1_clk_r_REG16_S1 ( .D(mult_x_1_n169), .CK(CLK), .Q(n1252) );
  DFFHQX4 mult_x_1_clk_r_REG30_S1 ( .D(mult_x_1_n569), .CK(CLK), .Q(n1295) );
  DFFHQX4 mult_x_1_clk_r_REG0_S1 ( .D(mult_x_1_n554), .CK(CLK), .Q(n1294) );
  DFFHQX4 mult_x_1_clk_r_REG3_S1 ( .D(mult_x_1_n537), .CK(CLK), .Q(n1293) );
  DFFHQX4 mult_x_1_clk_r_REG55_S1 ( .D(mult_x_1_n309), .CK(CLK), .Q(n1290) );
  DFFHQX4 mult_x_1_clk_r_REG48_S1 ( .D(mult_x_1_n291), .CK(CLK), .Q(n1287) );
  DFFHQX4 mult_x_1_clk_r_REG49_S1 ( .D(mult_x_1_n290), .CK(CLK), .Q(n1281) );
  DFFHQX4 mult_x_1_clk_r_REG45_S1 ( .D(mult_x_1_n287), .CK(CLK), .Q(n1280) );
  DFFHQX4 mult_x_1_clk_r_REG44_S1 ( .D(mult_x_1_n281), .CK(CLK), .Q(n1277) );
  DFFHQX4 mult_x_1_clk_r_REG40_S1 ( .D(mult_x_1_n273), .CK(CLK), .Q(n1273) );
  DFFHQX4 mult_x_1_clk_r_REG37_S1 ( .D(mult_x_1_n266), .CK(CLK), .Q(n1272) );
  DFFHQX4 mult_x_1_clk_r_REG36_S1 ( .D(mult_x_1_n262), .CK(CLK), .Q(n1269) );
  DFFHQXL mult_x_1_clk_r_REG5_S1 ( .D(mult_x_1_n207), .CK(CLK), .Q(n1263) );
  DFFHQXL clk_r_REG57_S1 ( .D(n1309), .CK(CLK), .Q(PRODUCT[12]) );
  DFFHQX4 mult_x_1_clk_r_REG43_S1 ( .D(mult_x_1_n282), .CK(CLK), .Q(n1278) );
  DFFHQXL mult_x_1_clk_r_REG51_S1 ( .D(mult_x_1_n294), .CK(CLK), .Q(n1288) );
  DFFHQXL mult_x_1_clk_r_REG13_S1 ( .D(mult_x_1_n177), .CK(CLK), .Q(n1255) );
  DFFHQXL clk_r_REG59_S1 ( .D(n1310), .CK(CLK), .Q(PRODUCT[11]) );
  DFFHQXL mult_x_1_clk_r_REG53_S1 ( .D(mult_x_1_n301), .CK(CLK), .Q(n1289) );
  DFFHQX4 mult_x_1_clk_r_REG39_S1 ( .D(mult_x_1_n274), .CK(CLK), .Q(n1274) );
  DFFHQXL clk_r_REG61_S1 ( .D(n1312), .CK(CLK), .Q(PRODUCT[9]) );
  DFFHQXL mult_x_1_clk_r_REG50_S1 ( .D(mult_x_1_n83), .CK(CLK), .Q(n1283) );
  DFFHQXL clk_r_REG60_S1 ( .D(n1311), .CK(CLK), .Q(PRODUCT[10]) );
  DFFHQXL mult_x_1_clk_r_REG8_S1 ( .D(mult_x_1_n197), .CK(CLK), .Q(n1260) );
  DFFHQXL mult_x_1_clk_r_REG17_S1 ( .D(mult_x_1_n161), .CK(CLK), .Q(n1251) );
  DFFHQXL mult_x_1_clk_r_REG47_S1 ( .D(mult_x_1_n82), .CK(CLK), .Q(n1282) );
  DFFHQXL mult_x_1_clk_r_REG21_S1 ( .D(mult_x_1_n137), .CK(CLK), .Q(n1247) );
  DFFHQX4 mult_x_1_clk_r_REG2_S1 ( .D(mult_x_1_n226), .CK(CLK), .Q(n1264) );
  DFFHQX4 mult_x_1_clk_r_REG35_S1 ( .D(mult_x_1_n263), .CK(CLK), .Q(n1270) );
  DFFHQXL mult_x_1_clk_r_REG31_S1 ( .D(mult_x_1_n245), .CK(CLK), .Q(n1267) );
  DFFHQXL mult_x_1_clk_r_REG1_S1 ( .D(mult_x_1_n227), .CK(CLK), .Q(n1265) );
  DFFHQXL clk_r_REG62_S1 ( .D(n1313), .CK(CLK), .Q(PRODUCT[8]) );
  DFFHQXL clk_r_REG63_S1 ( .D(n1314), .CK(CLK), .Q(PRODUCT[7]) );
  DFFHQXL clk_r_REG64_S1 ( .D(n1315), .CK(CLK), .Q(PRODUCT[6]) );
  DFFHQXL clk_r_REG65_S1 ( .D(n1316), .CK(CLK), .Q(PRODUCT[5]) );
  DFFHQXL clk_r_REG66_S1 ( .D(n1317), .CK(CLK), .Q(PRODUCT[4]) );
  DFFHQXL clk_r_REG67_S1 ( .D(n1318), .CK(CLK), .Q(PRODUCT[3]) );
  DFFHQXL clk_r_REG68_S1 ( .D(n1319), .CK(CLK), .Q(PRODUCT[2]) );
  DFFHQXL clk_r_REG69_S1 ( .D(n1320), .CK(CLK), .Q(PRODUCT[1]) );
  DFFHQXL clk_r_REG70_S1 ( .D(n1321), .CK(CLK), .Q(PRODUCT[0]) );
  DFFHQXL mult_x_1_clk_r_REG11_S1 ( .D(mult_x_1_n184), .CK(CLK), .Q(n1257) );
  DFFHQXL mult_x_1_clk_r_REG9_S1 ( .D(mult_x_1_n195), .CK(CLK), .Q(n1259) );
  DFFHQX1 mult_x_1_clk_r_REG54_S1 ( .D(mult_x_1_n85), .CK(CLK), .Q(n1285) );
  DFFHQXL mult_x_1_clk_r_REG12_S1 ( .D(mult_x_1_n183), .CK(CLK), .Q(n1256) );
  DFFHQXL mult_x_1_clk_r_REG15_S1 ( .D(mult_x_1_n170), .CK(CLK), .Q(n1253) );
  DFFHQXL mult_x_1_clk_r_REG19_S1 ( .D(mult_x_1_n152), .CK(CLK), .Q(n1249) );
  DFFHQXL mult_x_1_clk_r_REG23_S1 ( .D(mult_x_1_n130), .CK(CLK), .Q(n1245) );
  DFFHQXL mult_x_1_clk_r_REG24_S1 ( .D(mult_x_1_n129), .CK(CLK), .Q(n1244) );
  DFFHQXL mult_x_1_clk_r_REG25_S1 ( .D(mult_x_1_n121), .CK(CLK), .Q(n1243) );
  DFFHQXL mult_x_1_clk_r_REG26_S1 ( .D(mult_x_1_n120), .CK(CLK), .Q(n1242) );
  DFFHQXL mult_x_1_clk_r_REG27_S1 ( .D(mult_x_1_n110), .CK(CLK), .Q(n1241) );
  DFFHQXL mult_x_1_clk_r_REG28_S1 ( .D(mult_x_1_n109), .CK(CLK), .Q(n1240) );
  DFFHQXL mult_x_1_clk_r_REG29_S1 ( .D(mult_x_1_n58), .CK(CLK), .Q(n1239) );
  DFFHQX1 mult_x_1_clk_r_REG58_S1 ( .D(mult_x_1_n316), .CK(CLK), .Q(n1291) );
  DFFHQXL mult_x_1_clk_r_REG20_S1 ( .D(mult_x_1_n151), .CK(CLK), .Q(n1248) );
  DFFHQXL mult_x_1_clk_r_REG22_S1 ( .D(mult_x_1_n136), .CK(CLK), .Q(n1246) );
  DFFHQX1 mult_x_1_clk_r_REG52_S1 ( .D(mult_x_1_n84), .CK(CLK), .Q(n1284) );
  DFFHQXL mult_x_1_clk_r_REG56_S1 ( .D(mult_x_1_n308), .CK(CLK), .Q(n1238) );
  DFFHQXL mult_x_1_clk_r_REG7_S1 ( .D(mult_x_1_n198), .CK(CLK), .Q(n1261) );
  DFFHQX2 mult_x_1_clk_r_REG33_S1 ( .D(mult_x_1_n252), .CK(CLK), .Q(n1268) );
  DFFHQX2 mult_x_1_clk_r_REG46_S1 ( .D(mult_x_1_n286), .CK(CLK), .Q(n1279) );
  DFFHQX2 mult_x_1_clk_r_REG32_S1 ( .D(mult_x_1_n244), .CK(CLK), .Q(n1266) );
  DFFHQXL mult_x_1_clk_r_REG14_S1 ( .D(mult_x_1_n176), .CK(CLK), .Q(n1254) );
  DFFHQX1 mult_x_1_clk_r_REG6_S1 ( .D(mult_x_1_n206), .CK(CLK), .Q(n1262) );
  DFFHQX2 mult_x_1_clk_r_REG34_S1 ( .D(mult_x_1_n251), .CK(CLK), .Q(n1286) );
  DFFHQX2 mult_x_1_clk_r_REG42_S1 ( .D(mult_x_1_n276), .CK(CLK), .Q(n1275) );
  DFFHQX2 mult_x_1_clk_r_REG4_S1 ( .D(mult_x_1_n522), .CK(CLK), .Q(n1292) );
  DFFHQX1 mult_x_1_clk_r_REG38_S1 ( .D(mult_x_1_n265), .CK(CLK), .Q(n1271) );
  DFFHQX1 mult_x_1_clk_r_REG41_S1 ( .D(mult_x_1_n277), .CK(CLK), .Q(n1276) );
  DFFHQX1 mult_x_1_clk_r_REG10_S1 ( .D(mult_x_1_n194), .CK(CLK), .Q(n1258) );
  CMPR32X1 U1 ( .A(n932), .B(n931), .C(n930), .CO(n923), .S(n972) );
  ADDFHX1 U2 ( .A(n704), .B(n703), .CI(n702), .CO(n1069), .S(n729) );
  ADDFHX1 U3 ( .A(n690), .B(n689), .CI(n688), .CO(n1066), .S(n1068) );
  ADDFHX1 U4 ( .A(n798), .B(n797), .CI(n796), .CO(n765), .S(n803) );
  ADDFHX1 U5 ( .A(n820), .B(n819), .CI(n818), .CO(n804), .S(n844) );
  XNOR2X2 U6 ( .A(n550), .B(n551), .Y(n28) );
  ADDFHX2 U7 ( .A(n572), .B(n571), .CI(n570), .CO(n550), .S(n1059) );
  CMPR32X1 U8 ( .A(n621), .B(n620), .C(n619), .CO(n624), .S(n651) );
  CMPR32X1 U9 ( .A(n356), .B(n355), .C(n354), .CO(n398), .S(n393) );
  ADDFHX1 U10 ( .A(n720), .B(n719), .CI(n718), .CO(n704), .S(n758) );
  ADDFHX1 U11 ( .A(n1003), .B(n1002), .CI(n1001), .CO(n999), .S(n1020) );
  ADDFHX2 U12 ( .A(n531), .B(n530), .CI(n529), .CO(n551), .S(n571) );
  ADDFX2 U13 ( .A(n554), .B(n553), .CI(n552), .CO(n543), .S(n1061) );
  CMPR32X1 U14 ( .A(n678), .B(n677), .C(n676), .CO(n687), .S(n719) );
  CMPR32X1 U15 ( .A(n667), .B(n666), .C(n665), .CO(n647), .S(n683) );
  ADDFX2 U16 ( .A(n812), .B(n811), .CI(n810), .CO(n792), .S(n831) );
  ADDFHX1 U17 ( .A(n998), .B(n997), .CI(n996), .CO(n976), .S(n1001) );
  ADDFHX1 U18 ( .A(n1079), .B(n1078), .CI(n1077), .CO(n1080), .S(n1036) );
  ADDFHX1 U19 ( .A(n907), .B(n906), .CI(n905), .CO(n922), .S(n969) );
  ADDFHX2 U20 ( .A(n1027), .B(n1026), .CI(n1025), .CO(n1075), .S(n1078) );
  CMPR32X1 U21 ( .A(n467), .B(n466), .C(n465), .CO(n449), .S(n480) );
  ADDFX2 U22 ( .A(n600), .B(n599), .CI(n598), .CO(n569), .S(n617) );
  ADDFHX1 U23 ( .A(n947), .B(n946), .CI(n945), .CO(n970), .S(n997) );
  ADDFX2 U24 ( .A(n511), .B(n510), .CI(n509), .CO(n495), .S(n530) );
  CMPR32X1 U25 ( .A(n430), .B(n429), .C(n428), .CO(n448), .S(n465) );
  CMPR32X1 U26 ( .A(n427), .B(n426), .C(n425), .CO(n411), .S(n466) );
  ADDFHX1 U27 ( .A(n267), .B(n266), .CI(n265), .CO(n274), .S(n273) );
  CMPR32X1 U28 ( .A(n899), .B(n898), .C(n897), .CO(n907), .S(n946) );
  ADDFHX1 U29 ( .A(n461), .B(n460), .CI(n459), .CO(n452), .S(n494) );
  ADDFHX2 U30 ( .A(n264), .B(n263), .CI(n262), .CO(n1032), .S(n265) );
  ADDFHX1 U31 ( .A(n261), .B(n260), .CI(n259), .CO(n266), .S(n268) );
  ADDFHX2 U32 ( .A(n205), .B(n204), .CI(n203), .CO(n260), .S(n214) );
  BUFX8 U33 ( .A(n457), .Y(n11) );
  BUFX8 U34 ( .A(n859), .Y(n1143) );
  BUFX4 U35 ( .A(n244), .Y(n7) );
  ADDFX2 U36 ( .A(n255), .B(n254), .CI(n253), .CO(n1014), .S(n256) );
  BUFX8 U37 ( .A(B[13]), .Y(n225) );
  BUFX3 U38 ( .A(n35), .Y(n964) );
  CLKBUFX3 U39 ( .A(n118), .Y(n9) );
  BUFX4 U40 ( .A(n155), .Y(n949) );
  CLKINVX3 U41 ( .A(n156), .Y(n900) );
  BUFX3 U42 ( .A(n96), .Y(n12) );
  BUFX3 U43 ( .A(n484), .Y(n953) );
  NAND2X1 U44 ( .A(n146), .B(n155), .Y(n807) );
  INVX1 U45 ( .A(B[5]), .Y(n98) );
  INVX1 U46 ( .A(B[9]), .Y(n156) );
  XNOR2X2 U47 ( .A(B[10]), .B(B[9]), .Y(n484) );
  XOR2X1 U48 ( .A(n39), .B(n32), .Y(PRODUCT[31]) );
  XNOR2X1 U49 ( .A(n365), .B(n364), .Y(PRODUCT[33]) );
  OAI21XL U50 ( .A0(n1236), .A1(n441), .B0(n440), .Y(n39) );
  XOR2X1 U51 ( .A(n505), .B(n1236), .Y(PRODUCT[29]) );
  XNOR2X1 U52 ( .A(n727), .B(n726), .Y(PRODUCT[23]) );
  XNOR2X1 U53 ( .A(n594), .B(n593), .Y(PRODUCT[26]) );
  XNOR2X1 U54 ( .A(n763), .B(n762), .Y(PRODUCT[22]) );
  OAI21XL U55 ( .A0(n1264), .A1(n586), .B0(n1265), .Y(n83) );
  OAI21X1 U56 ( .A0(n1269), .A1(n1272), .B0(n1270), .Y(n657) );
  NOR2X1 U57 ( .A(n1295), .B(n1294), .Y(n584) );
  OAI22X1 U58 ( .A0(n951), .A1(n524), .B0(n949), .B1(n512), .Y(n540) );
  OAI21XL U59 ( .A0(n1232), .A1(n1158), .B0(n1157), .Y(n1196) );
  AND2X1 U60 ( .A(n470), .B(n1259), .Y(n33) );
  XNOR2XL U61 ( .A(n842), .B(n841), .Y(PRODUCT[20]) );
  XNOR2XL U62 ( .A(n936), .B(A[2]), .Y(n92) );
  XNOR2XL U63 ( .A(n910), .B(A[2]), .Y(n246) );
  XNOR2XL U64 ( .A(n707), .B(A[15]), .Y(n745) );
  XNOR2XL U65 ( .A(n908), .B(A[1]), .Y(n125) );
  XNOR2XL U66 ( .A(B[16]), .B(A[8]), .Y(n528) );
  XNOR2XL U67 ( .A(n781), .B(A[20]), .Y(n637) );
  XNOR2XL U68 ( .A(n912), .B(A[23]), .Y(n383) );
  XNOR2XL U69 ( .A(n601), .B(A[23]), .Y(n344) );
  BUFX1 U70 ( .A(B[16]), .Y(n1138) );
  XNOR2XL U71 ( .A(n910), .B(A[24]), .Y(n293) );
  XNOR2XL U72 ( .A(n225), .B(A[14]), .Y(n508) );
  XNOR2XL U73 ( .A(n225), .B(A[13]), .Y(n534) );
  XNOR2XL U74 ( .A(n910), .B(A[22]), .Y(n342) );
  BUFX4 U75 ( .A(n283), .Y(n1140) );
  ADDFX2 U76 ( .A(n919), .B(n918), .CI(n917), .CO(n935), .S(n978) );
  ADDFX2 U77 ( .A(n772), .B(n771), .CI(n770), .CO(n754), .S(n791) );
  OAI21XL U78 ( .A0(n1053), .A1(n181), .B0(n180), .Y(n1042) );
  XOR2XL U79 ( .A(n1188), .B(n1187), .Y(n1315) );
  XOR2XL U80 ( .A(n1058), .B(n1057), .Y(n1312) );
  OR2X2 U81 ( .A(n275), .B(n274), .Y(n5) );
  OR2X2 U82 ( .A(n1081), .B(n1080), .Y(n6) );
  NOR2XL U83 ( .A(n548), .B(n547), .Y(mult_x_1_n197) );
  NOR2X1 U84 ( .A(n924), .B(n923), .Y(mult_x_1_n276) );
  XNOR2X1 U85 ( .A(n1166), .B(n1165), .Y(n1313) );
  NAND2BXL U86 ( .AN(n969), .B(n15), .Y(n14) );
  NAND2X1 U87 ( .A(n969), .B(n970), .Y(n13) );
  INVX1 U88 ( .A(n970), .Y(n15) );
  XOR2X1 U89 ( .A(n969), .B(n970), .Y(n16) );
  NOR2X1 U90 ( .A(n1140), .B(n817), .Y(n851) );
  NOR2X1 U91 ( .A(n1140), .B(n635), .Y(n669) );
  OAI22XL U92 ( .A0(n8), .A1(n675), .B0(n12), .B1(n638), .Y(n676) );
  OAI22XL U93 ( .A0(n8), .A1(n808), .B0(n12), .B1(n745), .Y(n784) );
  NOR2BX1 U94 ( .AN(A[0]), .B(n953), .Y(n194) );
  OAI22XL U95 ( .A0(n8), .A1(n609), .B0(n12), .B1(n557), .Y(n610) );
  NAND2X1 U96 ( .A(n224), .B(n227), .Y(n244) );
  OR2XL U97 ( .A(n114), .B(n113), .Y(n1203) );
  NAND2BXL U98 ( .AN(n84), .B(n63), .Y(n62) );
  NAND2X1 U99 ( .A(n89), .B(n783), .Y(n118) );
  NAND2XL U100 ( .A(n58), .B(n1272), .Y(n763) );
  NAND2XL U101 ( .A(n82), .B(n59), .Y(n58) );
  INVXL U102 ( .A(n280), .Y(n585) );
  NAND2X1 U103 ( .A(n363), .B(n1253), .Y(n364) );
  AND2X2 U104 ( .A(n442), .B(n1257), .Y(n32) );
  AND2X2 U105 ( .A(n85), .B(n1263), .Y(n34) );
  INVX1 U106 ( .A(n401), .Y(n440) );
  INVX1 U107 ( .A(n1279), .Y(n926) );
  INVX1 U108 ( .A(n1287), .Y(n37) );
  INVX1 U109 ( .A(n1242), .Y(n1192) );
  INVX1 U110 ( .A(n1248), .Y(n1153) );
  XOR2X1 U111 ( .A(n1052), .B(n1051), .Y(n1311) );
  XNOR2X1 U112 ( .A(n1179), .B(n1178), .Y(n1314) );
  INVX1 U113 ( .A(n271), .Y(n1040) );
  INVX1 U114 ( .A(n1038), .Y(n1039) );
  NAND2X1 U115 ( .A(n1020), .B(n1019), .Y(n1086) );
  OAI2BB1X1 U116 ( .A0N(n14), .A1N(n968), .B0(n13), .Y(n931) );
  NAND2X1 U117 ( .A(n273), .B(n272), .Y(n1038) );
  NAND2X1 U118 ( .A(n221), .B(n220), .Y(n1044) );
  XOR2X1 U119 ( .A(n968), .B(n16), .Y(n975) );
  INVXL U120 ( .A(n922), .Y(n24) );
  NOR2X1 U121 ( .A(n141), .B(n140), .Y(n1184) );
  NAND2X1 U122 ( .A(n141), .B(n140), .Y(n1185) );
  ADDFHX1 U123 ( .A(n1024), .B(n1023), .CI(n1022), .CO(n1016), .S(n1079) );
  OAI2BB1XL U124 ( .A0N(n11), .A1N(n1143), .B0(n1142), .Y(n1144) );
  NOR2X1 U125 ( .A(n1140), .B(n1103), .Y(n1116) );
  NOR2X1 U126 ( .A(n1140), .B(n302), .Y(n1101) );
  NOR2X1 U127 ( .A(n1140), .B(n1127), .Y(n1137) );
  NOR2X1 U128 ( .A(n1140), .B(n284), .Y(n308) );
  NOR2X1 U129 ( .A(n1140), .B(n1118), .Y(n1131) );
  NOR2X1 U130 ( .A(n1140), .B(n847), .Y(n871) );
  NOR2X1 U131 ( .A(n1140), .B(n316), .Y(n331) );
  NOR2X1 U132 ( .A(n1140), .B(n317), .Y(n353) );
  NOR2X1 U133 ( .A(n1140), .B(n345), .Y(n372) );
  NOR2X1 U134 ( .A(n1140), .B(n287), .Y(n298) );
  NOR2X1 U135 ( .A(n1140), .B(n382), .Y(n426) );
  NOR2X1 U136 ( .A(n1140), .B(n366), .Y(n389) );
  NOR2X1 U137 ( .A(n1140), .B(n515), .Y(n525) );
  NOR2XL U138 ( .A(n149), .B(n12), .Y(n45) );
  NAND2X1 U139 ( .A(n484), .B(n53), .Y(n200) );
  BUFX8 U140 ( .A(n95), .Y(n8) );
  XNOR2X1 U141 ( .A(n80), .B(n79), .Y(PRODUCT[35]) );
  XNOR2X1 U142 ( .A(n1201), .B(n1200), .Y(PRODUCT[39]) );
  CLKINVX3 U143 ( .A(n82), .Y(n802) );
  NOR2X1 U144 ( .A(n1225), .B(n1158), .Y(n1190) );
  NAND2BXL U145 ( .AN(n1266), .B(n22), .Y(n21) );
  NAND2X1 U146 ( .A(n405), .B(n1255), .Y(n406) );
  XNOR2X1 U147 ( .A(n1288), .B(n1282), .Y(PRODUCT[16]) );
  INVX1 U148 ( .A(n1250), .Y(n1151) );
  INVX1 U149 ( .A(n1271), .Y(n59) );
  NAND2XL U150 ( .A(n548), .B(n547), .Y(mult_x_1_n198) );
  NAND2XL U151 ( .A(n924), .B(n923), .Y(mult_x_1_n277) );
  NOR2X1 U152 ( .A(n1036), .B(n1035), .Y(n1034) );
  NAND2XL U153 ( .A(n972), .B(n971), .Y(mult_x_1_n282) );
  NAND2X1 U154 ( .A(n275), .B(n274), .Y(n1082) );
  ADDFHX2 U155 ( .A(n1033), .B(n1032), .CI(n1031), .CO(n1035), .S(n275) );
  ADDFHX2 U156 ( .A(n889), .B(n888), .CI(n887), .CO(n882), .S(n924) );
  ADDFHX1 U157 ( .A(n546), .B(n545), .CI(n544), .CO(n503), .S(n547) );
  NAND2XL U158 ( .A(n57), .B(n443), .Y(n56) );
  NAND2XL U159 ( .A(n444), .B(n445), .Y(n55) );
  ADDFHX2 U160 ( .A(n1076), .B(n1075), .CI(n1074), .CO(n1019), .S(n1081) );
  NOR2X1 U161 ( .A(n221), .B(n220), .Y(n1043) );
  NAND2XL U162 ( .A(n50), .B(n49), .Y(n1028) );
  ADDFHX2 U163 ( .A(n1018), .B(n1017), .CI(n1016), .CO(n1002), .S(n1074) );
  ADDFHX1 U164 ( .A(n270), .B(n269), .CI(n268), .CO(n272), .S(n221) );
  ADDFHX1 U165 ( .A(n881), .B(n880), .CI(n879), .CO(n843), .S(n887) );
  ADDFHX2 U166 ( .A(n433), .B(n432), .CI(n431), .CO(n435), .S(n443) );
  OR2XL U167 ( .A(n1148), .B(n1147), .Y(n1150) );
  ADDFHX2 U168 ( .A(n618), .B(n617), .CI(n616), .CO(n1064), .S(n652) );
  NAND2XL U169 ( .A(n538), .B(n31), .Y(n30) );
  ADDFHX2 U170 ( .A(n566), .B(n565), .CI(n564), .CO(n572), .S(n623) );
  ADDFHX1 U171 ( .A(n191), .B(n190), .CI(n189), .CO(n209), .S(n217) );
  ADDFHX1 U172 ( .A(n236), .B(n235), .CI(n234), .CO(n264), .S(n259) );
  ADDFHX1 U173 ( .A(n630), .B(n629), .CI(n628), .CO(n618), .S(n646) );
  OR2XL U174 ( .A(n539), .B(n540), .Y(n31) );
  NAND2XL U175 ( .A(n539), .B(n540), .Y(n29) );
  ADDFHX1 U176 ( .A(n960), .B(n959), .CI(n958), .CO(n945), .S(n1005) );
  ADDFHX1 U177 ( .A(n995), .B(n994), .CI(n993), .CO(n1006), .S(n1022) );
  ADDFHX1 U178 ( .A(n696), .B(n695), .CI(n694), .CO(n684), .S(n716) );
  ADDFHX1 U179 ( .A(n737), .B(n736), .CI(n735), .CO(n717), .S(n753) );
  OR2X2 U180 ( .A(n130), .B(n129), .Y(n128) );
  ADDFHX1 U181 ( .A(n166), .B(n165), .CI(n164), .CO(n170), .S(n172) );
  OAI2BB1XL U182 ( .A0N(n1121), .A1N(n7), .B0(n1120), .Y(n1130) );
  OAI2BB1XL U183 ( .A0N(n964), .A1N(n732), .B0(n320), .Y(n351) );
  AND2XL U184 ( .A(n1209), .B(n1208), .Y(n1320) );
  BUFX8 U185 ( .A(n200), .Y(n10) );
  XNOR2X1 U186 ( .A(n1162), .B(n1161), .Y(PRODUCT[36]) );
  OR2XL U187 ( .A(n1207), .B(n1206), .Y(n1209) );
  CLKINVX3 U188 ( .A(n896), .Y(n1113) );
  NAND2X1 U189 ( .A(n88), .B(n96), .Y(n95) );
  XNOR2X1 U190 ( .A(n1173), .B(n1172), .Y(PRODUCT[37]) );
  XNOR2X1 U191 ( .A(n1183), .B(n1182), .Y(PRODUCT[38]) );
  OR2XL U192 ( .A(n1225), .B(n1231), .Y(n1235) );
  NAND3BX2 U193 ( .AN(n71), .B(n61), .C(n60), .Y(n82) );
  INVXL U194 ( .A(n1268), .Y(n22) );
  XOR2X1 U195 ( .A(n1291), .B(n1285), .Y(PRODUCT[13]) );
  OAI22X1 U196 ( .A0(n8), .A1(n472), .B0(n12), .B1(n419), .Y(n461) );
  INVX1 U197 ( .A(B[5]), .Y(n367) );
  XNOR2X4 U198 ( .A(B[14]), .B(B[13]), .Y(n457) );
  AOI21X1 U199 ( .A0(n6), .A1(n1091), .B0(n1085), .Y(n1088) );
  OAI22X1 U200 ( .A0(n1143), .A1(n896), .B0(n11), .B1(n895), .Y(n938) );
  XNOR2X2 U201 ( .A(B[7]), .B(B[8]), .Y(n155) );
  NAND3X1 U202 ( .A(n1267), .B(n23), .C(n21), .Y(n589) );
  INVXL U203 ( .A(n589), .Y(n279) );
  XOR2X2 U204 ( .A(n17), .B(n33), .Y(PRODUCT[30]) );
  OAI21X1 U205 ( .A0(n1236), .A1(n1260), .B0(n1261), .Y(n17) );
  NOR2X4 U206 ( .A(n20), .B(n18), .Y(n1236) );
  NAND2X2 U207 ( .A(n48), .B(n19), .Y(n18) );
  NAND2BX1 U208 ( .AN(n68), .B(n589), .Y(n19) );
  AND2X2 U209 ( .A(n66), .B(n82), .Y(n20) );
  NAND2X1 U210 ( .A(n657), .B(n73), .Y(n23) );
  NOR2X1 U211 ( .A(n1266), .B(n1286), .Y(n73) );
  XNOR3X2 U212 ( .A(n24), .B(n921), .C(n920), .Y(n930) );
  NAND2X1 U213 ( .A(n26), .B(n25), .Y(n888) );
  NAND2X1 U214 ( .A(n921), .B(n922), .Y(n25) );
  OAI21XL U215 ( .A0(n921), .A1(n922), .B0(n920), .Y(n26) );
  OAI2BB1X1 U216 ( .A0N(n551), .A1N(n550), .B0(n27), .Y(n548) );
  OAI21XL U217 ( .A0(n550), .A1(n551), .B0(n549), .Y(n27) );
  XNOR2X1 U218 ( .A(n28), .B(n549), .Y(n574) );
  NAND2X1 U219 ( .A(n30), .B(n29), .Y(n529) );
  XOR3X2 U220 ( .A(n540), .B(n539), .C(n538), .Y(n567) );
  OAI22X1 U221 ( .A0(n951), .A1(n901), .B0(n949), .B1(n861), .Y(n916) );
  CLKINVX3 U222 ( .A(B[11]), .Y(n285) );
  XNOR2X1 U223 ( .A(n1128), .B(A[14]), .Y(n420) );
  XNOR2X1 U224 ( .A(n707), .B(A[24]), .Y(n419) );
  CLKINVX3 U225 ( .A(n367), .Y(n707) );
  CLKINVX3 U226 ( .A(B[7]), .Y(n318) );
  XNOR2X1 U227 ( .A(n910), .B(A[16]), .Y(n483) );
  OAI22X1 U228 ( .A0(n10), .A1(n607), .B0(n953), .B1(n555), .Y(n612) );
  NOR2X1 U229 ( .A(n1140), .B(n672), .Y(n698) );
  NOR2X1 U230 ( .A(n1140), .B(n415), .Y(n475) );
  NOR2BX1 U231 ( .AN(A[0]), .B(n1140), .Y(n899) );
  NOR2X1 U232 ( .A(n1140), .B(n528), .Y(n603) );
  NOR2X2 U233 ( .A(n1140), .B(n456), .Y(n510) );
  XNOR2X1 U234 ( .A(n1128), .B(A[13]), .Y(n458) );
  XNOR2X1 U235 ( .A(n910), .B(A[15]), .Y(n518) );
  XNOR2X1 U236 ( .A(n517), .B(n516), .Y(n538) );
  OAI22X1 U237 ( .A0(n1143), .A1(n533), .B0(n11), .B1(n479), .Y(n516) );
  OAI22X1 U238 ( .A0(n10), .A1(n911), .B0(n953), .B1(n868), .Y(n918) );
  OAI22X1 U239 ( .A0(n859), .A1(n858), .B0(n11), .B1(n846), .Y(n872) );
  XNOR2X1 U240 ( .A(n912), .B(A[21]), .Y(n455) );
  OAI22X2 U241 ( .A0(n1143), .A1(n458), .B0(n11), .B1(n420), .Y(n460) );
  ADDFX2 U242 ( .A(n872), .B(n871), .CI(n870), .CO(n892), .S(n934) );
  OAI22X1 U243 ( .A0(n732), .A1(n478), .B0(n964), .B1(n455), .Y(n511) );
  OAI22X1 U244 ( .A0(n8), .A1(n937), .B0(n12), .B1(n867), .Y(n919) );
  XNOR2X1 U245 ( .A(n936), .B(A[12]), .Y(n867) );
  NAND2X1 U246 ( .A(n838), .B(n72), .Y(n60) );
  NAND3X1 U247 ( .A(n974), .B(n839), .C(n72), .Y(n61) );
  NAND2X1 U248 ( .A(n81), .B(n74), .Y(n68) );
  XNOR2XL U249 ( .A(n856), .B(A[16]), .Y(n857) );
  XNOR2XL U250 ( .A(n893), .B(A[9]), .Y(n186) );
  CLKINVX2 U251 ( .A(n513), .Y(n856) );
  NAND2XL U252 ( .A(n1151), .B(n1153), .Y(n1156) );
  AOI21XL U253 ( .A0(n1196), .A1(n1168), .B0(n1167), .Y(n1169) );
  INVXL U254 ( .A(n1247), .Y(n1167) );
  NOR2X1 U255 ( .A(n584), .B(n1264), .Y(n81) );
  NAND2XL U256 ( .A(n1294), .B(n1295), .Y(n586) );
  NAND2X1 U257 ( .A(n1292), .B(n1293), .Y(n580) );
  NAND2XL U258 ( .A(n504), .B(n1261), .Y(n505) );
  INVXL U259 ( .A(n1260), .Y(n504) );
  NAND2XL U260 ( .A(n1168), .B(n1247), .Y(n1161) );
  XNOR2XL U261 ( .A(n893), .B(A[12]), .Y(n228) );
  BUFX3 U262 ( .A(A[7]), .Y(n860) );
  INVX1 U263 ( .A(B[10]), .Y(n54) );
  XNOR2XL U264 ( .A(n1113), .B(A[17]), .Y(n346) );
  XNOR2XL U265 ( .A(n1113), .B(A[16]), .Y(n377) );
  AOI21X1 U266 ( .A0(n401), .A1(n76), .B0(n75), .Y(n1232) );
  NOR2XL U267 ( .A(n1156), .B(n1252), .Y(n1224) );
  NOR2XL U268 ( .A(n1223), .B(n1240), .Y(n1228) );
  AOI21XL U269 ( .A0(n1196), .A1(n1189), .B0(n1193), .Y(n1180) );
  OAI21XL U270 ( .A0(n802), .A1(n591), .B0(n590), .Y(n594) );
  XNOR2X1 U271 ( .A(n407), .B(n406), .Y(PRODUCT[32]) );
  OAI21XL U272 ( .A0(n1236), .A1(n404), .B0(n403), .Y(n407) );
  XNOR2XL U273 ( .A(n1113), .B(A[21]), .Y(n306) );
  ADDFX2 U274 ( .A(n239), .B(n238), .CI(n237), .CO(n263), .S(n270) );
  OAI22X1 U275 ( .A0(n951), .A1(n187), .B0(n949), .B1(n250), .Y(n238) );
  OAI22XL U276 ( .A0(n8), .A1(n196), .B0(n12), .B1(n233), .Y(n239) );
  XOR2X1 U277 ( .A(B[7]), .B(B[6]), .Y(n40) );
  XNOR2XL U278 ( .A(n893), .B(A[4]), .Y(n122) );
  INVX4 U279 ( .A(n98), .Y(n936) );
  BUFX3 U280 ( .A(n783), .Y(n956) );
  XNOR2XL U281 ( .A(n1113), .B(A[24]), .Y(n1129) );
  INVXL U282 ( .A(n1119), .Y(n1120) );
  XNOR2XL U283 ( .A(n1113), .B(A[23]), .Y(n1114) );
  OAI22XL U284 ( .A0(n1143), .A1(n1129), .B0(n11), .B1(n1141), .Y(n1146) );
  NOR2XL U285 ( .A(n121), .B(n120), .Y(n1218) );
  AOI21XL U286 ( .A0(n1203), .A1(n1204), .B0(n115), .Y(n1221) );
  INVXL U287 ( .A(n1202), .Y(n115) );
  NAND2XL U288 ( .A(n121), .B(n120), .Y(n1219) );
  NAND2XL U289 ( .A(n130), .B(n129), .Y(n1210) );
  INVXL U290 ( .A(n1246), .Y(n1168) );
  XNOR2XL U291 ( .A(n856), .B(A[15]), .Y(n894) );
  NAND2BXL U292 ( .AN(A[0]), .B(n225), .Y(n226) );
  XNOR2XL U293 ( .A(n893), .B(A[13]), .Y(n941) );
  XNOR2XL U294 ( .A(n856), .B(A[18]), .Y(n777) );
  XNOR2XL U295 ( .A(n856), .B(A[19]), .Y(n741) );
  INVXL U296 ( .A(n1251), .Y(n1154) );
  NAND2XL U297 ( .A(n1190), .B(n1168), .Y(n1170) );
  INVXL U298 ( .A(n1244), .Y(n1171) );
  NOR2XL U299 ( .A(n1246), .B(n1244), .Y(n1189) );
  AOI21XL U300 ( .A0(n589), .A1(n81), .B0(n83), .Y(n577) );
  INVXL U301 ( .A(n579), .Y(n581) );
  INVXL U302 ( .A(n1256), .Y(n442) );
  INVXL U303 ( .A(n1258), .Y(n470) );
  AOI21XL U304 ( .A0(n337), .A1(n1151), .B0(n1154), .Y(n77) );
  INVX1 U305 ( .A(B[15]), .Y(n896) );
  OAI22XL U306 ( .A0(n942), .A1(n857), .B0(n816), .B1(n1071), .Y(n852) );
  NAND2BXL U307 ( .AN(A[0]), .B(B[16]), .Y(n817) );
  OAI22XL U308 ( .A0(n732), .A1(n965), .B0(n964), .B1(n963), .Y(n1011) );
  OAI22XL U309 ( .A0(n942), .A1(n186), .B0(n185), .B1(n1071), .Y(n193) );
  OAI22XL U310 ( .A0(n951), .A1(n188), .B0(n949), .B1(n187), .Y(n192) );
  OAI22XL U311 ( .A0(n7), .A1(n245), .B0(n1121), .B1(n944), .Y(n1008) );
  ADDFX2 U312 ( .A(n992), .B(n991), .CI(n990), .CO(n1023), .S(n1029) );
  OAI22X1 U313 ( .A0(n9), .A1(n247), .B0(n956), .B1(n957), .Y(n991) );
  OAI22XL U314 ( .A0(n951), .A1(n249), .B0(n949), .B1(n950), .Y(n992) );
  OAI22XL U315 ( .A0(n9), .A1(n202), .B0(n956), .B1(n232), .Y(n234) );
  OAI22X1 U316 ( .A0(n10), .A1(n201), .B0(n953), .B1(n230), .Y(n235) );
  XNOR2XL U317 ( .A(n856), .B(A[24]), .Y(n527) );
  XNOR2XL U318 ( .A(n856), .B(A[22]), .Y(n634) );
  XNOR2XL U319 ( .A(n856), .B(A[20]), .Y(n700) );
  XNOR2X1 U320 ( .A(n910), .B(A[10]), .Y(n705) );
  XNOR2X1 U321 ( .A(n910), .B(A[13]), .Y(n607) );
  XNOR2XL U322 ( .A(n1138), .B(A[18]), .Y(n287) );
  XNOR2XL U323 ( .A(n1113), .B(A[19]), .Y(n294) );
  XNOR2XL U324 ( .A(n1113), .B(A[18]), .Y(n325) );
  XNOR2XL U325 ( .A(n908), .B(A[25]), .Y(n417) );
  XNOR2XL U326 ( .A(n1113), .B(A[15]), .Y(n385) );
  XNOR2XL U327 ( .A(n893), .B(A[5]), .Y(n94) );
  XNOR2XL U328 ( .A(n893), .B(A[6]), .Y(n87) );
  XNOR2XL U329 ( .A(n893), .B(n860), .Y(n158) );
  NAND2XL U330 ( .A(n1190), .B(n1189), .Y(n1181) );
  INVXL U331 ( .A(n1229), .Y(n1157) );
  INVXL U332 ( .A(n1223), .Y(n1195) );
  XNOR2X1 U333 ( .A(n974), .B(n973), .Y(PRODUCT[17]) );
  NAND2XL U334 ( .A(n926), .B(n1280), .Y(n973) );
  NAND2XL U335 ( .A(n660), .B(n1267), .Y(n661) );
  OAI22XL U336 ( .A0(n9), .A1(n198), .B0(n956), .B1(n202), .Y(n203) );
  XNOR2XL U337 ( .A(n1138), .B(A[20]), .Y(n302) );
  XNOR2XL U338 ( .A(n1113), .B(A[20]), .Y(n291) );
  NAND2BXL U339 ( .AN(A[0]), .B(n910), .Y(n182) );
  OAI22X1 U340 ( .A0(n951), .A1(n250), .B0(n949), .B1(n249), .Y(n258) );
  OAI22X1 U341 ( .A0(n10), .A1(n230), .B0(n953), .B1(n246), .Y(n253) );
  NOR2BX1 U342 ( .AN(A[0]), .B(n1121), .Y(n255) );
  OAI22X1 U343 ( .A0(n9), .A1(n485), .B0(n956), .B1(n417), .Y(n474) );
  XNOR2X1 U344 ( .A(n912), .B(A[19]), .Y(n532) );
  XNOR2X1 U345 ( .A(n912), .B(A[17]), .Y(n625) );
  INVXL U346 ( .A(A[8]), .Y(n70) );
  XNOR2X1 U347 ( .A(n912), .B(A[16]), .Y(n663) );
  XNOR2X1 U348 ( .A(n912), .B(A[15]), .Y(n691) );
  INVXL U349 ( .A(n319), .Y(n320) );
  OAI22XL U350 ( .A0(n10), .A1(n379), .B0(n484), .B1(n347), .Y(n370) );
  CMPR32X1 U351 ( .A(n375), .B(n374), .C(n373), .CO(n355), .S(n408) );
  INVXL U352 ( .A(n352), .Y(n373) );
  OAI22XL U353 ( .A0(n951), .A1(n378), .B0(n949), .B1(n344), .Y(n374) );
  OAI22XL U354 ( .A0(n7), .A1(n380), .B0(n1121), .B1(n343), .Y(n375) );
  AOI21XL U355 ( .A0(n1229), .A1(n1228), .B0(n1227), .Y(n1230) );
  NAND2XL U356 ( .A(n1224), .B(n1228), .Y(n1231) );
  AOI21XL U357 ( .A0(n1196), .A1(n1195), .B0(n1194), .Y(n1197) );
  INVXL U358 ( .A(n1226), .Y(n1194) );
  NAND2XL U359 ( .A(n1190), .B(n1195), .Y(n1198) );
  INVXL U360 ( .A(n1240), .Y(n1199) );
  NOR2X1 U361 ( .A(n68), .B(n280), .Y(n66) );
  NAND2BXL U362 ( .AN(n168), .B(n44), .Y(n42) );
  NAND2BXL U363 ( .AN(n44), .B(n168), .Y(n41) );
  OAI22XL U364 ( .A0(n7), .A1(n305), .B0(n1121), .B1(n1104), .Y(n1107) );
  OAI22XL U365 ( .A0(n1143), .A1(n306), .B0(n11), .B1(n1102), .Y(n1106) );
  INVXL U366 ( .A(n1132), .Y(n1115) );
  OAI22XL U367 ( .A0(n1143), .A1(n1102), .B0(n11), .B1(n1114), .Y(n1117) );
  OAI22XL U368 ( .A0(n9), .A1(n416), .B0(n783), .B1(n119), .Y(n120) );
  NAND2BXL U369 ( .AN(A[0]), .B(n908), .Y(n119) );
  OAI22XL U370 ( .A0(n9), .A1(n125), .B0(n956), .B1(n124), .Y(n135) );
  NOR2BXL U371 ( .AN(A[0]), .B(n12), .Y(n137) );
  OAI22XL U372 ( .A0(n9), .A1(n124), .B0(n956), .B1(n105), .Y(n134) );
  CMPR32X1 U373 ( .A(n104), .B(n103), .C(n102), .CO(n142), .S(n141) );
  OAI22XL U374 ( .A0(n9), .A1(n105), .B0(n956), .B1(n93), .Y(n104) );
  INVXL U375 ( .A(n1141), .Y(n1142) );
  NOR2XL U376 ( .A(n1140), .B(n1139), .Y(n1145) );
  XNOR2XL U377 ( .A(n1138), .B(A[24]), .Y(n1139) );
  INVXL U378 ( .A(n1146), .Y(n1136) );
  XNOR2XL U379 ( .A(n1138), .B(A[23]), .Y(n1127) );
  OAI22XL U380 ( .A0(n942), .A1(A[0]), .B0(n110), .B1(n1071), .Y(n1207) );
  NAND2XL U381 ( .A(n112), .B(n942), .Y(n1206) );
  NAND2BXL U382 ( .AN(A[0]), .B(n893), .Y(n112) );
  NAND2XL U383 ( .A(n1207), .B(n1206), .Y(n1208) );
  INVXL U384 ( .A(n1208), .Y(n1204) );
  INVXL U385 ( .A(n1210), .Y(n131) );
  NAND2XL U386 ( .A(n139), .B(n138), .Y(n1214) );
  INVXL U387 ( .A(n1174), .Y(n1187) );
  INVXL U388 ( .A(n1190), .Y(n1160) );
  INVXL U389 ( .A(n1196), .Y(n1159) );
  XNOR2XL U390 ( .A(n856), .B(A[17]), .Y(n816) );
  XNOR2XL U391 ( .A(n225), .B(A[0]), .Y(n245) );
  INVXL U392 ( .A(n1224), .Y(n1158) );
  NAND2XL U393 ( .A(n1189), .B(n1192), .Y(n1223) );
  INVXL U394 ( .A(n1277), .Y(n927) );
  INVXL U395 ( .A(n1269), .Y(n761) );
  INVX1 U396 ( .A(n1286), .Y(n725) );
  INVXL U397 ( .A(n1266), .Y(n660) );
  AOI21XL U398 ( .A0(n589), .A1(n588), .B0(n587), .Y(n590) );
  INVXL U399 ( .A(n1264), .Y(n592) );
  OAI21XL U400 ( .A0(n65), .A1(n589), .B0(n64), .Y(n63) );
  NOR2XL U401 ( .A(n575), .B(n579), .Y(n64) );
  NOR2BX1 U402 ( .AN(n585), .B(n802), .Y(n65) );
  OAI21XL U403 ( .A0(n576), .A1(n579), .B0(n580), .Y(n84) );
  INVXL U404 ( .A(n83), .Y(n576) );
  INVXL U405 ( .A(n1262), .Y(n85) );
  INVXL U406 ( .A(n439), .Y(n441) );
  INVXL U407 ( .A(n1252), .Y(n363) );
  NAND2XL U408 ( .A(n439), .B(n442), .Y(n404) );
  AOI21XL U409 ( .A0(n401), .A1(n442), .B0(n402), .Y(n403) );
  INVXL U410 ( .A(n1254), .Y(n405) );
  XNOR2XL U411 ( .A(n900), .B(A[0]), .Y(n147) );
  XNOR2XL U412 ( .A(n900), .B(A[1]), .Y(n188) );
  XNOR2XL U413 ( .A(n912), .B(A[4]), .Y(n199) );
  XNOR2XL U414 ( .A(n912), .B(A[12]), .Y(n813) );
  XNOR2XL U415 ( .A(n781), .B(A[16]), .Y(n782) );
  OAI22XL U416 ( .A0(n8), .A1(n867), .B0(n12), .B1(n823), .Y(n864) );
  XNOR2XL U417 ( .A(n908), .B(A[14]), .Y(n862) );
  XNOR2XL U418 ( .A(n225), .B(A[3]), .Y(n904) );
  XNOR2X1 U419 ( .A(n908), .B(A[13]), .Y(n909) );
  XNOR2XL U420 ( .A(n912), .B(A[9]), .Y(n913) );
  XNOR2XL U421 ( .A(n936), .B(A[10]), .Y(n961) );
  OAI22XL U422 ( .A0(n942), .A1(n941), .B0(n940), .B1(n1071), .Y(n988) );
  XNOR2XL U423 ( .A(n936), .B(A[11]), .Y(n937) );
  NAND2BXL U424 ( .AN(A[0]), .B(n1128), .Y(n895) );
  OAI22XL U425 ( .A0(n9), .A1(n957), .B0(n956), .B1(n955), .Y(n993) );
  OAI22X1 U426 ( .A0(n807), .A1(n156), .B0(n155), .B1(n154), .Y(n183) );
  NAND2BXL U427 ( .AN(A[0]), .B(n900), .Y(n154) );
  XNOR2XL U428 ( .A(n900), .B(A[2]), .Y(n187) );
  XNOR2XL U429 ( .A(n893), .B(A[10]), .Y(n185) );
  XNOR2XL U430 ( .A(n893), .B(A[11]), .Y(n229) );
  XNOR2XL U431 ( .A(n910), .B(A[1]), .Y(n230) );
  OAI22XL U432 ( .A0(n942), .A1(n228), .B0(n941), .B1(n1071), .Y(n967) );
  OAI22XL U433 ( .A0(n7), .A1(n286), .B0(n1121), .B1(n226), .Y(n966) );
  INVXL U434 ( .A(n225), .Y(n286) );
  OAI22XL U435 ( .A0(n8), .A1(n233), .B0(n12), .B1(n248), .Y(n240) );
  OAI22XL U436 ( .A0(n732), .A1(n231), .B0(n964), .B1(n243), .Y(n242) );
  XNOR2XL U437 ( .A(n856), .B(A[23]), .Y(n605) );
  XNOR2X1 U438 ( .A(n910), .B(A[14]), .Y(n555) );
  XNOR2XL U439 ( .A(n781), .B(A[22]), .Y(n556) );
  XNOR2XL U440 ( .A(n707), .B(A[20]), .Y(n557) );
  XNOR2XL U441 ( .A(n225), .B(n860), .Y(n769) );
  XNOR2XL U442 ( .A(n900), .B(A[11]), .Y(n773) );
  XNOR2XL U443 ( .A(n900), .B(A[12]), .Y(n738) );
  NOR2X1 U444 ( .A(n1140), .B(n742), .Y(n774) );
  NOR2X1 U445 ( .A(n1140), .B(n701), .Y(n739) );
  ADDFX2 U446 ( .A(n748), .B(n747), .CI(n746), .CO(n757), .S(n794) );
  OAI22XL U447 ( .A0(n9), .A1(n744), .B0(n956), .B1(n706), .Y(n747) );
  OAI22XL U448 ( .A0(n8), .A1(n745), .B0(n12), .B1(n708), .Y(n746) );
  XNOR2XL U449 ( .A(n912), .B(A[25]), .Y(n319) );
  XNOR2XL U450 ( .A(n1138), .B(A[16]), .Y(n317) );
  XNOR2XL U451 ( .A(n912), .B(A[22]), .Y(n421) );
  CMPR32X1 U452 ( .A(n464), .B(n463), .C(n462), .CO(n467), .S(n493) );
  OAI22XL U453 ( .A0(n951), .A1(n476), .B0(n949), .B1(n422), .Y(n464) );
  XNOR2XL U454 ( .A(n601), .B(A[20]), .Y(n422) );
  XNOR2XL U455 ( .A(n1138), .B(A[15]), .Y(n345) );
  OAI22XL U456 ( .A0(n7), .A1(n423), .B0(n1121), .B1(n381), .Y(n427) );
  XNOR2XL U457 ( .A(n912), .B(A[0]), .Y(n91) );
  XNOR2XL U458 ( .A(n912), .B(A[2]), .Y(n159) );
  XNOR2XL U459 ( .A(n893), .B(A[8]), .Y(n157) );
  XNOR2XL U460 ( .A(n936), .B(A[3]), .Y(n150) );
  XOR2XL U461 ( .A(n98), .B(A[4]), .Y(n149) );
  XNOR2X1 U462 ( .A(n908), .B(A[5]), .Y(n148) );
  XNOR2XL U463 ( .A(n908), .B(A[6]), .Y(n153) );
  AOI21XL U464 ( .A0(n1154), .A1(n1153), .B0(n1152), .Y(n1155) );
  INVXL U465 ( .A(n1249), .Y(n1152) );
  NAND2XL U466 ( .A(n1171), .B(n1245), .Y(n1172) );
  AOI21XL U467 ( .A0(n1193), .A1(n1192), .B0(n1191), .Y(n1226) );
  INVXL U468 ( .A(n1243), .Y(n1191) );
  XNOR2X1 U469 ( .A(n583), .B(n582), .Y(PRODUCT[27]) );
  OAI21XL U470 ( .A0(n802), .A1(n578), .B0(n577), .Y(n583) );
  NAND2XL U471 ( .A(n1151), .B(n1251), .Y(n340) );
  NAND2XL U472 ( .A(n1153), .B(n1249), .Y(n79) );
  OAI21XL U473 ( .A0(n1236), .A1(n78), .B0(n77), .Y(n80) );
  XNOR2XL U474 ( .A(n1138), .B(A[22]), .Y(n1118) );
  XNOR2XL U475 ( .A(n225), .B(A[24]), .Y(n1104) );
  XNOR2XL U476 ( .A(n1113), .B(A[22]), .Y(n1102) );
  XNOR2XL U477 ( .A(n1138), .B(A[21]), .Y(n1103) );
  XNOR2XL U478 ( .A(n225), .B(A[23]), .Y(n305) );
  ADDFX2 U479 ( .A(n826), .B(n825), .CI(n824), .CO(n832), .S(n877) );
  OAI22X1 U480 ( .A0(n8), .A1(n823), .B0(n12), .B1(n808), .Y(n825) );
  OAI22XL U481 ( .A0(n807), .A1(n850), .B0(n949), .B1(n806), .Y(n826) );
  OAI22XL U482 ( .A0(n7), .A1(n863), .B0(n1121), .B1(n848), .Y(n870) );
  OAI22XL U483 ( .A0(n732), .A1(n869), .B0(n35), .B1(n849), .Y(n875) );
  ADDFX2 U484 ( .A(n916), .B(n915), .CI(n914), .CO(n906), .S(n979) );
  OAI22X1 U485 ( .A0(n9), .A1(n909), .B0(n956), .B1(n862), .Y(n915) );
  OAI22XL U486 ( .A0(n7), .A1(n904), .B0(n1121), .B1(n863), .Y(n914) );
  OAI22XL U487 ( .A0(n732), .A1(n913), .B0(n35), .B1(n869), .Y(n917) );
  ADDFX2 U488 ( .A(n983), .B(n982), .CI(n981), .CO(n980), .S(n1018) );
  OAI22XL U489 ( .A0(n732), .A1(n963), .B0(n35), .B1(n913), .Y(n981) );
  OAI22XL U490 ( .A0(n9), .A1(n955), .B0(n956), .B1(n909), .Y(n983) );
  OAI22X1 U491 ( .A0(n10), .A1(n952), .B0(n953), .B1(n911), .Y(n982) );
  ADDFX2 U492 ( .A(n986), .B(n985), .CI(n984), .CO(n998), .S(n1017) );
  OAI22XL U493 ( .A0(n8), .A1(n961), .B0(n12), .B1(n937), .Y(n986) );
  NAND2XL U494 ( .A(n257), .B(n258), .Y(n49) );
  NAND2X1 U495 ( .A(n51), .B(n256), .Y(n50) );
  XNOR2XL U496 ( .A(n781), .B(A[23]), .Y(n519) );
  INVXL U497 ( .A(n514), .Y(n486) );
  XNOR2XL U498 ( .A(n601), .B(A[19]), .Y(n476) );
  OAI22XL U499 ( .A0(n7), .A1(n534), .B0(n1121), .B1(n508), .Y(n535) );
  OAI22XL U500 ( .A0(n8), .A1(n520), .B0(n12), .B1(n506), .Y(n537) );
  CMPR32X1 U501 ( .A(n560), .B(n559), .C(n558), .CO(n566), .S(n620) );
  OAI22XL U502 ( .A0(n8), .A1(n557), .B0(n12), .B1(n520), .Y(n558) );
  OAI22XL U503 ( .A0(n9), .A1(n556), .B0(n956), .B1(n519), .Y(n559) );
  OAI22X1 U504 ( .A0(n10), .A1(n555), .B0(n953), .B1(n518), .Y(n560) );
  XNOR2XL U505 ( .A(n900), .B(A[14]), .Y(n668) );
  XNOR2XL U506 ( .A(n900), .B(A[13]), .Y(n697) );
  OAI22XL U507 ( .A0(n942), .A1(n671), .B0(n634), .B1(n1071), .Y(n670) );
  OAI22XL U508 ( .A0(n8), .A1(n708), .B0(n12), .B1(n675), .Y(n709) );
  OAI22XL U509 ( .A0(n8), .A1(n638), .B0(n12), .B1(n609), .Y(n639) );
  OAI22X1 U510 ( .A0(n732), .A1(n731), .B0(n964), .B1(n691), .Y(n737) );
  OAI2BB1XL U511 ( .A0N(n949), .A1N(n951), .B0(n290), .Y(n296) );
  INVXL U512 ( .A(n289), .Y(n290) );
  OAI22XL U513 ( .A0(n10), .A1(n295), .B0(n484), .B1(n293), .Y(n299) );
  OAI22XL U514 ( .A0(n1143), .A1(n294), .B0(n11), .B1(n291), .Y(n301) );
  OAI22XL U515 ( .A0(n7), .A1(n315), .B0(n1121), .B1(n292), .Y(n300) );
  INVXL U516 ( .A(n297), .Y(n327) );
  OAI22XL U517 ( .A0(n1143), .A1(n325), .B0(n11), .B1(n294), .Y(n329) );
  OAI22XL U518 ( .A0(n951), .A1(n344), .B0(n949), .B1(n324), .Y(n350) );
  OAI22XL U519 ( .A0(n7), .A1(n343), .B0(n1121), .B1(n326), .Y(n348) );
  OAI22XL U520 ( .A0(n1143), .A1(n346), .B0(n11), .B1(n325), .Y(n349) );
  OAI2BB1XL U521 ( .A0N(n956), .A1N(n9), .B0(n418), .Y(n473) );
  INVXL U522 ( .A(n417), .Y(n418) );
  ADDFX2 U523 ( .A(n495), .B(n494), .CI(n493), .CO(n481), .S(n542) );
  OAI2BB1XL U524 ( .A0N(n12), .A1N(n8), .B0(n369), .Y(n387) );
  INVXL U525 ( .A(n368), .Y(n369) );
  OAI22XL U526 ( .A0(n951), .A1(n414), .B0(n949), .B1(n378), .Y(n390) );
  OAI22XL U527 ( .A0(n1143), .A1(n385), .B0(n11), .B1(n377), .Y(n391) );
  INVX1 U528 ( .A(B[1]), .Y(n513) );
  XNOR2XL U529 ( .A(n893), .B(A[2]), .Y(n116) );
  CLKINVX4 U530 ( .A(n416), .Y(n908) );
  XNOR2XL U531 ( .A(n908), .B(A[2]), .Y(n124) );
  XNOR2X1 U532 ( .A(n908), .B(A[3]), .Y(n105) );
  OAI22X1 U533 ( .A0(n8), .A1(n98), .B0(n12), .B1(n97), .Y(n108) );
  NAND2BXL U534 ( .AN(A[0]), .B(n936), .Y(n97) );
  OAI22XL U535 ( .A0(n111), .A1(n94), .B0(n87), .B1(n1071), .Y(n100) );
  OAI22XL U536 ( .A0(n8), .A1(n106), .B0(n12), .B1(n92), .Y(n99) );
  NOR2BXL U537 ( .AN(A[0]), .B(n964), .Y(n101) );
  NAND2BXL U538 ( .AN(A[0]), .B(n912), .Y(n86) );
  ADDFX2 U539 ( .A(n163), .B(n162), .CI(n161), .CO(n206), .S(n171) );
  OAI22XL U540 ( .A0(n111), .A1(n158), .B0(n157), .B1(n1071), .Y(n162) );
  OAI22XL U541 ( .A0(n732), .A1(n160), .B0(n964), .B1(n159), .Y(n161) );
  NOR2BXL U542 ( .AN(A[0]), .B(n949), .Y(n163) );
  AOI2BB1X1 U543 ( .A0N(n150), .A1N(n8), .B0(n45), .Y(n44) );
  NAND2XL U544 ( .A(n1192), .B(n1243), .Y(n1182) );
  OAI2BB1XL U545 ( .A0N(n484), .A1N(n10), .B0(n304), .Y(n1099) );
  INVXL U546 ( .A(n303), .Y(n304) );
  OAI22XL U547 ( .A0(n1143), .A1(n291), .B0(n11), .B1(n306), .Y(n309) );
  INVXL U548 ( .A(n1100), .Y(n307) );
  ADDFX2 U549 ( .A(n312), .B(n311), .CI(n310), .CO(n1096), .S(n334) );
  OAI22XL U550 ( .A0(n7), .A1(n292), .B0(n1121), .B1(n305), .Y(n312) );
  ADDFX2 U551 ( .A(n935), .B(n934), .CI(n933), .CO(n921), .S(n977) );
  ADDFX2 U552 ( .A(n980), .B(n979), .CI(n978), .CO(n968), .S(n1003) );
  XNOR3X2 U553 ( .A(n258), .B(n256), .C(n52), .Y(n267) );
  INVXL U554 ( .A(n257), .Y(n52) );
  ADDFX2 U555 ( .A(n523), .B(n522), .CI(n521), .CO(n554), .S(n565) );
  OAI2BB1XL U556 ( .A0N(n1071), .A1N(n942), .B0(n486), .Y(n521) );
  OAI22X1 U557 ( .A0(n9), .A1(n519), .B0(n783), .B1(n485), .Y(n522) );
  OAI22XL U558 ( .A0(n10), .A1(n518), .B0(n484), .B1(n483), .Y(n523) );
  OAI22XL U559 ( .A0(n7), .A1(n508), .B0(n1121), .B1(n471), .Y(n489) );
  OAI22XL U560 ( .A0(n732), .A1(n595), .B0(n964), .B1(n532), .Y(n600) );
  OAI22X1 U561 ( .A0(n1143), .A1(n596), .B0(n11), .B1(n533), .Y(n599) );
  OAI22X1 U562 ( .A0(n732), .A1(n663), .B0(n964), .B1(n625), .Y(n667) );
  OAI22X1 U563 ( .A0(n732), .A1(n691), .B0(n964), .B1(n663), .Y(n696) );
  OAI22X1 U564 ( .A0(n1143), .A1(n692), .B0(n11), .B1(n69), .Y(n695) );
  OAI22XL U565 ( .A0(n10), .A1(n347), .B0(n484), .B1(n342), .Y(n356) );
  OAI22XL U566 ( .A0(n7), .A1(n326), .B0(n1121), .B1(n315), .Y(n332) );
  XNOR2XL U567 ( .A(n1138), .B(A[17]), .Y(n316) );
  ADDFX2 U568 ( .A(n359), .B(n358), .CI(n357), .CO(n360), .S(n396) );
  ADDFX2 U569 ( .A(n543), .B(n542), .CI(n541), .CO(n544), .S(n549) );
  ADDFX2 U570 ( .A(n482), .B(n481), .CI(n480), .CO(n499), .S(n545) );
  OAI22XL U571 ( .A0(n942), .A1(n110), .B0(n116), .B1(n1071), .Y(n114) );
  NOR2BXL U572 ( .AN(A[0]), .B(n956), .Y(n113) );
  INVXL U573 ( .A(n1233), .Y(n1234) );
  NAND2XL U574 ( .A(n1199), .B(n1241), .Y(n1200) );
  NAND2X1 U575 ( .A(n56), .B(n55), .Y(n438) );
  OR2X2 U576 ( .A(n444), .B(n445), .Y(n57) );
  OAI22XL U577 ( .A0(n1143), .A1(n1114), .B0(n11), .B1(n1129), .Y(n1126) );
  NOR2X1 U578 ( .A(n1020), .B(n1019), .Y(n1087) );
  ADDFX2 U579 ( .A(n362), .B(n361), .CI(n360), .CO(n1095), .S(n1092) );
  XOR3X2 U580 ( .A(n445), .B(n443), .C(n444), .Y(n469) );
  NAND2XL U581 ( .A(n114), .B(n113), .Y(n1202) );
  NAND2XL U582 ( .A(n1056), .B(n1055), .Y(n1057) );
  NOR2XL U583 ( .A(n1095), .B(n1094), .Y(mult_x_1_n151) );
  OAI21XL U584 ( .A0(n1052), .A1(n1048), .B0(n1049), .Y(n1047) );
  AND2XL U585 ( .A(n1040), .B(n1038), .Y(n36) );
  NAND2XL U586 ( .A(n1150), .B(n1149), .Y(mult_x_1_n58) );
  NAND2XL U587 ( .A(n1148), .B(n1147), .Y(n1149) );
  NOR2XL U588 ( .A(n1134), .B(n1133), .Y(mult_x_1_n109) );
  NAND2XL U589 ( .A(n1134), .B(n1133), .Y(mult_x_1_n110) );
  NOR2XL U590 ( .A(n1123), .B(n1122), .Y(mult_x_1_n120) );
  NAND2XL U591 ( .A(n1123), .B(n1122), .Y(mult_x_1_n121) );
  NOR2XL U592 ( .A(n1109), .B(n1108), .Y(mult_x_1_n129) );
  NAND2XL U593 ( .A(n1109), .B(n1108), .Y(mult_x_1_n130) );
  NOR2XL U594 ( .A(n574), .B(n573), .Y(mult_x_1_n206) );
  NAND2XL U595 ( .A(n574), .B(n573), .Y(mult_x_1_n207) );
  NOR2XL U596 ( .A(n1093), .B(n1092), .Y(mult_x_1_n160) );
  NOR2BXL U597 ( .AN(A[0]), .B(n1071), .Y(n1321) );
  XNOR2XL U598 ( .A(n1205), .B(n1204), .Y(n1319) );
  NAND2XL U599 ( .A(n1203), .B(n1202), .Y(n1205) );
  NAND2XL U600 ( .A(n1220), .B(n1219), .Y(n1222) );
  INVXL U601 ( .A(n1218), .Y(n1220) );
  NAND2XL U602 ( .A(n128), .B(n1210), .Y(n1212) );
  NAND2XL U603 ( .A(n1215), .B(n1214), .Y(n1217) );
  INVXL U604 ( .A(n1213), .Y(n1215) );
  NAND2XL U605 ( .A(n1186), .B(n1185), .Y(n1188) );
  INVXL U606 ( .A(n1184), .Y(n1186) );
  NAND2XL U607 ( .A(n1177), .B(n1176), .Y(n1178) );
  NAND2XL U608 ( .A(n1164), .B(n1163), .Y(n1165) );
  XNOR2X4 U609 ( .A(B[5]), .B(B[6]), .Y(n35) );
  XNOR2X1 U610 ( .A(n936), .B(A[14]), .Y(n808) );
  CMPR22X1 U611 ( .A(n109), .B(n108), .CO(n103), .S(n132) );
  CMPR22X1 U612 ( .A(n526), .B(n525), .CO(n539), .S(n562) );
  OAI22X1 U613 ( .A0(n942), .A1(n157), .B0(n186), .B1(n1071), .Y(n184) );
  OR2X2 U614 ( .A(n257), .B(n258), .Y(n51) );
  CMPR22X1 U615 ( .A(n252), .B(n251), .CO(n257), .S(n237) );
  CMPR22X1 U616 ( .A(n152), .B(n151), .CO(n167), .S(n174) );
  OAI22X1 U617 ( .A0(n732), .A1(n318), .B0(n964), .B1(n86), .Y(n151) );
  OAI22X1 U618 ( .A0(n732), .A1(n376), .B0(n964), .B1(n319), .Y(n352) );
  OAI22X1 U619 ( .A0(n951), .A1(n324), .B0(n949), .B1(n289), .Y(n297) );
  NOR2X1 U620 ( .A(n1256), .B(n1254), .Y(n76) );
  XNOR2XL U621 ( .A(n900), .B(A[4]), .Y(n249) );
  XNOR2XL U622 ( .A(n908), .B(A[8]), .Y(n202) );
  XNOR2XL U623 ( .A(n936), .B(A[8]), .Y(n248) );
  XNOR2XL U624 ( .A(n225), .B(A[8]), .Y(n734) );
  XNOR2X1 U625 ( .A(n910), .B(A[8]), .Y(n779) );
  NAND2X1 U626 ( .A(n1081), .B(n1080), .Y(n1084) );
  AOI21X1 U627 ( .A0(n1042), .A1(n223), .B0(n222), .Y(n1037) );
  NOR2X1 U628 ( .A(n1275), .B(n1273), .Y(n72) );
  NOR2X1 U629 ( .A(n1279), .B(n1277), .Y(n839) );
  NAND2X2 U630 ( .A(n38), .B(n37), .Y(n974) );
  NAND2X1 U631 ( .A(n1281), .B(n1290), .Y(n38) );
  XOR2X1 U632 ( .A(n1041), .B(n36), .Y(n1309) );
  INVX1 U633 ( .A(n177), .Y(n46) );
  NAND2X4 U634 ( .A(n35), .B(n40), .Y(n732) );
  OAI2BB1X1 U635 ( .A0N(n42), .A1N(n167), .B0(n41), .Y(n216) );
  XOR2X1 U636 ( .A(n167), .B(n43), .Y(n169) );
  XNOR2X1 U637 ( .A(n168), .B(n44), .Y(n43) );
  NAND2BX1 U638 ( .AN(n178), .B(n46), .Y(n1056) );
  NOR2X1 U639 ( .A(n143), .B(n142), .Y(n1175) );
  XOR2X1 U640 ( .A(B[15]), .B(B[14]), .Y(n47) );
  NAND2X2 U641 ( .A(n47), .B(n457), .Y(n859) );
  AOI21X1 U642 ( .A0(n83), .A1(n74), .B0(n67), .Y(n48) );
  XNOR2X1 U643 ( .A(B[11]), .B(n54), .Y(n53) );
  XNOR2X1 U644 ( .A(B[15]), .B(B[16]), .Y(n283) );
  XOR2X2 U645 ( .A(n62), .B(n34), .Y(PRODUCT[28]) );
  OAI21XL U646 ( .A0(n580), .A1(n1262), .B0(n1263), .Y(n67) );
  CLKINVX3 U647 ( .A(B[15]), .Y(n384) );
  OAI22X1 U648 ( .A0(n1143), .A1(n69), .B0(n11), .B1(n626), .Y(n666) );
  XOR2X1 U649 ( .A(n1128), .B(n70), .Y(n69) );
  OAI21XL U650 ( .A0(n1088), .A1(n1087), .B0(n1086), .Y(mult_x_1_n291) );
  XNOR2X2 U651 ( .A(B[12]), .B(B[11]), .Y(n227) );
  CMPR22X1 U652 ( .A(n633), .B(n632), .CO(n613), .S(n643) );
  CMPR22X1 U653 ( .A(n815), .B(n814), .CO(n787), .S(n828) );
  NAND2X1 U654 ( .A(n1036), .B(n1035), .Y(n1083) );
  NOR2X1 U655 ( .A(n579), .B(n1262), .Y(n74) );
  OAI22X1 U656 ( .A0(n1143), .A1(n420), .B0(n11), .B1(n385), .Y(n429) );
  OAI21X2 U657 ( .A0(n1277), .A1(n1280), .B0(n1278), .Y(n838) );
  CMPR22X1 U658 ( .A(n939), .B(n938), .CO(n947), .S(n985) );
  CMPR22X1 U659 ( .A(n775), .B(n774), .CO(n749), .S(n788) );
  OAI22X1 U660 ( .A0(n7), .A1(n471), .B0(n1121), .B1(n423), .Y(n463) );
  XNOR2X1 U661 ( .A(n1128), .B(A[3]), .Y(n846) );
  NOR2X1 U662 ( .A(n1140), .B(n778), .Y(n814) );
  CMPR22X1 U663 ( .A(n740), .B(n739), .CO(n712), .S(n750) );
  NOR2X1 U664 ( .A(n1140), .B(n606), .Y(n632) );
  XNOR2X1 U665 ( .A(n1128), .B(A[12]), .Y(n479) );
  XNOR2X1 U666 ( .A(n1128), .B(A[11]), .Y(n533) );
  CMPR22X1 U667 ( .A(n699), .B(n698), .CO(n679), .S(n713) );
  CMPR22X1 U668 ( .A(n604), .B(n603), .CO(n561), .S(n614) );
  OAI22X1 U669 ( .A0(n1143), .A1(n902), .B0(n11), .B1(n858), .Y(n897) );
  XNOR2X1 U670 ( .A(n1128), .B(A[2]), .Y(n858) );
  NAND2X1 U671 ( .A(n439), .B(n76), .Y(n1225) );
  NOR2X1 U672 ( .A(n1260), .B(n1258), .Y(n439) );
  AOI21X1 U673 ( .A0(n974), .A1(n839), .B0(n838), .Y(n886) );
  OAI21XL U674 ( .A0(n1258), .A1(n1261), .B0(n1259), .Y(n401) );
  XNOR2XL U675 ( .A(n893), .B(A[14]), .Y(n940) );
  OAI22X1 U676 ( .A0(n732), .A1(n159), .B0(n964), .B1(n195), .Y(n191) );
  XNOR2XL U677 ( .A(n781), .B(A[15]), .Y(n822) );
  XNOR2XL U678 ( .A(n707), .B(A[18]), .Y(n638) );
  XNOR2XL U679 ( .A(n856), .B(A[21]), .Y(n671) );
  XNOR2XL U680 ( .A(n908), .B(A[4]), .Y(n93) );
  XNOR2XL U681 ( .A(n893), .B(A[1]), .Y(n110) );
  NOR2X1 U682 ( .A(n1271), .B(n1269), .Y(n656) );
  NAND2X1 U683 ( .A(n656), .B(n73), .Y(n280) );
  NOR2X2 U684 ( .A(n1292), .B(n1293), .Y(n579) );
  OAI21XL U685 ( .A0(n1273), .A1(n1276), .B0(n1274), .Y(n71) );
  NOR2XL U686 ( .A(n1225), .B(n1252), .Y(n336) );
  NAND2XL U687 ( .A(n336), .B(n1151), .Y(n78) );
  OAI21XL U688 ( .A0(n1254), .A1(n1257), .B0(n1255), .Y(n75) );
  OAI21XL U689 ( .A0(n1232), .A1(n1252), .B0(n1253), .Y(n337) );
  INVXL U690 ( .A(n81), .Y(n575) );
  INVX1 U691 ( .A(B[0]), .Y(n776) );
  NAND2XL U692 ( .A(B[1]), .B(n776), .Y(n111) );
  CLKINVX3 U693 ( .A(n513), .Y(n893) );
  BUFX3 U694 ( .A(n776), .Y(n1071) );
  OAI22X1 U695 ( .A0(n942), .A1(n87), .B0(n158), .B1(n1071), .Y(n152) );
  INVX8 U696 ( .A(n318), .Y(n912) );
  XOR2X1 U697 ( .A(B[4]), .B(B[5]), .Y(n88) );
  XNOR2X1 U698 ( .A(B[4]), .B(B[3]), .Y(n96) );
  XNOR2XL U699 ( .A(n936), .B(A[1]), .Y(n106) );
  XOR2X1 U700 ( .A(B[2]), .B(B[3]), .Y(n89) );
  XNOR2X1 U701 ( .A(B[2]), .B(B[1]), .Y(n783) );
  BUFX3 U702 ( .A(B[3]), .Y(n90) );
  INVX4 U703 ( .A(n90), .Y(n416) );
  OAI22X1 U704 ( .A0(n9), .A1(n93), .B0(n956), .B1(n148), .Y(n166) );
  XNOR2X1 U705 ( .A(n912), .B(A[1]), .Y(n160) );
  OAI22X1 U706 ( .A0(n732), .A1(n91), .B0(n964), .B1(n160), .Y(n165) );
  OAI22XL U707 ( .A0(n8), .A1(n92), .B0(n12), .B1(n150), .Y(n164) );
  OAI22X1 U708 ( .A0(n942), .A1(n122), .B0(n94), .B1(n1071), .Y(n109) );
  CMPR32X1 U709 ( .A(n101), .B(n100), .C(n99), .CO(n173), .S(n102) );
  XNOR2X1 U710 ( .A(n936), .B(A[0]), .Y(n107) );
  OAI22XL U711 ( .A0(n8), .A1(n107), .B0(n12), .B1(n106), .Y(n133) );
  NOR2XL U712 ( .A(n1175), .B(n1184), .Y(n145) );
  BUFX3 U713 ( .A(n111), .Y(n942) );
  XNOR2XL U714 ( .A(n893), .B(A[3]), .Y(n123) );
  OAI22X1 U715 ( .A0(n942), .A1(n116), .B0(n123), .B1(n1071), .Y(n127) );
  XNOR2X1 U716 ( .A(n908), .B(A[0]), .Y(n117) );
  OAI22X1 U717 ( .A0(n9), .A1(n117), .B0(n956), .B1(n125), .Y(n126) );
  OAI21XL U718 ( .A0(n1221), .A1(n1218), .B0(n1219), .Y(n1211) );
  OAI22XL U719 ( .A0(n111), .A1(n123), .B0(n122), .B1(n1071), .Y(n136) );
  CMPR22X1 U720 ( .A(n127), .B(n126), .CO(n129), .S(n121) );
  AOI21XL U721 ( .A0(n1211), .A1(n128), .B0(n131), .Y(n1216) );
  CMPR32X1 U722 ( .A(n134), .B(n133), .C(n132), .CO(n140), .S(n139) );
  CMPR32X1 U723 ( .A(n137), .B(n136), .C(n135), .CO(n138), .S(n130) );
  NOR2XL U724 ( .A(n139), .B(n138), .Y(n1213) );
  OAI21XL U725 ( .A0(n1216), .A1(n1213), .B0(n1214), .Y(n1174) );
  NAND2XL U726 ( .A(n143), .B(n142), .Y(n1176) );
  OAI21XL U727 ( .A0(n1175), .A1(n1185), .B0(n1176), .Y(n144) );
  AOI21XL U728 ( .A0(n145), .A1(n1174), .B0(n144), .Y(n1053) );
  XNOR2X1 U729 ( .A(n912), .B(A[3]), .Y(n195) );
  XOR2X1 U730 ( .A(B[8]), .B(B[9]), .Y(n146) );
  BUFX8 U731 ( .A(n807), .Y(n951) );
  OAI22X1 U732 ( .A0(n951), .A1(n147), .B0(n949), .B1(n188), .Y(n190) );
  XNOR2XL U733 ( .A(n936), .B(A[5]), .Y(n197) );
  OAI22XL U734 ( .A0(n8), .A1(n149), .B0(n12), .B1(n197), .Y(n189) );
  OAI22X1 U735 ( .A0(n9), .A1(n148), .B0(n956), .B1(n153), .Y(n168) );
  XNOR2XL U736 ( .A(n908), .B(n860), .Y(n198) );
  OAI22XL U737 ( .A0(n9), .A1(n153), .B0(n956), .B1(n198), .Y(n208) );
  CMPR32X1 U738 ( .A(n171), .B(n170), .C(n169), .CO(n177), .S(n176) );
  CMPR32X1 U739 ( .A(n174), .B(n173), .C(n172), .CO(n175), .S(n143) );
  OR2X2 U740 ( .A(n176), .B(n175), .Y(n1164) );
  NAND2X1 U741 ( .A(n1056), .B(n1164), .Y(n181) );
  NAND2XL U742 ( .A(n176), .B(n175), .Y(n1163) );
  INVXL U743 ( .A(n1163), .Y(n1054) );
  NAND2XL U744 ( .A(n178), .B(n177), .Y(n1055) );
  INVXL U745 ( .A(n1055), .Y(n179) );
  AOI21XL U746 ( .A0(n1056), .A1(n1054), .B0(n179), .Y(n180) );
  XNOR2XL U747 ( .A(n936), .B(A[6]), .Y(n196) );
  XNOR2XL U748 ( .A(n936), .B(n860), .Y(n233) );
  XNOR2X1 U749 ( .A(n900), .B(A[3]), .Y(n250) );
  OAI22X1 U750 ( .A0(n942), .A1(n185), .B0(n229), .B1(n1071), .Y(n252) );
  INVX8 U751 ( .A(n285), .Y(n910) );
  OAI22X1 U752 ( .A0(n10), .A1(n285), .B0(n953), .B1(n182), .Y(n251) );
  CMPR22X1 U753 ( .A(n184), .B(n183), .CO(n211), .S(n207) );
  CMPR32X1 U754 ( .A(n194), .B(n193), .C(n192), .CO(n261), .S(n210) );
  OAI22X1 U755 ( .A0(n732), .A1(n195), .B0(n35), .B1(n199), .Y(n205) );
  OAI22X2 U756 ( .A0(n8), .A1(n197), .B0(n12), .B1(n196), .Y(n204) );
  XNOR2X1 U757 ( .A(n912), .B(A[5]), .Y(n231) );
  OAI22X1 U758 ( .A0(n732), .A1(n199), .B0(n35), .B1(n231), .Y(n236) );
  XNOR2XL U759 ( .A(n910), .B(A[0]), .Y(n201) );
  XNOR2XL U760 ( .A(n908), .B(A[9]), .Y(n232) );
  CMPR32X1 U761 ( .A(n208), .B(n207), .C(n206), .CO(n213), .S(n215) );
  ADDFHX1 U762 ( .A(n211), .B(n210), .CI(n209), .CO(n269), .S(n212) );
  CMPR32X1 U763 ( .A(n214), .B(n213), .C(n212), .CO(n220), .S(n219) );
  CMPR32X1 U764 ( .A(n217), .B(n216), .C(n215), .CO(n218), .S(n178) );
  NOR2X1 U765 ( .A(n219), .B(n218), .Y(n1048) );
  NOR2XL U766 ( .A(n1043), .B(n1048), .Y(n223) );
  NAND2XL U767 ( .A(n219), .B(n218), .Y(n1049) );
  OAI21XL U768 ( .A0(n1043), .A1(n1049), .B0(n1044), .Y(n222) );
  XOR2X1 U769 ( .A(B[12]), .B(B[13]), .Y(n224) );
  BUFX3 U770 ( .A(n227), .Y(n1121) );
  OAI22X2 U771 ( .A0(n942), .A1(n229), .B0(n228), .B1(n1071), .Y(n254) );
  XNOR2X1 U772 ( .A(n912), .B(A[6]), .Y(n243) );
  XNOR2X1 U773 ( .A(n908), .B(A[10]), .Y(n247) );
  OAI22XL U774 ( .A0(n9), .A1(n232), .B0(n956), .B1(n247), .Y(n241) );
  CMPR32X1 U775 ( .A(n242), .B(n241), .C(n240), .CO(n1013), .S(n262) );
  XNOR2X1 U776 ( .A(n912), .B(n860), .Y(n965) );
  OAI22XL U777 ( .A0(n732), .A1(n243), .B0(n964), .B1(n965), .Y(n1009) );
  XNOR2X1 U778 ( .A(n225), .B(A[1]), .Y(n944) );
  XNOR2X1 U779 ( .A(n910), .B(A[3]), .Y(n954) );
  OAI22XL U780 ( .A0(n10), .A1(n246), .B0(n953), .B1(n954), .Y(n1007) );
  XNOR2X1 U781 ( .A(n900), .B(A[5]), .Y(n950) );
  XNOR2X1 U782 ( .A(n908), .B(A[11]), .Y(n957) );
  XNOR2XL U783 ( .A(n936), .B(A[9]), .Y(n962) );
  OAI22XL U784 ( .A0(n8), .A1(n248), .B0(n12), .B1(n962), .Y(n990) );
  NOR2XL U785 ( .A(n273), .B(n272), .Y(n271) );
  NAND2X1 U786 ( .A(n5), .B(n1040), .Y(n278) );
  INVXL U787 ( .A(n1082), .Y(n276) );
  AOI21X1 U788 ( .A0(n5), .A1(n1039), .B0(n276), .Y(n277) );
  OAI21X1 U789 ( .A0(n1037), .A1(n278), .B0(n277), .Y(mult_x_1_n309) );
  OAI21XL U790 ( .A0(n802), .A1(n280), .B0(n279), .Y(n282) );
  NAND2XL U791 ( .A(n588), .B(n586), .Y(n281) );
  XNOR2X1 U792 ( .A(n282), .B(n281), .Y(PRODUCT[25]) );
  XNOR2XL U793 ( .A(n1138), .B(A[19]), .Y(n284) );
  XNOR2XL U794 ( .A(n910), .B(A[25]), .Y(n303) );
  OAI22X1 U795 ( .A0(n10), .A1(n293), .B0(n484), .B1(n303), .Y(n1100) );
  XNOR2X1 U796 ( .A(n225), .B(A[22]), .Y(n292) );
  INVX1 U797 ( .A(B[9]), .Y(n288) );
  CLKINVX3 U798 ( .A(n288), .Y(n601) );
  XNOR2XL U799 ( .A(n601), .B(A[24]), .Y(n324) );
  XNOR2X1 U800 ( .A(n900), .B(A[25]), .Y(n289) );
  XNOR2X1 U801 ( .A(n225), .B(A[21]), .Y(n315) );
  XNOR2XL U802 ( .A(n910), .B(A[23]), .Y(n295) );
  OAI22XL U803 ( .A0(n10), .A1(n342), .B0(n484), .B1(n295), .Y(n328) );
  CMPR32X1 U804 ( .A(n298), .B(n297), .C(n296), .CO(n311), .S(n322) );
  CMPR32X1 U805 ( .A(n301), .B(n300), .C(n299), .CO(n310), .S(n321) );
  CMPR32X1 U806 ( .A(n309), .B(n308), .C(n307), .CO(n1105), .S(n335) );
  NOR2XL U807 ( .A(n314), .B(n313), .Y(mult_x_1_n136) );
  NAND2XL U808 ( .A(n314), .B(n313), .Y(mult_x_1_n137) );
  XNOR2X1 U809 ( .A(n225), .B(A[20]), .Y(n326) );
  XNOR2XL U810 ( .A(n912), .B(A[24]), .Y(n376) );
  CMPR32X1 U811 ( .A(n323), .B(n322), .C(n321), .CO(n333), .S(n361) );
  XNOR2X1 U812 ( .A(n225), .B(A[19]), .Y(n343) );
  CMPR32X1 U813 ( .A(n329), .B(n328), .C(n327), .CO(n323), .S(n358) );
  CMPR32X1 U814 ( .A(n332), .B(n331), .C(n330), .CO(n362), .S(n357) );
  CMPR32X1 U815 ( .A(n335), .B(n334), .C(n333), .CO(n314), .S(n1094) );
  NAND2XL U816 ( .A(n1095), .B(n1094), .Y(mult_x_1_n152) );
  INVXL U817 ( .A(n336), .Y(n339) );
  INVXL U818 ( .A(n337), .Y(n338) );
  OAI21XL U819 ( .A0(n1236), .A1(n339), .B0(n338), .Y(n341) );
  XNOR2X1 U820 ( .A(n341), .B(n340), .Y(PRODUCT[34]) );
  XNOR2X1 U821 ( .A(n910), .B(A[21]), .Y(n347) );
  XNOR2XL U822 ( .A(n225), .B(A[18]), .Y(n380) );
  XNOR2X1 U823 ( .A(n601), .B(A[22]), .Y(n378) );
  OAI22XL U824 ( .A0(n1143), .A1(n377), .B0(n11), .B1(n346), .Y(n371) );
  XNOR2XL U825 ( .A(n910), .B(A[20]), .Y(n379) );
  CMPR32X1 U826 ( .A(n350), .B(n349), .C(n348), .CO(n359), .S(n395) );
  CMPR32X1 U827 ( .A(n353), .B(n352), .C(n351), .CO(n330), .S(n394) );
  NAND2XL U828 ( .A(n1093), .B(n1092), .Y(mult_x_1_n161) );
  OAI21XL U829 ( .A0(n1236), .A1(n1225), .B0(n1232), .Y(n365) );
  XNOR2XL U830 ( .A(n1138), .B(A[14]), .Y(n366) );
  XNOR2X1 U831 ( .A(n936), .B(A[25]), .Y(n368) );
  OAI22X1 U832 ( .A0(n8), .A1(n419), .B0(n12), .B1(n368), .Y(n388) );
  CMPR32X1 U833 ( .A(n372), .B(n371), .C(n370), .CO(n354), .S(n409) );
  OAI22XL U834 ( .A0(n732), .A1(n383), .B0(n964), .B1(n376), .Y(n392) );
  XNOR2XL U835 ( .A(n601), .B(A[21]), .Y(n414) );
  XNOR2X1 U836 ( .A(n910), .B(A[19]), .Y(n386) );
  OAI22XL U837 ( .A0(n10), .A1(n386), .B0(n484), .B1(n379), .Y(n413) );
  XNOR2X1 U838 ( .A(n225), .B(A[17]), .Y(n381) );
  OAI22XL U839 ( .A0(n7), .A1(n381), .B0(n1121), .B1(n380), .Y(n412) );
  XNOR2X1 U840 ( .A(n225), .B(A[16]), .Y(n423) );
  XNOR2X1 U841 ( .A(B[16]), .B(A[13]), .Y(n382) );
  INVXL U842 ( .A(n388), .Y(n425) );
  OAI22XL U843 ( .A0(n732), .A1(n421), .B0(n964), .B1(n383), .Y(n430) );
  INVX8 U844 ( .A(n384), .Y(n1128) );
  XNOR2X1 U845 ( .A(n910), .B(A[18]), .Y(n424) );
  OAI22XL U846 ( .A0(n10), .A1(n424), .B0(n484), .B1(n386), .Y(n428) );
  CMPR32X1 U847 ( .A(n389), .B(n388), .C(n387), .CO(n410), .S(n447) );
  CMPR32X1 U848 ( .A(n392), .B(n391), .C(n390), .CO(n433), .S(n446) );
  CMPR32X1 U849 ( .A(n395), .B(n394), .C(n393), .CO(n397), .S(n434) );
  CMPR32X1 U850 ( .A(n398), .B(n397), .C(n396), .CO(n1093), .S(n399) );
  NOR2XL U851 ( .A(n400), .B(n399), .Y(mult_x_1_n169) );
  NAND2XL U852 ( .A(n400), .B(n399), .Y(mult_x_1_n170) );
  INVXL U853 ( .A(n1257), .Y(n402) );
  CMPR32X1 U854 ( .A(n410), .B(n409), .C(n408), .CO(n436), .S(n445) );
  CMPR32X1 U855 ( .A(n413), .B(n412), .C(n411), .CO(n432), .S(n451) );
  OAI22XL U856 ( .A0(n951), .A1(n422), .B0(n949), .B1(n414), .Y(n454) );
  XNOR2XL U857 ( .A(B[16]), .B(A[12]), .Y(n415) );
  CLKINVX3 U858 ( .A(n416), .Y(n781) );
  XNOR2X1 U859 ( .A(n781), .B(A[24]), .Y(n485) );
  XNOR2XL U860 ( .A(n707), .B(A[23]), .Y(n472) );
  OAI22XL U861 ( .A0(n732), .A1(n455), .B0(n964), .B1(n421), .Y(n459) );
  XNOR2X1 U862 ( .A(n225), .B(A[15]), .Y(n471) );
  XNOR2XL U863 ( .A(n910), .B(A[17]), .Y(n477) );
  OAI22XL U864 ( .A0(n10), .A1(n477), .B0(n484), .B1(n424), .Y(n462) );
  CMPR32X1 U865 ( .A(n436), .B(n435), .C(n434), .CO(n400), .S(n437) );
  NOR2XL U866 ( .A(n438), .B(n437), .Y(mult_x_1_n176) );
  NAND2XL U867 ( .A(n438), .B(n437), .Y(mult_x_1_n177) );
  CMPR32X1 U868 ( .A(n448), .B(n447), .C(n446), .CO(n431), .S(n501) );
  CMPR32X1 U869 ( .A(n451), .B(n450), .C(n449), .CO(n444), .S(n500) );
  ADDFHX1 U870 ( .A(n454), .B(n453), .CI(n452), .CO(n450), .S(n482) );
  XNOR2X1 U871 ( .A(n912), .B(A[20]), .Y(n478) );
  XNOR2X1 U872 ( .A(B[16]), .B(A[11]), .Y(n456) );
  OAI22XL U873 ( .A0(n1143), .A1(n479), .B0(n11), .B1(n458), .Y(n509) );
  NOR2XL U874 ( .A(n469), .B(n468), .Y(mult_x_1_n183) );
  NAND2XL U875 ( .A(n469), .B(n468), .Y(mult_x_1_n184) );
  XNOR2X1 U876 ( .A(n707), .B(A[22]), .Y(n506) );
  OAI22XL U877 ( .A0(n8), .A1(n506), .B0(n12), .B1(n472), .Y(n488) );
  INVXL U878 ( .A(n474), .Y(n487) );
  CMPR32X1 U879 ( .A(n475), .B(n474), .C(n473), .CO(n453), .S(n497) );
  XNOR2XL U880 ( .A(n601), .B(A[18]), .Y(n512) );
  OAI22XL U881 ( .A0(n951), .A1(n512), .B0(n949), .B1(n476), .Y(n492) );
  OAI22XL U882 ( .A0(n10), .A1(n483), .B0(n484), .B1(n477), .Y(n491) );
  OAI22XL U883 ( .A0(n732), .A1(n532), .B0(n964), .B1(n478), .Y(n517) );
  OR2X2 U884 ( .A(n517), .B(n516), .Y(n490) );
  XNOR2XL U885 ( .A(n893), .B(A[25]), .Y(n514) );
  CMPR32X1 U886 ( .A(n489), .B(n488), .C(n487), .CO(n498), .S(n553) );
  CMPR32X1 U887 ( .A(n492), .B(n491), .C(n490), .CO(n496), .S(n552) );
  CMPR32X1 U888 ( .A(n498), .B(n497), .C(n496), .CO(n546), .S(n541) );
  CMPR32X1 U889 ( .A(n501), .B(n500), .C(n499), .CO(n468), .S(n502) );
  NOR2XL U890 ( .A(n503), .B(n502), .Y(mult_x_1_n194) );
  NAND2XL U891 ( .A(n503), .B(n502), .Y(mult_x_1_n195) );
  XNOR2X1 U892 ( .A(n707), .B(A[21]), .Y(n520) );
  XNOR2X1 U893 ( .A(B[16]), .B(A[10]), .Y(n507) );
  NOR2XL U894 ( .A(n1140), .B(n507), .Y(n536) );
  XNOR2XL U895 ( .A(n601), .B(A[17]), .Y(n524) );
  OAI22X1 U896 ( .A0(n942), .A1(n527), .B0(n514), .B1(n776), .Y(n526) );
  XNOR2X1 U897 ( .A(B[16]), .B(A[9]), .Y(n515) );
  XNOR2XL U898 ( .A(n601), .B(A[16]), .Y(n602) );
  OAI22XL U899 ( .A0(n951), .A1(n602), .B0(n949), .B1(n524), .Y(n563) );
  OAI22X1 U900 ( .A0(n942), .A1(n605), .B0(n527), .B1(n776), .Y(n604) );
  XNOR2X1 U901 ( .A(n912), .B(A[18]), .Y(n595) );
  XNOR2X1 U902 ( .A(n1128), .B(A[10]), .Y(n596) );
  XNOR2X1 U903 ( .A(n225), .B(A[12]), .Y(n597) );
  OAI22XL U904 ( .A0(n7), .A1(n597), .B0(n1121), .B1(n534), .Y(n598) );
  CMPR32X1 U905 ( .A(n537), .B(n536), .C(n535), .CO(n531), .S(n568) );
  XNOR2X1 U906 ( .A(n781), .B(A[21]), .Y(n608) );
  OAI22XL U907 ( .A0(n9), .A1(n608), .B0(n956), .B1(n556), .Y(n611) );
  XNOR2X1 U908 ( .A(n707), .B(A[19]), .Y(n609) );
  CMPR32X1 U909 ( .A(n563), .B(n561), .C(n562), .CO(n564), .S(n619) );
  CMPR32X1 U910 ( .A(n569), .B(n568), .C(n567), .CO(n570), .S(n622) );
  NAND2XL U911 ( .A(n585), .B(n81), .Y(n578) );
  NAND2XL U912 ( .A(n581), .B(n580), .Y(n582) );
  INVXL U913 ( .A(n584), .Y(n588) );
  NAND2XL U914 ( .A(n585), .B(n588), .Y(n591) );
  INVXL U915 ( .A(n586), .Y(n587) );
  NAND2X1 U916 ( .A(n592), .B(n1265), .Y(n593) );
  OAI22X1 U917 ( .A0(n732), .A1(n625), .B0(n964), .B1(n595), .Y(n630) );
  XNOR2X1 U918 ( .A(n1128), .B(A[9]), .Y(n626) );
  OAI22X1 U919 ( .A0(n1143), .A1(n626), .B0(n11), .B1(n596), .Y(n629) );
  XNOR2X1 U920 ( .A(n225), .B(A[11]), .Y(n627) );
  OAI22XL U921 ( .A0(n7), .A1(n627), .B0(n1121), .B1(n597), .Y(n628) );
  XNOR2XL U922 ( .A(n601), .B(A[15]), .Y(n631) );
  OAI22XL U923 ( .A0(n951), .A1(n631), .B0(n949), .B1(n602), .Y(n615) );
  OAI22X1 U924 ( .A0(n942), .A1(n634), .B0(n605), .B1(n1071), .Y(n633) );
  XNOR2X1 U925 ( .A(B[16]), .B(n860), .Y(n606) );
  XNOR2X1 U926 ( .A(n910), .B(A[12]), .Y(n636) );
  OAI22X1 U927 ( .A0(n10), .A1(n636), .B0(n953), .B1(n607), .Y(n641) );
  OAI22XL U928 ( .A0(n9), .A1(n637), .B0(n956), .B1(n608), .Y(n640) );
  CMPR32X1 U929 ( .A(n612), .B(n611), .C(n610), .CO(n621), .S(n649) );
  CMPR32X1 U930 ( .A(n615), .B(n614), .C(n613), .CO(n616), .S(n648) );
  ADDFHX1 U931 ( .A(n624), .B(n623), .CI(n622), .CO(n1060), .S(n1062) );
  XNOR2X1 U932 ( .A(n225), .B(A[10]), .Y(n664) );
  OAI22XL U933 ( .A0(n7), .A1(n664), .B0(n1121), .B1(n627), .Y(n665) );
  OAI22XL U934 ( .A0(n951), .A1(n668), .B0(n949), .B1(n631), .Y(n644) );
  XNOR2X1 U935 ( .A(B[16]), .B(A[6]), .Y(n635) );
  XNOR2X1 U936 ( .A(n910), .B(A[11]), .Y(n673) );
  OAI22X1 U937 ( .A0(n10), .A1(n673), .B0(n953), .B1(n636), .Y(n678) );
  XNOR2X1 U938 ( .A(n781), .B(A[19]), .Y(n674) );
  OAI22X1 U939 ( .A0(n9), .A1(n674), .B0(n956), .B1(n637), .Y(n677) );
  XNOR2X1 U940 ( .A(n707), .B(A[17]), .Y(n675) );
  CMPR32X1 U941 ( .A(n641), .B(n640), .C(n639), .CO(n650), .S(n686) );
  CMPR32X1 U942 ( .A(n644), .B(n643), .C(n642), .CO(n645), .S(n685) );
  CMPR32X1 U943 ( .A(n647), .B(n646), .C(n645), .CO(n1067), .S(n689) );
  CMPR32X1 U944 ( .A(n650), .B(n649), .C(n648), .CO(n653), .S(n688) );
  CMPR32X1 U945 ( .A(n653), .B(n652), .C(n651), .CO(n1063), .S(n1065) );
  NOR2XL U946 ( .A(n655), .B(n654), .Y(mult_x_1_n226) );
  NAND2XL U947 ( .A(n655), .B(n654), .Y(mult_x_1_n227) );
  NAND2XL U948 ( .A(n656), .B(n725), .Y(n659) );
  AOI21XL U949 ( .A0(n657), .A1(n725), .B0(n22), .Y(n658) );
  OAI21XL U950 ( .A0(n802), .A1(n659), .B0(n658), .Y(n662) );
  XNOR2X1 U951 ( .A(n662), .B(n661), .Y(PRODUCT[24]) );
  XNOR2X1 U952 ( .A(n1128), .B(n860), .Y(n692) );
  XNOR2X1 U953 ( .A(n225), .B(A[9]), .Y(n693) );
  OAI22XL U954 ( .A0(n7), .A1(n693), .B0(n1121), .B1(n664), .Y(n694) );
  OAI22XL U955 ( .A0(n951), .A1(n697), .B0(n949), .B1(n668), .Y(n681) );
  ADDHXL U956 ( .A(n670), .B(n669), .CO(n642), .S(n680) );
  OAI22X1 U957 ( .A0(n942), .A1(n700), .B0(n671), .B1(n1071), .Y(n699) );
  XNOR2X1 U958 ( .A(B[16]), .B(A[5]), .Y(n672) );
  OAI22X1 U959 ( .A0(n10), .A1(n705), .B0(n953), .B1(n673), .Y(n711) );
  XNOR2X1 U960 ( .A(n781), .B(A[18]), .Y(n706) );
  OAI22XL U961 ( .A0(n9), .A1(n706), .B0(n956), .B1(n674), .Y(n710) );
  XNOR2X1 U962 ( .A(n707), .B(A[16]), .Y(n708) );
  CMPR32X1 U963 ( .A(n681), .B(n679), .C(n680), .CO(n682), .S(n718) );
  CMPR32X1 U964 ( .A(n684), .B(n683), .C(n682), .CO(n1070), .S(n703) );
  CMPR32X1 U965 ( .A(n687), .B(n686), .C(n685), .CO(n690), .S(n702) );
  XNOR2X1 U966 ( .A(n912), .B(A[14]), .Y(n731) );
  XNOR2X1 U967 ( .A(n1128), .B(A[6]), .Y(n733) );
  OAI22X1 U968 ( .A0(n1143), .A1(n733), .B0(n11), .B1(n692), .Y(n736) );
  OAI22XL U969 ( .A0(n7), .A1(n734), .B0(n1121), .B1(n693), .Y(n735) );
  OAI22XL U970 ( .A0(n951), .A1(n738), .B0(n949), .B1(n697), .Y(n714) );
  OAI22X1 U971 ( .A0(n942), .A1(n741), .B0(n700), .B1(n776), .Y(n740) );
  XNOR2X1 U972 ( .A(B[16]), .B(A[4]), .Y(n701) );
  XNOR2X1 U973 ( .A(n910), .B(A[9]), .Y(n743) );
  OAI22X1 U974 ( .A0(n10), .A1(n743), .B0(n953), .B1(n705), .Y(n748) );
  XNOR2X1 U975 ( .A(n781), .B(A[17]), .Y(n744) );
  CMPR32X1 U976 ( .A(n711), .B(n710), .C(n709), .CO(n720), .S(n756) );
  CMPR32X1 U977 ( .A(n714), .B(n713), .C(n712), .CO(n715), .S(n755) );
  CMPR32X1 U978 ( .A(n717), .B(n716), .C(n715), .CO(n730), .S(n759) );
  NOR2XL U979 ( .A(n722), .B(n721), .Y(mult_x_1_n244) );
  NAND2XL U980 ( .A(n722), .B(n721), .Y(mult_x_1_n245) );
  INVXL U981 ( .A(n656), .Y(n724) );
  INVXL U982 ( .A(n657), .Y(n723) );
  OAI21XL U983 ( .A0(n802), .A1(n724), .B0(n723), .Y(n727) );
  NAND2X1 U984 ( .A(n725), .B(n1268), .Y(n726) );
  ADDFHX1 U985 ( .A(n730), .B(n729), .CI(n728), .CO(n721), .S(n1073) );
  XNOR2X1 U986 ( .A(n912), .B(A[13]), .Y(n767) );
  OAI22X1 U987 ( .A0(n732), .A1(n767), .B0(n964), .B1(n731), .Y(n772) );
  XNOR2X1 U988 ( .A(n1128), .B(A[5]), .Y(n768) );
  OAI22X1 U989 ( .A0(n1143), .A1(n768), .B0(n11), .B1(n733), .Y(n771) );
  OAI22XL U990 ( .A0(n7), .A1(n769), .B0(n1121), .B1(n734), .Y(n770) );
  OAI22XL U991 ( .A0(n951), .A1(n773), .B0(n949), .B1(n738), .Y(n751) );
  OAI22X1 U992 ( .A0(n942), .A1(n777), .B0(n741), .B1(n1071), .Y(n775) );
  XNOR2X1 U993 ( .A(B[16]), .B(A[3]), .Y(n742) );
  OAI22X1 U994 ( .A0(n10), .A1(n779), .B0(n953), .B1(n743), .Y(n786) );
  OAI22X1 U995 ( .A0(n9), .A1(n782), .B0(n956), .B1(n744), .Y(n785) );
  CMPR32X1 U996 ( .A(n751), .B(n750), .C(n749), .CO(n752), .S(n793) );
  CMPR32X1 U997 ( .A(n754), .B(n753), .C(n752), .CO(n766), .S(n797) );
  CMPR32X1 U998 ( .A(n757), .B(n756), .C(n755), .CO(n760), .S(n796) );
  CMPR32X1 U999 ( .A(n760), .B(n759), .C(n758), .CO(n728), .S(n764) );
  NAND2XL U1000 ( .A(n1073), .B(n1072), .Y(mult_x_1_n252) );
  NAND2X1 U1001 ( .A(n761), .B(n1270), .Y(n762) );
  ADDFHX1 U1002 ( .A(n766), .B(n765), .CI(n764), .CO(n1072), .S(n800) );
  OAI22X1 U1003 ( .A0(n732), .A1(n813), .B0(n35), .B1(n767), .Y(n812) );
  XNOR2X1 U1004 ( .A(n1128), .B(A[4]), .Y(n780) );
  OAI22X1 U1005 ( .A0(n1143), .A1(n780), .B0(n11), .B1(n768), .Y(n811) );
  XNOR2X1 U1006 ( .A(n225), .B(A[6]), .Y(n809) );
  OAI22XL U1007 ( .A0(n7), .A1(n809), .B0(n1121), .B1(n769), .Y(n810) );
  XNOR2X1 U1008 ( .A(n900), .B(A[10]), .Y(n806) );
  OAI22XL U1009 ( .A0(n951), .A1(n806), .B0(n949), .B1(n773), .Y(n789) );
  OAI22X1 U1010 ( .A0(n942), .A1(n816), .B0(n777), .B1(n776), .Y(n815) );
  XNOR2X1 U1011 ( .A(B[16]), .B(A[2]), .Y(n778) );
  XNOR2X1 U1012 ( .A(n910), .B(n860), .Y(n821) );
  OAI22X1 U1013 ( .A0(n10), .A1(n821), .B0(n953), .B1(n779), .Y(n855) );
  OAI22X1 U1014 ( .A0(n859), .A1(n846), .B0(n11), .B1(n780), .Y(n854) );
  OAI22XL U1015 ( .A0(n9), .A1(n822), .B0(n783), .B1(n782), .Y(n853) );
  CMPR32X1 U1016 ( .A(n786), .B(n785), .C(n784), .CO(n795), .S(n834) );
  CMPR32X1 U1017 ( .A(n789), .B(n788), .C(n787), .CO(n790), .S(n833) );
  CMPR32X1 U1018 ( .A(n792), .B(n791), .C(n790), .CO(n805), .S(n819) );
  CMPR32X1 U1019 ( .A(n795), .B(n794), .C(n793), .CO(n798), .S(n818) );
  NOR2XL U1020 ( .A(n800), .B(n799), .Y(mult_x_1_n262) );
  NAND2XL U1021 ( .A(n800), .B(n799), .Y(mult_x_1_n263) );
  NAND2X1 U1022 ( .A(n59), .B(n1272), .Y(n801) );
  XOR2X1 U1023 ( .A(n802), .B(n801), .Y(PRODUCT[21]) );
  ADDFHX1 U1024 ( .A(n805), .B(n804), .CI(n803), .CO(n799), .S(n837) );
  XNOR2X1 U1025 ( .A(n900), .B(A[9]), .Y(n850) );
  XNOR2XL U1026 ( .A(n936), .B(A[13]), .Y(n823) );
  XNOR2X1 U1027 ( .A(n225), .B(A[5]), .Y(n848) );
  OAI22XL U1028 ( .A0(n7), .A1(n848), .B0(n1121), .B1(n809), .Y(n824) );
  XNOR2X1 U1029 ( .A(n912), .B(A[11]), .Y(n849) );
  OAI22XL U1030 ( .A0(n732), .A1(n849), .B0(n35), .B1(n813), .Y(n829) );
  XNOR2X1 U1031 ( .A(n910), .B(A[6]), .Y(n868) );
  OAI22X1 U1032 ( .A0(n10), .A1(n868), .B0(n953), .B1(n821), .Y(n866) );
  OAI22XL U1033 ( .A0(n9), .A1(n862), .B0(n956), .B1(n822), .Y(n865) );
  CMPR32X1 U1034 ( .A(n829), .B(n828), .C(n827), .CO(n830), .S(n876) );
  CMPR32X1 U1035 ( .A(n832), .B(n831), .C(n830), .CO(n845), .S(n880) );
  CMPR32X1 U1036 ( .A(n835), .B(n834), .C(n833), .CO(n820), .S(n879) );
  NOR2XL U1037 ( .A(n837), .B(n836), .Y(mult_x_1_n265) );
  NAND2XL U1038 ( .A(n837), .B(n836), .Y(mult_x_1_n266) );
  OAI21XL U1039 ( .A0(n886), .A1(n1275), .B0(n1276), .Y(n842) );
  INVXL U1040 ( .A(n1273), .Y(n840) );
  NAND2XL U1041 ( .A(n840), .B(n1274), .Y(n841) );
  ADDFHX1 U1042 ( .A(n845), .B(n844), .CI(n843), .CO(n836), .S(n883) );
  XNOR2X1 U1043 ( .A(B[16]), .B(A[1]), .Y(n847) );
  XNOR2X1 U1044 ( .A(n225), .B(A[4]), .Y(n863) );
  XNOR2X1 U1045 ( .A(n912), .B(A[10]), .Y(n869) );
  XNOR2X1 U1046 ( .A(n900), .B(A[8]), .Y(n861) );
  OAI22XL U1047 ( .A0(n951), .A1(n861), .B0(n949), .B1(n850), .Y(n874) );
  ADDHXL U1048 ( .A(n852), .B(n851), .CO(n827), .S(n873) );
  CMPR32X1 U1049 ( .A(n855), .B(n854), .C(n853), .CO(n835), .S(n890) );
  OAI22X2 U1050 ( .A0(n942), .A1(n894), .B0(n857), .B1(n1071), .Y(n898) );
  XNOR2X1 U1051 ( .A(n1128), .B(A[1]), .Y(n902) );
  XNOR2X1 U1052 ( .A(n900), .B(n860), .Y(n901) );
  CMPR32X1 U1053 ( .A(n866), .B(n865), .C(n864), .CO(n878), .S(n905) );
  XNOR2X1 U1054 ( .A(n910), .B(A[5]), .Y(n911) );
  CMPR32X1 U1055 ( .A(n875), .B(n874), .C(n873), .CO(n891), .S(n933) );
  CMPR32X1 U1056 ( .A(n878), .B(n877), .C(n876), .CO(n881), .S(n920) );
  NOR2XL U1057 ( .A(n883), .B(n882), .Y(mult_x_1_n273) );
  NAND2XL U1058 ( .A(n883), .B(n882), .Y(mult_x_1_n274) );
  INVXL U1059 ( .A(n1275), .Y(n884) );
  NAND2XL U1060 ( .A(n884), .B(n1276), .Y(n885) );
  XOR2X1 U1061 ( .A(n886), .B(n885), .Y(PRODUCT[19]) );
  CMPR32X1 U1062 ( .A(n892), .B(n891), .C(n890), .CO(n889), .S(n932) );
  OAI22X1 U1063 ( .A0(n942), .A1(n940), .B0(n894), .B1(n1071), .Y(n939) );
  XNOR2X1 U1064 ( .A(n900), .B(A[6]), .Y(n948) );
  OAI22X1 U1065 ( .A0(n951), .A1(n948), .B0(n949), .B1(n901), .Y(n960) );
  XNOR2XL U1066 ( .A(n1128), .B(A[0]), .Y(n903) );
  OAI22X1 U1067 ( .A0(n1143), .A1(n903), .B0(n11), .B1(n902), .Y(n959) );
  XNOR2X1 U1068 ( .A(n225), .B(A[2]), .Y(n943) );
  OAI22XL U1069 ( .A0(n7), .A1(n943), .B0(n1121), .B1(n904), .Y(n958) );
  XNOR2X1 U1070 ( .A(n908), .B(A[12]), .Y(n955) );
  XNOR2X1 U1071 ( .A(n910), .B(A[4]), .Y(n952) );
  XNOR2X1 U1072 ( .A(n912), .B(A[8]), .Y(n963) );
  INVXL U1073 ( .A(n1280), .Y(n925) );
  AOI21X1 U1074 ( .A0(n974), .A1(n926), .B0(n925), .Y(n929) );
  NAND2XL U1075 ( .A(n927), .B(n1278), .Y(n928) );
  XOR2X1 U1076 ( .A(n929), .B(n928), .Y(PRODUCT[18]) );
  NOR2BX1 U1077 ( .AN(A[0]), .B(n11), .Y(n989) );
  OAI22XL U1078 ( .A0(n7), .A1(n944), .B0(n1121), .B1(n943), .Y(n987) );
  OAI22X1 U1079 ( .A0(n951), .A1(n950), .B0(n949), .B1(n948), .Y(n995) );
  OAI22X1 U1080 ( .A0(n10), .A1(n954), .B0(n953), .B1(n952), .Y(n994) );
  OAI22XL U1081 ( .A0(n8), .A1(n962), .B0(n12), .B1(n961), .Y(n1012) );
  ADDHXL U1082 ( .A(n967), .B(n966), .CO(n1010), .S(n1015) );
  NOR2XL U1083 ( .A(n972), .B(n971), .Y(mult_x_1_n281) );
  CMPR32X1 U1084 ( .A(n977), .B(n976), .C(n975), .CO(n971), .S(n1000) );
  CMPR32X1 U1085 ( .A(n989), .B(n988), .C(n987), .CO(n984), .S(n1024) );
  NOR2XL U1086 ( .A(n1000), .B(n999), .Y(mult_x_1_n286) );
  NAND2XL U1087 ( .A(n1000), .B(n999), .Y(mult_x_1_n287) );
  CMPR32X1 U1088 ( .A(n1006), .B(n1005), .C(n1004), .CO(n996), .S(n1076) );
  CMPR32X1 U1089 ( .A(n1009), .B(n1008), .C(n1007), .CO(n1027), .S(n1030) );
  CMPR32X1 U1090 ( .A(n1012), .B(n1011), .C(n1010), .CO(n1004), .S(n1026) );
  ADDFHX1 U1091 ( .A(n1015), .B(n1014), .CI(n1013), .CO(n1025), .S(n1033) );
  INVXL U1092 ( .A(n1087), .Y(n1021) );
  NAND2XL U1093 ( .A(n1021), .B(n1086), .Y(mult_x_1_n82) );
  XNOR2X1 U1094 ( .A(n1289), .B(n1283), .Y(PRODUCT[15]) );
  XOR2X1 U1095 ( .A(n1238), .B(n1284), .Y(PRODUCT[14]) );
  CMPR32X1 U1096 ( .A(n1030), .B(n1029), .C(n1028), .CO(n1077), .S(n1031) );
  INVXL U1097 ( .A(n1034), .Y(n1090) );
  NAND2XL U1098 ( .A(n1090), .B(n1083), .Y(mult_x_1_n84) );
  INVXL U1099 ( .A(n1037), .Y(n1041) );
  AOI21XL U1100 ( .A0(n1041), .A1(n1040), .B0(n1039), .Y(mult_x_1_n316) );
  INVXL U1101 ( .A(n1042), .Y(n1052) );
  INVXL U1102 ( .A(n1043), .Y(n1045) );
  NAND2XL U1103 ( .A(n1045), .B(n1044), .Y(n1046) );
  XNOR2X1 U1104 ( .A(n1047), .B(n1046), .Y(n1310) );
  INVXL U1105 ( .A(n1048), .Y(n1050) );
  NAND2XL U1106 ( .A(n1050), .B(n1049), .Y(n1051) );
  INVXL U1107 ( .A(n1053), .Y(n1166) );
  AOI21XL U1108 ( .A0(n1166), .A1(n1164), .B0(n1054), .Y(n1058) );
  ADDFHX1 U1109 ( .A(n1061), .B(n1060), .CI(n1059), .CO(n573), .S(
        mult_x_1_n522) );
  ADDFHX1 U1110 ( .A(n1064), .B(n1063), .CI(n1062), .CO(mult_x_1_n537), .S(
        n655) );
  ADDFHX1 U1111 ( .A(n1067), .B(n1066), .CI(n1065), .CO(n654), .S(
        mult_x_1_n554) );
  ADDFHX1 U1112 ( .A(n1070), .B(n1069), .CI(n1068), .CO(mult_x_1_n569), .S(
        n722) );
  NOR2XL U1113 ( .A(n1073), .B(n1072), .Y(mult_x_1_n251) );
  NAND2XL U1114 ( .A(n6), .B(n1084), .Y(mult_x_1_n83) );
  NAND2XL U1115 ( .A(n5), .B(n1082), .Y(mult_x_1_n85) );
  INVXL U1116 ( .A(n1083), .Y(n1091) );
  INVXL U1117 ( .A(n1084), .Y(n1085) );
  NAND2XL U1118 ( .A(n6), .B(n1090), .Y(n1089) );
  NOR2XL U1119 ( .A(n1089), .B(n1087), .Y(mult_x_1_n290) );
  CLKINVX2 U1120 ( .A(mult_x_1_n309), .Y(mult_x_1_n308) );
  OAI21XL U1121 ( .A0(mult_x_1_n308), .A1(n1089), .B0(n1088), .Y(mult_x_1_n294) );
  OAI21XL U1122 ( .A0(mult_x_1_n308), .A1(n1034), .B0(n1083), .Y(mult_x_1_n301) );
  CMPR32X1 U1123 ( .A(n1098), .B(n1097), .C(n1096), .CO(n1109), .S(n313) );
  CMPR32X1 U1124 ( .A(n1101), .B(n1100), .C(n1099), .CO(n1112), .S(n1098) );
  XNOR2XL U1125 ( .A(n225), .B(A[25]), .Y(n1119) );
  OAI22X1 U1126 ( .A0(n7), .A1(n1104), .B0(n1121), .B1(n1119), .Y(n1132) );
  CMPR32X1 U1127 ( .A(n1107), .B(n1106), .C(n1105), .CO(n1110), .S(n1097) );
  CMPR32X1 U1128 ( .A(n1112), .B(n1111), .C(n1110), .CO(n1123), .S(n1108) );
  CMPR32X1 U1129 ( .A(n1117), .B(n1116), .C(n1115), .CO(n1125), .S(n1111) );
  CMPR32X1 U1130 ( .A(n1126), .B(n1125), .C(n1124), .CO(n1134), .S(n1122) );
  XNOR2XL U1131 ( .A(n1128), .B(A[25]), .Y(n1141) );
  CMPR32X1 U1132 ( .A(n1132), .B(n1131), .C(n1130), .CO(n1135), .S(n1124) );
  CMPR32X1 U1133 ( .A(n1137), .B(n1136), .C(n1135), .CO(n1148), .S(n1133) );
  XOR3X2 U1134 ( .A(n1146), .B(n1145), .C(n1144), .Y(n1147) );
  OAI21XL U1135 ( .A0(n1156), .A1(n1253), .B0(n1155), .Y(n1229) );
  OAI21XL U1136 ( .A0(n1236), .A1(n1160), .B0(n1159), .Y(n1162) );
  OAI21XL U1137 ( .A0(n1236), .A1(n1170), .B0(n1169), .Y(n1173) );
  OAI21XL U1138 ( .A0(n1187), .A1(n1184), .B0(n1185), .Y(n1179) );
  INVXL U1139 ( .A(n1175), .Y(n1177) );
  OAI21XL U1140 ( .A0(n1244), .A1(n1247), .B0(n1245), .Y(n1193) );
  OAI21XL U1141 ( .A0(n1236), .A1(n1181), .B0(n1180), .Y(n1183) );
  OAI21XL U1142 ( .A0(n1236), .A1(n1198), .B0(n1197), .Y(n1201) );
  XNOR2XL U1143 ( .A(n1212), .B(n1211), .Y(n1317) );
  XOR2XL U1144 ( .A(n1217), .B(n1216), .Y(n1316) );
  XOR2XL U1145 ( .A(n1222), .B(n1221), .Y(n1318) );
  OAI21XL U1146 ( .A0(n1226), .A1(n1240), .B0(n1241), .Y(n1227) );
  OAI21XL U1147 ( .A0(n1232), .A1(n1231), .B0(n1230), .Y(n1233) );
  OAI21XL U1148 ( .A0(n1236), .A1(n1235), .B0(n1234), .Y(n1237) );
  XNOR2XL U1149 ( .A(n1237), .B(n1239), .Y(PRODUCT[40]) );
endmodule


module FFT2048_DW02_mult_2_stage_J1_5 ( A, B, TC, CLK, PRODUCT );
  input [25:0] A;
  input [16:0] B;
  output [42:0] PRODUCT;
  input TC, CLK;
  wire   n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, mult_x_1_n665, mult_x_1_n650, mult_x_1_n649,
         mult_x_1_n634, mult_x_1_n633, mult_x_1_n618, mult_x_1_n617,
         mult_x_1_n602, mult_x_1_n601, mult_x_1_n586, mult_x_1_n585,
         mult_x_1_n570, mult_x_1_n569, mult_x_1_n554, mult_x_1_n553,
         mult_x_1_n538, mult_x_1_n537, mult_x_1_n522, mult_x_1_n521,
         mult_x_1_n508, mult_x_1_n507, mult_x_1_n494, mult_x_1_n493,
         mult_x_1_n482, mult_x_1_n481, mult_x_1_n470, mult_x_1_n321,
         mult_x_1_n318, mult_x_1_n317, mult_x_1_n309, mult_x_1_n305,
         mult_x_1_n304, mult_x_1_n298, mult_x_1_n293, mult_x_1_n292,
         mult_x_1_n287, mult_x_1_n286, mult_x_1_n282, mult_x_1_n281,
         mult_x_1_n177, mult_x_1_n176, mult_x_1_n170, mult_x_1_n169,
         mult_x_1_n161, mult_x_1_n160, mult_x_1_n152, mult_x_1_n151,
         mult_x_1_n137, mult_x_1_n136, mult_x_1_n130, mult_x_1_n129,
         mult_x_1_n121, mult_x_1_n120, mult_x_1_n110, mult_x_1_n109,
         mult_x_1_n86, mult_x_1_n85, mult_x_1_n84, mult_x_1_n83, mult_x_1_n58,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321;

  DFFHQXL mult_x_1_clk_r_REG16_S1 ( .D(mult_x_1_n169), .CK(CLK), .Q(n1280) );
  DFFHQXL mult_x_1_clk_r_REG18_S1 ( .D(mult_x_1_n160), .CK(CLK), .Q(n1278) );
  DFFHQXL mult_x_1_clk_r_REG20_S1 ( .D(mult_x_1_n151), .CK(CLK), .Q(n1276) );
  DFFHQX4 mult_x_1_clk_r_REG42_S1 ( .D(mult_x_1_n665), .CK(CLK), .Q(n1320) );
  DFFHQX4 mult_x_1_clk_r_REG41_S1 ( .D(mult_x_1_n650), .CK(CLK), .Q(n1319) );
  DFFHQX4 mult_x_1_clk_r_REG40_S1 ( .D(mult_x_1_n649), .CK(CLK), .Q(n1318) );
  DFFHQX4 mult_x_1_clk_r_REG39_S1 ( .D(mult_x_1_n634), .CK(CLK), .Q(n1317) );
  DFFHQX4 mult_x_1_clk_r_REG38_S1 ( .D(mult_x_1_n633), .CK(CLK), .Q(n1316) );
  DFFHQX4 mult_x_1_clk_r_REG37_S1 ( .D(mult_x_1_n618), .CK(CLK), .Q(n1315) );
  DFFHQX4 mult_x_1_clk_r_REG36_S1 ( .D(mult_x_1_n617), .CK(CLK), .Q(n1314) );
  DFFHQX4 mult_x_1_clk_r_REG35_S1 ( .D(mult_x_1_n602), .CK(CLK), .Q(n1313) );
  DFFHQX4 mult_x_1_clk_r_REG32_S1 ( .D(mult_x_1_n585), .CK(CLK), .Q(n1310) );
  DFFHQX4 mult_x_1_clk_r_REG31_S1 ( .D(mult_x_1_n570), .CK(CLK), .Q(n1309) );
  DFFHQX4 mult_x_1_clk_r_REG56_S1 ( .D(mult_x_1_n309), .CK(CLK), .Q(n1294) );
  DFFHQX1 mult_x_1_clk_r_REG47_S1 ( .D(mult_x_1_n293), .CK(CLK), .Q(n1289) );
  DFFHQX2 mult_x_1_clk_r_REG48_S1 ( .D(mult_x_1_n292), .CK(CLK), .Q(n1288) );
  DFFHQX4 mult_x_1_clk_r_REG53_S1 ( .D(mult_x_1_n305), .CK(CLK), .Q(n1263) );
  DFFHQX4 mult_x_1_clk_r_REG54_S1 ( .D(mult_x_1_n304), .CK(CLK), .Q(n1262) );
  DFFHQX4 mult_x_1_clk_r_REG51_S1 ( .D(n1321), .CK(CLK), .Q(n1260) );
  DFFHQXL mult_x_1_clk_r_REG15_S1 ( .D(mult_x_1_n170), .CK(CLK), .Q(n1281) );
  DFFHQXL mult_x_1_clk_r_REG19_S1 ( .D(mult_x_1_n152), .CK(CLK), .Q(n1277) );
  DFFHQXL mult_x_1_clk_r_REG14_S1 ( .D(mult_x_1_n176), .CK(CLK), .Q(n1282) );
  DFFHQXL mult_x_1_clk_r_REG13_S1 ( .D(mult_x_1_n177), .CK(CLK), .Q(n1283) );
  DFFHQXL clk_r_REG63_S1 ( .D(n1336), .CK(CLK), .Q(PRODUCT[9]) );
  DFFHQXL mult_x_1_clk_r_REG17_S1 ( .D(mult_x_1_n161), .CK(CLK), .Q(n1279) );
  DFFHQXL mult_x_1_clk_r_REG10_S1 ( .D(mult_x_1_n481), .CK(CLK), .Q(n1296) );
  DFFHQXL mult_x_1_clk_r_REG49_S1 ( .D(mult_x_1_n83), .CK(CLK), .Q(n1290) );
  DFFHQXL clk_r_REG71_S1 ( .D(n1344), .CK(CLK), .Q(PRODUCT[1]) );
  DFFHQXL mult_x_1_clk_r_REG22_S1 ( .D(mult_x_1_n136), .CK(CLK), .Q(n1274) );
  DFFHQXL clk_r_REG60_S1 ( .D(n1334), .CK(CLK), .Q(PRODUCT[11]) );
  DFFHQXL mult_x_1_clk_r_REG9_S1 ( .D(mult_x_1_n494), .CK(CLK), .Q(n1299) );
  DFFHQXL clk_r_REG62_S1 ( .D(n1335), .CK(CLK), .Q(PRODUCT[10]) );
  DFFHQXL clk_r_REG64_S1 ( .D(n1337), .CK(CLK), .Q(PRODUCT[8]) );
  DFFHQXL clk_r_REG65_S1 ( .D(n1338), .CK(CLK), .Q(PRODUCT[7]) );
  DFFHQXL clk_r_REG66_S1 ( .D(n1339), .CK(CLK), .Q(PRODUCT[6]) );
  DFFHQXL clk_r_REG67_S1 ( .D(n1340), .CK(CLK), .Q(PRODUCT[5]) );
  DFFHQXL clk_r_REG68_S1 ( .D(n1341), .CK(CLK), .Q(PRODUCT[4]) );
  DFFHQXL clk_r_REG69_S1 ( .D(n1342), .CK(CLK), .Q(PRODUCT[3]) );
  DFFHQXL clk_r_REG70_S1 ( .D(n1343), .CK(CLK), .Q(PRODUCT[2]) );
  DFFHQXL clk_r_REG72_S1 ( .D(n1345), .CK(CLK), .Q(PRODUCT[0]) );
  DFFHQXL mult_x_1_clk_r_REG8_S1 ( .D(mult_x_1_n493), .CK(CLK), .Q(n1298) );
  DFFHQXL mult_x_1_clk_r_REG11_S1 ( .D(mult_x_1_n482), .CK(CLK), .Q(n1297) );
  DFFHQXL mult_x_1_clk_r_REG12_S1 ( .D(mult_x_1_n470), .CK(CLK), .Q(n1295) );
  DFFHQXL mult_x_1_clk_r_REG57_S1 ( .D(mult_x_1_n86), .CK(CLK), .Q(n1293) );
  DFFHQX1 mult_x_1_clk_r_REG55_S1 ( .D(mult_x_1_n85), .CK(CLK), .Q(n1292) );
  DFFHQX2 mult_x_1_clk_r_REG44_S1 ( .D(mult_x_1_n281), .CK(CLK), .Q(n1284) );
  DFFHQXL mult_x_1_clk_r_REG21_S1 ( .D(mult_x_1_n137), .CK(CLK), .Q(n1275) );
  DFFHQXL mult_x_1_clk_r_REG23_S1 ( .D(mult_x_1_n130), .CK(CLK), .Q(n1273) );
  DFFHQXL mult_x_1_clk_r_REG24_S1 ( .D(mult_x_1_n129), .CK(CLK), .Q(n1272) );
  DFFHQXL mult_x_1_clk_r_REG25_S1 ( .D(mult_x_1_n121), .CK(CLK), .Q(n1271) );
  DFFHQXL mult_x_1_clk_r_REG26_S1 ( .D(mult_x_1_n120), .CK(CLK), .Q(n1270) );
  DFFHQXL mult_x_1_clk_r_REG27_S1 ( .D(mult_x_1_n110), .CK(CLK), .Q(n1269) );
  DFFHQXL mult_x_1_clk_r_REG28_S1 ( .D(mult_x_1_n109), .CK(CLK), .Q(n1268) );
  DFFHQXL mult_x_1_clk_r_REG29_S1 ( .D(mult_x_1_n58), .CK(CLK), .Q(n1267) );
  DFFHQX1 mult_x_1_clk_r_REG61_S1 ( .D(mult_x_1_n321), .CK(CLK), .Q(n1266) );
  DFFHQX1 mult_x_1_clk_r_REG58_S1 ( .D(mult_x_1_n318), .CK(CLK), .Q(n1265) );
  DFFHQX1 mult_x_1_clk_r_REG43_S1 ( .D(mult_x_1_n282), .CK(CLK), .Q(n1285) );
  DFFHQX1 mult_x_1_clk_r_REG52_S1 ( .D(mult_x_1_n84), .CK(CLK), .Q(n1291) );
  DFFHQX2 mult_x_1_clk_r_REG46_S1 ( .D(mult_x_1_n286), .CK(CLK), .Q(n1286) );
  DFFHQXL mult_x_1_clk_r_REG7_S1 ( .D(mult_x_1_n508), .CK(CLK), .Q(n1301) );
  DFFHQXL mult_x_1_clk_r_REG4_S1 ( .D(mult_x_1_n521), .CK(CLK), .Q(n1302) );
  DFFHQXL mult_x_1_clk_r_REG59_S1 ( .D(mult_x_1_n317), .CK(CLK), .Q(n1264) );
  DFFHQX2 mult_x_1_clk_r_REG50_S1 ( .D(mult_x_1_n298), .CK(CLK), .Q(n1261) );
  DFFHQX2 mult_x_1_clk_r_REG45_S1 ( .D(mult_x_1_n287), .CK(CLK), .Q(n1287) );
  DFFHQX2 mult_x_1_clk_r_REG34_S1 ( .D(mult_x_1_n601), .CK(CLK), .Q(n1312) );
  DFFHQX2 mult_x_1_clk_r_REG33_S1 ( .D(mult_x_1_n586), .CK(CLK), .Q(n1311) );
  DFFHQX1 mult_x_1_clk_r_REG2_S1 ( .D(mult_x_1_n537), .CK(CLK), .Q(n1304) );
  DFFHQX1 mult_x_1_clk_r_REG5_S1 ( .D(mult_x_1_n522), .CK(CLK), .Q(n1303) );
  DFFHQX2 mult_x_1_clk_r_REG0_S1 ( .D(mult_x_1_n553), .CK(CLK), .Q(n1306) );
  DFFHQX2 mult_x_1_clk_r_REG30_S1 ( .D(mult_x_1_n569), .CK(CLK), .Q(n1308) );
  DFFHQX2 mult_x_1_clk_r_REG1_S1 ( .D(mult_x_1_n554), .CK(CLK), .Q(n1307) );
  DFFHQX2 mult_x_1_clk_r_REG3_S1 ( .D(mult_x_1_n538), .CK(CLK), .Q(n1305) );
  DFFHQX1 mult_x_1_clk_r_REG6_S1 ( .D(mult_x_1_n507), .CK(CLK), .Q(n1300) );
  ADDFHX1 U1 ( .A(n1050), .B(n1049), .CI(n1048), .CO(mult_x_1_n633), .S(
        mult_x_1_n634) );
  ADDFHX2 U2 ( .A(n987), .B(n986), .CI(n985), .CO(n944), .S(n988) );
  ADDFHX2 U3 ( .A(n901), .B(n900), .CI(n899), .CO(n868), .S(n902) );
  XOR2X1 U4 ( .A(n13), .B(n1058), .Y(n1060) );
  ADDFHX1 U5 ( .A(n866), .B(n865), .CI(n864), .CO(n836), .S(n867) );
  ADDFHX2 U6 ( .A(n834), .B(n833), .CI(n832), .CO(n803), .S(n835) );
  ADDFHX2 U7 ( .A(n272), .B(n271), .CI(n270), .CO(n274), .S(n683) );
  ADDFX2 U8 ( .A(n898), .B(n897), .CI(n896), .CO(n901), .S(n940) );
  ADDFX2 U9 ( .A(n863), .B(n862), .CI(n861), .CO(n866), .S(n899) );
  XOR2X1 U10 ( .A(n1057), .B(n1059), .Y(n13) );
  ADDFHX1 U11 ( .A(n1056), .B(n1055), .CI(n1054), .CO(n1061), .S(n1063) );
  ADDFHX1 U12 ( .A(n1047), .B(n1046), .CI(n1045), .CO(n1026), .S(n1048) );
  ADDFX2 U13 ( .A(n984), .B(n983), .CI(n982), .CO(n987), .S(n1022) );
  ADDFHX1 U14 ( .A(n911), .B(n910), .CI(n909), .CO(n895), .S(n935) );
  ADDFHX1 U15 ( .A(n876), .B(n875), .CI(n874), .CO(n860), .S(n894) );
  ADDFHX1 U16 ( .A(n688), .B(n687), .CI(n686), .CO(n270), .S(n709) );
  ADDFHX1 U17 ( .A(n1082), .B(n1081), .CI(n1080), .CO(n555), .S(n1087) );
  ADDFHX2 U18 ( .A(n445), .B(n444), .CI(n443), .CO(n423), .S(n452) );
  ADDFHX2 U19 ( .A(n395), .B(n394), .CI(n393), .CO(n1055), .S(n424) );
  CMPR32X1 U20 ( .A(n364), .B(n363), .C(n362), .CO(n371), .S(n426) );
  XOR2X1 U21 ( .A(n1031), .B(n17), .Y(n16) );
  CMPR32X1 U22 ( .A(n669), .B(n668), .C(n667), .CO(n1081), .S(n1083) );
  CMPR32X1 U23 ( .A(n457), .B(n456), .C(n455), .CO(n443), .S(n479) );
  CMPR32X1 U24 ( .A(n623), .B(n622), .C(n621), .CO(n667), .S(n672) );
  ADDFX2 U25 ( .A(n576), .B(n575), .CI(n574), .CO(n652), .S(n577) );
  INVX1 U26 ( .A(n994), .Y(n6) );
  BUFX4 U27 ( .A(n335), .Y(n994) );
  BUFX3 U28 ( .A(n335), .Y(n1180) );
  CLKBUFX8 U29 ( .A(B[11]), .Y(n920) );
  NAND2X2 U30 ( .A(n335), .B(n57), .Y(n719) );
  XOR2X1 U31 ( .A(B[10]), .B(B[11]), .Y(n27) );
  BUFX3 U32 ( .A(n337), .Y(n9) );
  XNOR2X1 U33 ( .A(B[10]), .B(B[9]), .Y(n341) );
  BUFX3 U34 ( .A(n968), .Y(n41) );
  BUFX3 U35 ( .A(n255), .Y(n966) );
  CLKINVX3 U36 ( .A(n594), .Y(n624) );
  BUFX4 U37 ( .A(n338), .Y(n7) );
  NAND2X1 U38 ( .A(n254), .B(n255), .Y(n968) );
  XNOR2X1 U39 ( .A(n283), .B(n282), .Y(PRODUCT[31]) );
  OAI21XL U40 ( .A0(n5), .A1(n279), .B0(n241), .Y(n283) );
  XOR2X1 U41 ( .A(n79), .B(n34), .Y(PRODUCT[23]) );
  XNOR2X1 U42 ( .A(n326), .B(n325), .Y(PRODUCT[20]) );
  OAI21XL U43 ( .A0(n62), .A1(n321), .B0(n327), .Y(n326) );
  OAI21XL U44 ( .A0(n58), .A1(n121), .B0(n120), .Y(n124) );
  INVX2 U45 ( .A(n58), .Y(n68) );
  INVXL U46 ( .A(n421), .Y(n318) );
  AOI21XL U47 ( .A0(n421), .A1(n331), .B0(n330), .Y(n334) );
  NOR2X1 U48 ( .A(n1314), .B(n1313), .Y(n109) );
  NAND2X1 U49 ( .A(n1316), .B(n1315), .Y(n1069) );
  NOR2X2 U50 ( .A(n322), .B(n321), .Y(n96) );
  OAI22X1 U51 ( .A0(n1155), .A1(n997), .B0(n9), .B1(n996), .Y(n1031) );
  NAND2BX1 U52 ( .AN(n84), .B(n83), .Y(n308) );
  XNOR2X1 U53 ( .A(n124), .B(n123), .Y(PRODUCT[27]) );
  XNOR2XL U54 ( .A(B[1]), .B(n919), .Y(n541) );
  XNOR2XL U55 ( .A(n920), .B(n1067), .Y(n508) );
  XOR2XL U56 ( .A(B[2]), .B(B[3]), .Y(n254) );
  XNOR2XL U57 ( .A(n955), .B(n917), .Y(n489) );
  XNOR2XL U58 ( .A(B[1]), .B(A[25]), .Y(n748) );
  XNOR2XL U59 ( .A(B[1]), .B(n1138), .Y(n880) );
  BUFX1 U60 ( .A(A[23]), .Y(n1156) );
  INVX1 U61 ( .A(B[3]), .Y(n594) );
  XNOR2XL U62 ( .A(n955), .B(n1115), .Y(n261) );
  XNOR2XL U63 ( .A(n920), .B(A[19]), .Y(n224) );
  XNOR2XL U64 ( .A(n955), .B(n925), .Y(n844) );
  XNOR2XL U65 ( .A(n955), .B(n946), .Y(n913) );
  XNOR2XL U66 ( .A(n955), .B(n919), .Y(n385) );
  XNOR2XL U67 ( .A(n1140), .B(n1151), .Y(n171) );
  XNOR2XL U68 ( .A(n920), .B(n1151), .Y(n181) );
  ADDFX2 U69 ( .A(n1085), .B(n1084), .CI(n1083), .CO(n1086), .S(n674) );
  ADDFX2 U70 ( .A(n537), .B(n536), .CI(n535), .CO(n558), .S(n560) );
  ADDFX2 U71 ( .A(n939), .B(n938), .CI(n937), .CO(n942), .S(n985) );
  ADDFX2 U72 ( .A(n801), .B(n800), .CI(n799), .CO(n779), .S(n802) );
  XOR2XL U73 ( .A(n682), .B(n681), .Y(n1336) );
  AND3X4 U74 ( .A(n90), .B(n101), .C(n89), .Y(n5) );
  XNOR2X1 U75 ( .A(n1196), .B(n1195), .Y(n1337) );
  NOR2XL U76 ( .A(n419), .B(n418), .Y(mult_x_1_n281) );
  NAND2XL U77 ( .A(n422), .B(n20), .Y(n19) );
  ADDFHX2 U78 ( .A(n1024), .B(n1023), .CI(n1022), .CO(n989), .S(n1025) );
  ADDFHX1 U79 ( .A(n1065), .B(n1064), .CI(n1063), .CO(mult_x_1_n665), .S(n419)
         );
  NAND2X1 U80 ( .A(n21), .B(n22), .Y(n20) );
  ADDFHX1 U81 ( .A(n945), .B(n944), .CI(n943), .CO(mult_x_1_n585), .S(
        mult_x_1_n586) );
  ADDFHX1 U82 ( .A(n869), .B(n868), .CI(n867), .CO(mult_x_1_n553), .S(
        mult_x_1_n554) );
  INVX1 U83 ( .A(n803), .Y(n25) );
  ADDFHX2 U84 ( .A(n942), .B(n941), .CI(n940), .CO(n903), .S(n943) );
  INVX1 U85 ( .A(n424), .Y(n22) );
  INVX1 U86 ( .A(n804), .Y(n26) );
  NAND2X1 U87 ( .A(n1087), .B(n1086), .Y(n1104) );
  XNOR2X1 U88 ( .A(n751), .B(n750), .Y(n772) );
  NOR2X1 U89 ( .A(n1176), .B(n848), .Y(n878) );
  OR2XL U90 ( .A(n589), .B(n588), .Y(n1248) );
  OAI2BB1XL U91 ( .A0N(n9), .A1N(n1155), .B0(n1154), .Y(n1159) );
  NOR2X1 U92 ( .A(n1176), .B(n390), .Y(n1005) );
  NOR2X1 U93 ( .A(n1176), .B(n918), .Y(n957) );
  OAI22XL U94 ( .A0(n961), .A1(n467), .B0(n412), .B1(n1066), .Y(n466) );
  XNOR2XL U95 ( .A(B[15]), .B(n1151), .Y(n1137) );
  NOR2X1 U96 ( .A(n1227), .B(n129), .Y(n1213) );
  NAND2X1 U97 ( .A(n278), .B(n104), .Y(n1227) );
  AND2X2 U98 ( .A(n1073), .B(n1071), .Y(n34) );
  AND2XL U99 ( .A(n245), .B(n1283), .Y(n36) );
  INVX1 U100 ( .A(n301), .Y(n311) );
  INVX1 U101 ( .A(n1287), .Y(n330) );
  BUFX2 U102 ( .A(A[21]), .Y(n1138) );
  NAND2X1 U103 ( .A(n1305), .B(n1306), .Y(n306) );
  INVX1 U104 ( .A(n1270), .Y(n1215) );
  INVX1 U105 ( .A(n1090), .Y(n1102) );
  OAI2BB1X1 U106 ( .A0N(n424), .A1N(n423), .B0(n19), .Y(n418) );
  XNOR2X1 U107 ( .A(n1206), .B(n1205), .Y(n1338) );
  ADDFHX1 U108 ( .A(n990), .B(n989), .CI(n988), .CO(mult_x_1_n601), .S(
        mult_x_1_n602) );
  ADDFHX1 U109 ( .A(n904), .B(n903), .CI(n902), .CO(mult_x_1_n569), .S(
        mult_x_1_n570) );
  OAI21XL U110 ( .A0(n26), .A1(n25), .B0(n24), .Y(mult_x_1_n521) );
  ADDFHX1 U111 ( .A(n837), .B(n836), .CI(n835), .CO(mult_x_1_n537), .S(
        mult_x_1_n538) );
  INVX1 U112 ( .A(n423), .Y(n21) );
  XNOR3X2 U113 ( .A(n22), .B(n423), .C(n422), .Y(n447) );
  OAI21XL U114 ( .A0(n803), .A1(n804), .B0(n802), .Y(n24) );
  NAND2BXL U115 ( .AN(n416), .B(n30), .Y(n29) );
  INVX1 U116 ( .A(n563), .Y(n46) );
  NAND2X1 U117 ( .A(n674), .B(n673), .Y(n1100) );
  INVXL U118 ( .A(n417), .Y(n30) );
  NAND2X1 U119 ( .A(n616), .B(n615), .Y(n1208) );
  NOR2X1 U120 ( .A(n616), .B(n615), .Y(n1207) );
  ADDFHX1 U121 ( .A(n953), .B(n952), .CI(n951), .CO(n936), .S(n980) );
  NAND2BXL U122 ( .AN(n873), .B(n45), .Y(n43) );
  NAND2BXL U123 ( .AN(n908), .B(n45), .Y(n44) );
  ADDHXL U124 ( .A(n466), .B(n465), .CO(n462), .S(n505) );
  ADDFHX1 U125 ( .A(n700), .B(n699), .CI(n698), .CO(n692), .S(n733) );
  NAND2BX1 U126 ( .AN(n993), .B(n6), .Y(n18) );
  XNOR2XL U127 ( .A(B[16]), .B(A[19]), .Y(n169) );
  OAI22XL U128 ( .A0(n41), .A1(n358), .B0(n966), .B1(n967), .Y(n1007) );
  XNOR2X1 U129 ( .A(n1224), .B(n1223), .Y(PRODUCT[39]) );
  XOR2X1 U130 ( .A(n246), .B(n36), .Y(PRODUCT[32]) );
  XNOR2X1 U131 ( .A(n135), .B(n134), .Y(PRODUCT[37]) );
  XNOR2X1 U132 ( .A(n1200), .B(n1199), .Y(PRODUCT[38]) );
  XNOR2XL U133 ( .A(n920), .B(A[24]), .Y(n170) );
  BUFX8 U134 ( .A(n339), .Y(n8) );
  NOR2BX1 U135 ( .AN(n1067), .B(n10), .Y(n545) );
  NAND2BXL U136 ( .AN(n1067), .B(n955), .Y(n542) );
  NAND2XL U137 ( .A(n73), .B(n1074), .Y(n72) );
  NAND2X1 U138 ( .A(n298), .B(n297), .Y(n299) );
  AND2X2 U139 ( .A(n115), .B(n114), .Y(n35) );
  NAND2X1 U140 ( .A(n111), .B(n110), .Y(n112) );
  NAND2X1 U141 ( .A(n122), .B(n289), .Y(n123) );
  AND2X2 U142 ( .A(n307), .B(n306), .Y(n38) );
  NOR2X1 U143 ( .A(n301), .B(n305), .Y(n118) );
  XOR2X1 U144 ( .A(n1290), .B(n69), .Y(PRODUCT[15]) );
  XOR2X1 U145 ( .A(n499), .B(n1291), .Y(PRODUCT[14]) );
  XOR2X1 U146 ( .A(n523), .B(n1292), .Y(PRODUCT[13]) );
  BUFX2 U147 ( .A(A[9]), .Y(n919) );
  BUFX2 U148 ( .A(A[2]), .Y(n585) );
  NAND2X1 U149 ( .A(n1300), .B(n1299), .Y(n285) );
  INVX1 U150 ( .A(n1276), .Y(n142) );
  INVX1 U151 ( .A(n1278), .Y(n138) );
  NAND2X1 U152 ( .A(n1317), .B(n1318), .Y(n323) );
  BUFX2 U153 ( .A(A[18]), .Y(n883) );
  BUFX2 U154 ( .A(A[20]), .Y(n1115) );
  OAI21XL U155 ( .A0(n1026), .A1(n1027), .B0(n1025), .Y(n49) );
  XNOR3X2 U156 ( .A(n26), .B(n803), .C(n802), .Y(mult_x_1_n522) );
  NAND2X1 U157 ( .A(n556), .B(n555), .Y(n1128) );
  ADDFHX1 U158 ( .A(n479), .B(n478), .CI(n477), .CO(n475), .S(n1098) );
  OR2XL U159 ( .A(n1185), .B(n1184), .Y(n1187) );
  ADDFHX1 U160 ( .A(n474), .B(n473), .CI(n472), .CO(n453), .S(n477) );
  ADDFHX2 U161 ( .A(n672), .B(n671), .CI(n670), .CO(n673), .S(n657) );
  ADDFHX1 U162 ( .A(n562), .B(n561), .CI(n560), .CO(n563), .S(n556) );
  ADDFHX1 U163 ( .A(n505), .B(n504), .CI(n503), .CO(n496), .S(n559) );
  INVXL U164 ( .A(n693), .Y(n94) );
  ADDFHX1 U165 ( .A(n810), .B(n809), .CI(n808), .CO(n798), .S(n827) );
  NAND2XL U166 ( .A(n67), .B(n66), .Y(n65) );
  ADDFHX1 U167 ( .A(n843), .B(n842), .CI(n841), .CO(n828), .S(n859) );
  AND2XL U168 ( .A(n1254), .B(n1253), .Y(n1344) );
  OR2X2 U169 ( .A(n605), .B(n604), .Y(n603) );
  ADDFHX1 U170 ( .A(n644), .B(n643), .CI(n642), .CO(n649), .S(n651) );
  NAND2XL U171 ( .A(n66), .B(n64), .Y(n63) );
  OAI2BB1XL U172 ( .A0N(n1001), .A1N(n8), .B0(n155), .Y(n172) );
  INVXL U173 ( .A(n8), .Y(n67) );
  NOR2X1 U174 ( .A(n749), .B(n1176), .Y(n759) );
  OR2XL U175 ( .A(n1252), .B(n1251), .Y(n1254) );
  NOR2XL U176 ( .A(n1176), .B(n1175), .Y(n1182) );
  XNOR2X1 U177 ( .A(n144), .B(n143), .Y(PRODUCT[35]) );
  OAI2BB1XL U178 ( .A0N(n966), .A1N(n968), .B0(n257), .Y(n712) );
  OAI22X1 U179 ( .A0(n636), .A1(n634), .B0(n541), .B1(n1066), .Y(n633) );
  INVXL U180 ( .A(n1001), .Y(n64) );
  XNOR2XL U181 ( .A(B[16]), .B(A[24]), .Y(n1175) );
  XNOR2XL U182 ( .A(B[16]), .B(n1156), .Y(n1157) );
  OAI2BB1XL U183 ( .A0N(n7), .A1N(n948), .B0(n149), .Y(n190) );
  XNOR2XL U184 ( .A(B[15]), .B(A[25]), .Y(n1177) );
  XNOR2XL U185 ( .A(B[15]), .B(A[24]), .Y(n1158) );
  NAND2X1 U186 ( .A(B[1]), .B(n814), .Y(n636) );
  BUFX8 U187 ( .A(n341), .Y(n10) );
  INVXL U188 ( .A(n139), .Y(n105) );
  INVXL U189 ( .A(n1079), .Y(n76) );
  INVX1 U190 ( .A(B[0]), .Y(n814) );
  BUFX2 U191 ( .A(A[22]), .Y(n1151) );
  BUFX2 U192 ( .A(A[13]), .Y(n946) );
  BUFX2 U193 ( .A(A[16]), .Y(n885) );
  BUFX2 U194 ( .A(A[17]), .Y(n922) );
  NOR2X1 U195 ( .A(n1303), .B(n1304), .Y(n290) );
  NOR2X1 U196 ( .A(n1301), .B(n1302), .Y(n296) );
  BUFX2 U197 ( .A(A[4]), .Y(n917) );
  BUFX2 U198 ( .A(A[8]), .Y(n907) );
  BUFX2 U199 ( .A(A[11]), .Y(n954) );
  BUFX2 U200 ( .A(A[12]), .Y(n912) );
  INVXL U201 ( .A(A[6]), .Y(n33) );
  OAI22X1 U202 ( .A0(n1179), .A1(n342), .B0(n994), .B1(n995), .Y(n1008) );
  NOR2BX1 U203 ( .AN(n1067), .B(n994), .Y(n436) );
  NAND2X4 U204 ( .A(n341), .B(n27), .Y(n1119) );
  OAI22X1 U205 ( .A0(n1119), .A1(n367), .B0(n10), .B1(n366), .Y(n374) );
  NAND2BX1 U206 ( .AN(n102), .B(n308), .Y(n89) );
  NOR2X1 U207 ( .A(n296), .B(n290), .Y(n100) );
  NOR2X4 U208 ( .A(n1319), .B(n1320), .Y(n321) );
  NOR2X4 U209 ( .A(n1318), .B(n1317), .Y(n322) );
  NAND2X2 U210 ( .A(n12), .B(n11), .Y(n1049) );
  NAND2X1 U211 ( .A(n1058), .B(n1059), .Y(n11) );
  OAI21X1 U212 ( .A0(n1058), .A1(n1059), .B0(n1057), .Y(n12) );
  NAND2X1 U213 ( .A(n15), .B(n14), .Y(n1018) );
  NAND2X1 U214 ( .A(n1032), .B(n17), .Y(n14) );
  OAI21XL U215 ( .A0(n1032), .A1(n17), .B0(n1031), .Y(n15) );
  XOR2X1 U216 ( .A(n16), .B(n1032), .Y(n1040) );
  OAI21X2 U217 ( .A0(n1179), .A1(n995), .B0(n18), .Y(n17) );
  INVX1 U218 ( .A(n564), .Y(n47) );
  NAND2X4 U219 ( .A(n23), .B(n338), .Y(n948) );
  XNOR2X1 U220 ( .A(B[6]), .B(B[5]), .Y(n338) );
  XOR2X1 U221 ( .A(B[6]), .B(B[7]), .Y(n23) );
  XNOR2X4 U222 ( .A(B[15]), .B(B[16]), .Y(n1176) );
  OAI2BB1X1 U223 ( .A0N(n29), .A1N(n415), .B0(n28), .Y(n1064) );
  NAND2X1 U224 ( .A(n416), .B(n417), .Y(n28) );
  XOR3X2 U225 ( .A(n417), .B(n416), .C(n415), .Y(n422) );
  AOI21X1 U226 ( .A0(n1264), .A1(n1266), .B0(n1265), .Y(n523) );
  INVX8 U227 ( .A(B[15]), .Y(n344) );
  OAI22X2 U228 ( .A0(n993), .A1(n1179), .B0(n994), .B1(n32), .Y(n56) );
  OAI21X1 U229 ( .A0(n1179), .A1(n32), .B0(n31), .Y(n952) );
  NAND2BX1 U230 ( .AN(n906), .B(n6), .Y(n31) );
  XOR2X1 U231 ( .A(n949), .B(n33), .Y(n32) );
  ADDFX2 U232 ( .A(n442), .B(n441), .CI(n440), .CO(n457), .S(n480) );
  OAI22X1 U233 ( .A0(n8), .A1(n437), .B0(n1001), .B1(n404), .Y(n442) );
  OAI22X1 U234 ( .A0(n1179), .A1(n349), .B0(n994), .B1(n348), .Y(n408) );
  OAI22X1 U235 ( .A0(n8), .A1(n354), .B0(n1001), .B1(n353), .Y(n364) );
  CLKINVX3 U236 ( .A(n594), .Y(n923) );
  XOR2X1 U237 ( .A(n5), .B(n287), .Y(PRODUCT[29]) );
  XNOR2X1 U238 ( .A(n923), .B(A[24]), .Y(n724) );
  XNOR2X1 U239 ( .A(B[11]), .B(B[12]), .Y(n337) );
  OAI22X1 U240 ( .A0(n1179), .A1(n348), .B0(n994), .B1(n347), .Y(n350) );
  XNOR2X1 U241 ( .A(n920), .B(A[14]), .Y(n784) );
  XNOR2X1 U242 ( .A(n920), .B(n925), .Y(n752) );
  OAI22X1 U243 ( .A0(n41), .A1(n753), .B0(n966), .B1(n724), .Y(n756) );
  OAI22X1 U244 ( .A0(n1119), .A1(n752), .B0(n10), .B1(n723), .Y(n757) );
  AOI21X1 U245 ( .A0(n421), .A1(n320), .B0(n319), .Y(n62) );
  OAI21X1 U246 ( .A0(n1284), .A1(n1287), .B0(n1285), .Y(n319) );
  XOR2X2 U247 ( .A(B[15]), .B(B[14]), .Y(n57) );
  OAI22XL U248 ( .A0(n961), .A1(n960), .B0(n959), .B1(n1066), .Y(n1004) );
  XNOR2XL U249 ( .A(n949), .B(A[5]), .Y(n993) );
  NOR2X1 U250 ( .A(n1315), .B(n1316), .Y(n1068) );
  INVXL U251 ( .A(n1274), .Y(n1190) );
  XNOR2XL U252 ( .A(n926), .B(n954), .Y(n396) );
  BUFX3 U253 ( .A(A[15]), .Y(n925) );
  OAI21XL U254 ( .A0(n1234), .A1(n129), .B0(n128), .Y(n1219) );
  INVXL U255 ( .A(n1231), .Y(n128) );
  INVXL U256 ( .A(n1225), .Y(n1218) );
  NAND2X1 U257 ( .A(n206), .B(n360), .Y(n550) );
  XNOR2XL U258 ( .A(n1140), .B(A[19]), .Y(n182) );
  XNOR2XL U259 ( .A(n624), .B(A[25]), .Y(n256) );
  CMPR32X1 U260 ( .A(n266), .B(n265), .C(n264), .CO(n250), .S(n705) );
  OAI22X1 U261 ( .A0(n1155), .A1(n262), .B0(n9), .B1(n220), .Y(n266) );
  NOR2XL U262 ( .A(n1176), .B(n221), .Y(n265) );
  XNOR2XL U263 ( .A(n926), .B(n1156), .Y(n711) );
  XNOR2XL U264 ( .A(n870), .B(A[14]), .Y(n947) );
  XNOR2XL U265 ( .A(n624), .B(A[1]), .Y(n600) );
  BUFX3 U266 ( .A(n550), .Y(n972) );
  XNOR2XL U267 ( .A(n926), .B(A[1]), .Y(n581) );
  XNOR2XL U268 ( .A(n624), .B(n917), .Y(n570) );
  NOR2XL U269 ( .A(n1176), .B(n1152), .Y(n1160) );
  INVXL U270 ( .A(n1153), .Y(n1154) );
  OAI22XL U271 ( .A0(n948), .A1(n991), .B0(n7), .B1(n947), .Y(n999) );
  OAI22XL U272 ( .A0(n8), .A1(n1002), .B0(n1001), .B1(n1000), .Y(n1015) );
  OAI22XL U273 ( .A0(n1179), .A1(n1158), .B0(n1180), .B1(n1177), .Y(n1183) );
  AOI21XL U274 ( .A0(n118), .A1(n308), .B0(n119), .Y(n120) );
  OAI21XL U275 ( .A0(n1234), .A1(n1280), .B0(n1281), .Y(n139) );
  INVXL U276 ( .A(n1219), .Y(n1188) );
  INVXL U277 ( .A(n1213), .Y(n1189) );
  INVXL U278 ( .A(n1279), .Y(n137) );
  NOR2XL U279 ( .A(n1274), .B(n1272), .Y(n1212) );
  NOR2X1 U280 ( .A(n317), .B(n1076), .Y(n98) );
  NAND2BX1 U281 ( .AN(n304), .B(n68), .Y(n82) );
  INVXL U282 ( .A(n305), .Y(n307) );
  INVX1 U283 ( .A(n1069), .Y(n78) );
  NAND2X1 U284 ( .A(n1314), .B(n1313), .Y(n110) );
  NAND2XL U285 ( .A(n59), .B(n314), .Y(n80) );
  XOR2X1 U286 ( .A(n58), .B(n1070), .Y(PRODUCT[21]) );
  INVXL U287 ( .A(n1280), .Y(n202) );
  INVX1 U288 ( .A(n1294), .Y(n499) );
  NAND2BXL U289 ( .AN(n1067), .B(n1140), .Y(n413) );
  XNOR2XL U290 ( .A(n624), .B(A[10]), .Y(n470) );
  XNOR2XL U291 ( .A(n926), .B(n907), .Y(n471) );
  XNOR2XL U292 ( .A(n624), .B(n919), .Y(n509) );
  XNOR2XL U293 ( .A(n870), .B(A[6]), .Y(n469) );
  XNOR2XL U294 ( .A(n1140), .B(n1067), .Y(n460) );
  XNOR2XL U295 ( .A(n1140), .B(A[1]), .Y(n459) );
  XNOR2XL U296 ( .A(n624), .B(n954), .Y(n438) );
  INVX1 U297 ( .A(n1155), .Y(n45) );
  XNOR2XL U298 ( .A(n624), .B(n912), .Y(n406) );
  XNOR2XL U299 ( .A(n1140), .B(n585), .Y(n400) );
  XNOR2XL U300 ( .A(n624), .B(n946), .Y(n361) );
  XNOR2XL U301 ( .A(n1140), .B(A[3]), .Y(n356) );
  XNOR2XL U302 ( .A(n624), .B(A[14]), .Y(n359) );
  XNOR2XL U303 ( .A(n926), .B(n912), .Y(n365) );
  NAND2BXL U304 ( .AN(n1067), .B(n926), .Y(n572) );
  INVX2 U305 ( .A(B[7]), .Y(n566) );
  XNOR2XL U306 ( .A(n926), .B(n585), .Y(n569) );
  XNOR2XL U307 ( .A(n624), .B(n907), .Y(n531) );
  XNOR2XL U308 ( .A(n624), .B(A[5]), .Y(n625) );
  XNOR2XL U309 ( .A(n926), .B(A[3]), .Y(n627) );
  XNOR2XL U310 ( .A(n926), .B(A[5]), .Y(n549) );
  XNOR2XL U311 ( .A(n624), .B(A[6]), .Y(n631) );
  XNOR2XL U312 ( .A(n624), .B(A[7]), .Y(n630) );
  NOR2XL U313 ( .A(n1225), .B(n1268), .Y(n1230) );
  NAND2XL U314 ( .A(n133), .B(n1273), .Y(n134) );
  NAND2XL U315 ( .A(n1213), .B(n1212), .Y(n1198) );
  NAND2XL U316 ( .A(n100), .B(n118), .Y(n102) );
  CMPR32X1 U317 ( .A(n495), .B(n494), .C(n493), .CO(n504), .S(n524) );
  OAI22XL U318 ( .A0(n1119), .A1(n507), .B0(n10), .B1(n468), .Y(n493) );
  NOR2BXL U319 ( .AN(n1067), .B(n9), .Y(n495) );
  OAI22XL U320 ( .A0(n636), .A1(n490), .B0(n467), .B1(n1066), .Y(n494) );
  OAI22X1 U321 ( .A0(n1119), .A1(n492), .B0(n10), .B1(n491), .Y(n48) );
  INVXL U322 ( .A(n920), .Y(n492) );
  NAND2BXL U323 ( .AN(n1067), .B(n920), .Y(n491) );
  OAI22XL U324 ( .A0(n961), .A1(n527), .B0(n490), .B1(n1066), .Y(n512) );
  XNOR2XL U325 ( .A(n926), .B(A[6]), .Y(n530) );
  XNOR2XL U326 ( .A(n926), .B(A[7]), .Y(n510) );
  XNOR2XL U327 ( .A(n955), .B(n585), .Y(n528) );
  OAI22X1 U328 ( .A0(n8), .A1(n151), .B0(n1001), .B1(n542), .Y(n632) );
  INVXL U329 ( .A(n1117), .Y(n1118) );
  OAI22XL U330 ( .A0(n972), .A1(n410), .B0(n970), .B1(n396), .Y(n433) );
  XNOR2XL U331 ( .A(n926), .B(n1138), .Y(n754) );
  OAI22X1 U332 ( .A0(n1155), .A1(n710), .B0(n9), .B1(n262), .Y(n702) );
  OAI22XL U333 ( .A0(n8), .A1(n715), .B0(n1001), .B1(n261), .Y(n703) );
  XNOR2X1 U334 ( .A(n1140), .B(n925), .Y(n710) );
  XNOR2XL U335 ( .A(n1140), .B(A[14]), .Y(n743) );
  OAI22XL U336 ( .A0(n948), .A1(n766), .B0(n7), .B1(n717), .Y(n751) );
  XNOR2XL U337 ( .A(n1140), .B(n946), .Y(n768) );
  XNOR2XL U338 ( .A(n1140), .B(n912), .Y(n807) );
  OAI22XL U339 ( .A0(n961), .A1(n847), .B0(n815), .B1(n814), .Y(n846) );
  XNOR2XL U340 ( .A(n1140), .B(n954), .Y(n840) );
  XNOR2XL U341 ( .A(n1140), .B(A[10]), .Y(n873) );
  OAI22XL U342 ( .A0(n961), .A1(n916), .B0(n880), .B1(n1066), .Y(n915) );
  XNOR2XL U343 ( .A(n1140), .B(n919), .Y(n908) );
  XNOR2XL U344 ( .A(n926), .B(A[14]), .Y(n971) );
  XNOR2XL U345 ( .A(n926), .B(n946), .Y(n386) );
  XNOR2XL U346 ( .A(n1140), .B(A[6]), .Y(n997) );
  XNOR2XL U347 ( .A(n1140), .B(n917), .Y(n355) );
  XNOR2XL U348 ( .A(n1140), .B(A[5]), .Y(n387) );
  NOR2XL U349 ( .A(n1176), .B(n340), .Y(n391) );
  OAI22XL U350 ( .A0(n961), .A1(n345), .B0(n389), .B1(n1066), .Y(n392) );
  NAND2BXL U351 ( .AN(n1067), .B(B[16]), .Y(n340) );
  XNOR2XL U352 ( .A(n1140), .B(n1115), .Y(n161) );
  NOR2XL U353 ( .A(n1176), .B(n153), .Y(n174) );
  OAI22XL U354 ( .A0(n1119), .A1(n158), .B0(n10), .B1(n170), .Y(n175) );
  OAI22XL U355 ( .A0(n1179), .A1(n156), .B0(n1180), .B1(n168), .Y(n177) );
  OAI22XL U356 ( .A0(n1155), .A1(n157), .B0(n9), .B1(n171), .Y(n176) );
  NOR2XL U357 ( .A(n1176), .B(n147), .Y(n192) );
  INVXL U358 ( .A(n148), .Y(n149) );
  NOR2BXL U359 ( .AN(n1067), .B(n1001), .Y(n641) );
  NAND2XL U360 ( .A(n1226), .B(n1230), .Y(n1233) );
  INVXL U361 ( .A(n1228), .Y(n1217) );
  NAND2XL U362 ( .A(n1213), .B(n1218), .Y(n1221) );
  INVXL U363 ( .A(n1268), .Y(n1222) );
  ADDFX2 U364 ( .A(n518), .B(n517), .CI(n516), .CO(n501), .S(n557) );
  NOR2XL U365 ( .A(n1176), .B(n1139), .Y(n1149) );
  INVXL U366 ( .A(n1161), .Y(n1148) );
  OAI22XL U367 ( .A0(n1179), .A1(n1137), .B0(n1180), .B1(n1147), .Y(n1150) );
  OAI22XL U368 ( .A0(n1155), .A1(n1120), .B0(n9), .B1(n1141), .Y(n1144) );
  OAI22XL U369 ( .A0(n1179), .A1(n1121), .B0(n1180), .B1(n1137), .Y(n1143) );
  INVXL U370 ( .A(n191), .Y(n212) );
  OAI22XL U371 ( .A0(n1155), .A1(n219), .B0(n9), .B1(n182), .Y(n214) );
  OAI22XL U372 ( .A0(n8), .A1(n217), .B0(n1001), .B1(n183), .Y(n213) );
  ADDFX2 U373 ( .A(n211), .B(n210), .CI(n209), .CO(n193), .S(n248) );
  OAI22XL U374 ( .A0(n1119), .A1(n218), .B0(n10), .B1(n186), .Y(n209) );
  NOR2XL U375 ( .A(n1176), .B(n184), .Y(n211) );
  OAI22XL U376 ( .A0(n1179), .A1(n216), .B0(n1180), .B1(n185), .Y(n210) );
  OAI22XL U377 ( .A0(n1155), .A1(n220), .B0(n9), .B1(n219), .Y(n251) );
  OAI22XL U378 ( .A0(n1119), .A1(n224), .B0(n10), .B1(n218), .Y(n252) );
  OAI22XL U379 ( .A0(n948), .A1(n695), .B0(n7), .B1(n260), .Y(n698) );
  OAI22X2 U380 ( .A0(n1179), .A1(n697), .B0(n1180), .B1(n259), .Y(n699) );
  OAI21XL U381 ( .A0(n261), .A1(n8), .B0(n63), .Y(n694) );
  NOR2XL U382 ( .A(n1176), .B(n253), .Y(n714) );
  CMPR32X1 U383 ( .A(n746), .B(n745), .C(n744), .CO(n734), .S(n764) );
  INVXL U384 ( .A(n56), .Y(n54) );
  OAI22XL U385 ( .A0(n8), .A1(n1000), .B0(n1001), .B1(n956), .Y(n978) );
  ADDFX2 U386 ( .A(n1021), .B(n1020), .CI(n1019), .CO(n1024), .S(n1045) );
  ADDFX2 U387 ( .A(n1044), .B(n1043), .CI(n1042), .CO(n1047), .S(n1057) );
  NOR2BXL U388 ( .AN(n1067), .B(n970), .Y(n612) );
  OAI22XL U389 ( .A0(n961), .A1(n598), .B0(n597), .B1(n1066), .Y(n611) );
  OAI22XL U390 ( .A0(n41), .A1(n600), .B0(n966), .B1(n599), .Y(n610) );
  OAI22XL U391 ( .A0(n972), .A1(n582), .B0(n970), .B1(n581), .Y(n608) );
  OAI22XL U392 ( .A0(n41), .A1(n599), .B0(n966), .B1(n580), .Y(n609) );
  XNOR2XL U393 ( .A(n926), .B(n1067), .Y(n582) );
  OAI22XL U394 ( .A0(n41), .A1(n580), .B0(n966), .B1(n570), .Y(n579) );
  OAI22XL U395 ( .A0(n961), .A1(n1067), .B0(n586), .B1(n1066), .Y(n1252) );
  NAND2XL U396 ( .A(n587), .B(n961), .Y(n1251) );
  NAND2BXL U397 ( .AN(n1067), .B(B[1]), .Y(n587) );
  NAND2XL U398 ( .A(n1252), .B(n1251), .Y(n1253) );
  INVXL U399 ( .A(n1177), .Y(n1178) );
  NOR2XL U400 ( .A(n1176), .B(n1157), .Y(n1174) );
  INVXL U401 ( .A(n1183), .Y(n1173) );
  XOR2X1 U402 ( .A(n998), .B(n56), .Y(n55) );
  AOI21XL U403 ( .A0(n1240), .A1(n603), .B0(n606), .Y(n1258) );
  INVXL U404 ( .A(n1239), .Y(n606) );
  NOR2XL U405 ( .A(n614), .B(n613), .Y(n1255) );
  NAND2XL U406 ( .A(n614), .B(n613), .Y(n1256) );
  NOR2X1 U407 ( .A(n618), .B(n617), .Y(n1202) );
  INVXL U408 ( .A(n1201), .Y(n1210) );
  NOR2X1 U409 ( .A(n1284), .B(n1286), .Y(n320) );
  NAND2XL U410 ( .A(n314), .B(n1073), .Y(n1075) );
  NOR2XL U411 ( .A(n1295), .B(n1296), .Y(n239) );
  INVXL U412 ( .A(n1275), .Y(n130) );
  INVXL U413 ( .A(n1272), .Y(n133) );
  NAND2XL U414 ( .A(n1212), .B(n1215), .Y(n1225) );
  NAND2XL U415 ( .A(n286), .B(n285), .Y(n287) );
  INVXL U416 ( .A(n284), .Y(n286) );
  AOI21XL U417 ( .A0(n1262), .A1(n1294), .B0(n1263), .Y(n69) );
  INVXL U418 ( .A(n239), .Y(n281) );
  INVXL U419 ( .A(n113), .Y(n115) );
  NAND2X1 U420 ( .A(n1320), .B(n1319), .Y(n327) );
  XNOR2X1 U421 ( .A(n313), .B(n312), .Y(PRODUCT[25]) );
  OAI21XL U422 ( .A0(n58), .A1(n117), .B0(n309), .Y(n313) );
  NAND2XL U423 ( .A(n1075), .B(n76), .Y(n73) );
  NOR2XL U424 ( .A(n1075), .B(n76), .Y(n74) );
  INVXL U425 ( .A(n1282), .Y(n245) );
  NAND2X1 U426 ( .A(n1262), .B(n1260), .Y(n449) );
  CLKINVX3 U427 ( .A(B[9]), .Y(n151) );
  XNOR2XL U428 ( .A(n926), .B(n919), .Y(n439) );
  XNOR2XL U429 ( .A(n926), .B(A[10]), .Y(n410) );
  XNOR2XL U430 ( .A(B[16]), .B(n946), .Y(n221) );
  XNOR2X1 U431 ( .A(n1140), .B(n885), .Y(n262) );
  XNOR2XL U432 ( .A(n923), .B(n1151), .Y(n785) );
  XNOR2XL U433 ( .A(n926), .B(n1115), .Y(n786) );
  XNOR2XL U434 ( .A(n923), .B(n1138), .Y(n818) );
  XNOR2XL U435 ( .A(n920), .B(n946), .Y(n817) );
  XNOR2XL U436 ( .A(n926), .B(A[19]), .Y(n819) );
  XNOR2XL U437 ( .A(n923), .B(n1115), .Y(n850) );
  XNOR2XL U438 ( .A(n920), .B(n912), .Y(n849) );
  XNOR2XL U439 ( .A(n926), .B(n883), .Y(n851) );
  XNOR2XL U440 ( .A(n923), .B(A[19]), .Y(n884) );
  XNOR2XL U441 ( .A(n920), .B(n954), .Y(n882) );
  XNOR2XL U442 ( .A(n926), .B(n922), .Y(n886) );
  XNOR2XL U443 ( .A(n923), .B(n883), .Y(n924) );
  XNOR2X1 U444 ( .A(n920), .B(A[10]), .Y(n921) );
  XNOR2XL U445 ( .A(n926), .B(n885), .Y(n927) );
  XNOR2XL U446 ( .A(n923), .B(n922), .Y(n965) );
  XNOR2XL U447 ( .A(n920), .B(n919), .Y(n963) );
  XNOR2XL U448 ( .A(n926), .B(n925), .Y(n969) );
  INVXL U449 ( .A(n154), .Y(n155) );
  XNOR2XL U450 ( .A(B[16]), .B(n885), .Y(n147) );
  XNOR2XL U451 ( .A(B[7]), .B(n585), .Y(n637) );
  XNOR2XL U452 ( .A(n955), .B(n1067), .Y(n548) );
  XNOR2XL U453 ( .A(n926), .B(n917), .Y(n626) );
  NAND2XL U454 ( .A(n1190), .B(n1275), .Y(n1191) );
  AOI21XL U455 ( .A0(n137), .A1(n142), .B0(n125), .Y(n126) );
  INVXL U456 ( .A(n1277), .Y(n125) );
  AOI21XL U457 ( .A0(n1216), .A1(n1215), .B0(n1214), .Y(n1228) );
  INVXL U458 ( .A(n1271), .Y(n1214) );
  INVXL U459 ( .A(n102), .Y(n85) );
  XOR2X2 U460 ( .A(n77), .B(n112), .Y(PRODUCT[22]) );
  NAND2X1 U461 ( .A(n80), .B(n316), .Y(n79) );
  OAI21XL U462 ( .A0(n68), .A1(n75), .B0(n70), .Y(PRODUCT[24]) );
  NAND2XL U463 ( .A(n1074), .B(n76), .Y(n75) );
  AOI22X1 U464 ( .A0(n68), .A1(n74), .B0(n72), .B1(n71), .Y(n70) );
  NAND2XL U465 ( .A(n202), .B(n1281), .Y(n203) );
  NAND2XL U466 ( .A(n142), .B(n1277), .Y(n143) );
  XNOR2X1 U467 ( .A(n108), .B(n107), .Y(PRODUCT[34]) );
  NAND2XL U468 ( .A(n138), .B(n1279), .Y(n107) );
  OAI21XL U469 ( .A0(n5), .A1(n106), .B0(n105), .Y(n108) );
  OAI22XL U470 ( .A0(n1155), .A1(n459), .B0(n9), .B1(n400), .Y(n434) );
  INVXL U471 ( .A(n1140), .Y(n414) );
  CMPR32X1 U472 ( .A(n488), .B(n487), .C(n486), .CO(n481), .S(n517) );
  OAI22XL U473 ( .A0(n972), .A1(n471), .B0(n970), .B1(n439), .Y(n486) );
  OAI22XL U474 ( .A0(n8), .A1(n489), .B0(n1001), .B1(n437), .Y(n488) );
  OAI22XL U475 ( .A0(n41), .A1(n470), .B0(n966), .B1(n438), .Y(n487) );
  OAI22XL U476 ( .A0(n972), .A1(n510), .B0(n970), .B1(n471), .Y(n513) );
  OAI22XL U477 ( .A0(n41), .A1(n509), .B0(n966), .B1(n470), .Y(n514) );
  OAI22XL U478 ( .A0(n41), .A1(n531), .B0(n966), .B1(n509), .Y(n532) );
  OAI22XL U479 ( .A0(n1119), .A1(n508), .B0(n10), .B1(n507), .Y(n533) );
  CMPR32X1 U480 ( .A(n545), .B(n544), .C(n543), .CO(n553), .S(n668) );
  OAI22XL U481 ( .A0(n8), .A1(n547), .B0(n1001), .B1(n528), .Y(n543) );
  XNOR2XL U482 ( .A(B[16]), .B(n1151), .Y(n1152) );
  XNOR2XL U483 ( .A(B[16]), .B(n1138), .Y(n1139) );
  XNOR2XL U484 ( .A(n1140), .B(A[24]), .Y(n1141) );
  OAI22XL U485 ( .A0(n1119), .A1(n468), .B0(n10), .B1(n461), .Y(n483) );
  OAI22XL U486 ( .A0(n1155), .A1(n460), .B0(n9), .B1(n459), .Y(n484) );
  ADDFX2 U487 ( .A(n464), .B(n463), .CI(n462), .CO(n455), .S(n497) );
  OAI22XL U488 ( .A0(n550), .A1(n439), .B0(n970), .B1(n410), .Y(n464) );
  OAI22X1 U489 ( .A0(n948), .A1(n458), .B0(n7), .B1(n411), .Y(n463) );
  OAI22XL U490 ( .A0(n41), .A1(n438), .B0(n966), .B1(n406), .Y(n440) );
  OAI22XL U491 ( .A0(n1119), .A1(n461), .B0(n10), .B1(n405), .Y(n441) );
  XNOR2XL U492 ( .A(B[16]), .B(n925), .Y(n184) );
  XNOR2XL U493 ( .A(n920), .B(n883), .Y(n263) );
  XNOR2XL U494 ( .A(n926), .B(A[25]), .Y(n207) );
  XNOR2XL U495 ( .A(B[16]), .B(A[14]), .Y(n205) );
  XNOR2X1 U496 ( .A(n1140), .B(n922), .Y(n220) );
  XNOR2XL U497 ( .A(n920), .B(n1115), .Y(n218) );
  XNOR2XL U498 ( .A(n1140), .B(n883), .Y(n219) );
  XNOR2X1 U499 ( .A(n949), .B(A[14]), .Y(n259) );
  XNOR2XL U500 ( .A(n926), .B(A[24]), .Y(n258) );
  INVXL U501 ( .A(n748), .Y(n725) );
  XNOR2XL U502 ( .A(n923), .B(n1156), .Y(n753) );
  OAI22XL U503 ( .A0(n8), .A1(n811), .B0(n1001), .B1(n758), .Y(n792) );
  ADDFX2 U504 ( .A(n789), .B(n788), .CI(n787), .CO(n795), .S(n830) );
  OAI22XL U505 ( .A0(n972), .A1(n786), .B0(n970), .B1(n754), .Y(n787) );
  OAI22XL U506 ( .A0(n1119), .A1(n784), .B0(n10), .B1(n752), .Y(n789) );
  OAI22XL U507 ( .A0(n41), .A1(n785), .B0(n966), .B1(n753), .Y(n788) );
  ADDFX2 U508 ( .A(n822), .B(n821), .CI(n820), .CO(n831), .S(n862) );
  OAI22XL U509 ( .A0(n972), .A1(n819), .B0(n970), .B1(n786), .Y(n820) );
  OAI22X1 U510 ( .A0(n41), .A1(n818), .B0(n966), .B1(n785), .Y(n821) );
  OAI22XL U511 ( .A0(n1119), .A1(n817), .B0(n10), .B1(n784), .Y(n822) );
  CMPR32X1 U512 ( .A(n854), .B(n853), .C(n852), .CO(n863), .S(n897) );
  OAI22XL U513 ( .A0(n972), .A1(n851), .B0(n970), .B1(n819), .Y(n852) );
  OAI22XL U514 ( .A0(n1119), .A1(n849), .B0(n10), .B1(n817), .Y(n854) );
  OAI22XL U515 ( .A0(n41), .A1(n850), .B0(n966), .B1(n818), .Y(n853) );
  CMPR32X1 U516 ( .A(n889), .B(n888), .C(n887), .CO(n898), .S(n938) );
  OAI22XL U517 ( .A0(n972), .A1(n886), .B0(n970), .B1(n851), .Y(n887) );
  OAI22XL U518 ( .A0(n1119), .A1(n882), .B0(n10), .B1(n849), .Y(n889) );
  OAI22XL U519 ( .A0(n41), .A1(n884), .B0(n966), .B1(n850), .Y(n888) );
  XNOR2XL U520 ( .A(n955), .B(n954), .Y(n1000) );
  CMPR32X1 U521 ( .A(n930), .B(n929), .C(n928), .CO(n939), .S(n983) );
  OAI22XL U522 ( .A0(n972), .A1(n927), .B0(n970), .B1(n886), .Y(n928) );
  OAI22XL U523 ( .A0(n1119), .A1(n921), .B0(n10), .B1(n882), .Y(n930) );
  OAI22XL U524 ( .A0(n41), .A1(n924), .B0(n966), .B1(n884), .Y(n929) );
  CMPR32X1 U525 ( .A(n975), .B(n974), .C(n973), .CO(n984), .S(n1020) );
  OAI22XL U526 ( .A0(n972), .A1(n969), .B0(n970), .B1(n927), .Y(n973) );
  OAI22XL U527 ( .A0(n1119), .A1(n963), .B0(n10), .B1(n921), .Y(n975) );
  OAI22XL U528 ( .A0(n41), .A1(n965), .B0(n966), .B1(n924), .Y(n974) );
  CMPR32X1 U529 ( .A(n1012), .B(n1011), .C(n1010), .CO(n1021), .S(n1043) );
  OAI22XL U530 ( .A0(n972), .A1(n971), .B0(n970), .B1(n969), .Y(n1010) );
  OAI22XL U531 ( .A0(n1119), .A1(n964), .B0(n10), .B1(n963), .Y(n1012) );
  OAI22XL U532 ( .A0(n41), .A1(n967), .B0(n966), .B1(n965), .Y(n1011) );
  OAI22XL U533 ( .A0(n948), .A1(n411), .B0(n7), .B1(n369), .Y(n428) );
  OAI22XL U534 ( .A0(n1119), .A1(n405), .B0(n10), .B1(n367), .Y(n429) );
  OAI22XL U535 ( .A0(n41), .A1(n406), .B0(n966), .B1(n361), .Y(n430) );
  ADDFX2 U536 ( .A(n409), .B(n408), .CI(n407), .CO(n401), .S(n456) );
  OAI22XL U537 ( .A0(n1155), .A1(n400), .B0(n9), .B1(n356), .Y(n407) );
  OAI22XL U538 ( .A0(n8), .A1(n404), .B0(n1001), .B1(n354), .Y(n409) );
  OAI22X1 U539 ( .A0(n1179), .A1(n344), .B0(n1180), .B1(n343), .Y(n397) );
  NAND2BXL U540 ( .AN(n1067), .B(n949), .Y(n343) );
  NOR2BXL U541 ( .AN(n1067), .B(n1176), .Y(n352) );
  OAI22XL U542 ( .A0(n961), .A1(n346), .B0(n345), .B1(n1066), .Y(n351) );
  OAI22XL U543 ( .A0(n550), .A1(n396), .B0(n970), .B1(n365), .Y(n375) );
  OAI22XL U544 ( .A0(n948), .A1(n369), .B0(n7), .B1(n368), .Y(n373) );
  ADDFX2 U545 ( .A(n384), .B(n383), .CI(n382), .CO(n1038), .S(n370) );
  OAI22XL U546 ( .A0(n972), .A1(n365), .B0(n970), .B1(n386), .Y(n382) );
  OAI22XL U547 ( .A0(n1119), .A1(n366), .B0(n10), .B1(n357), .Y(n384) );
  OAI22X1 U548 ( .A0(n41), .A1(n359), .B0(n966), .B1(n358), .Y(n383) );
  XNOR2XL U549 ( .A(n920), .B(A[7]), .Y(n357) );
  XNOR2XL U550 ( .A(n923), .B(n925), .Y(n358) );
  XNOR2XL U551 ( .A(n923), .B(n885), .Y(n967) );
  XNOR2XL U552 ( .A(n920), .B(n907), .Y(n964) );
  INVXL U553 ( .A(n173), .Y(n162) );
  OAI22XL U554 ( .A0(n1155), .A1(n182), .B0(n9), .B1(n161), .Y(n187) );
  OAI22XL U555 ( .A0(n8), .A1(n183), .B0(n1001), .B1(n159), .Y(n189) );
  XNOR2XL U556 ( .A(n624), .B(n585), .Y(n599) );
  XNOR2XL U557 ( .A(n624), .B(A[3]), .Y(n580) );
  INVXL U558 ( .A(n926), .Y(n573) );
  OAI22XL U559 ( .A0(n961), .A1(n567), .B0(n635), .B1(n1066), .Y(n629) );
  NAND2BXL U560 ( .AN(n1067), .B(n870), .Y(n565) );
  OAI22XL U561 ( .A0(n972), .A1(n581), .B0(n970), .B1(n569), .Y(n574) );
  OAI22XL U562 ( .A0(n972), .A1(n569), .B0(n970), .B1(n627), .Y(n642) );
  OAI22XL U563 ( .A0(n972), .A1(n549), .B0(n970), .B1(n530), .Y(n662) );
  OAI22XL U564 ( .A0(n41), .A1(n630), .B0(n966), .B1(n531), .Y(n661) );
  CMPR32X1 U565 ( .A(n647), .B(n646), .C(n645), .CO(n671), .S(n648) );
  OAI22XL U566 ( .A0(n972), .A1(n627), .B0(n970), .B1(n626), .Y(n646) );
  OAI22XL U567 ( .A0(n41), .A1(n625), .B0(n966), .B1(n631), .Y(n647) );
  OAI22XL U568 ( .A0(n41), .A1(n631), .B0(n966), .B1(n630), .Y(n666) );
  NAND2XL U569 ( .A(n1215), .B(n1271), .Y(n1199) );
  OAI22XL U570 ( .A0(n8), .A1(n511), .B0(n1001), .B1(n489), .Y(n526) );
  AND2X1 U571 ( .A(n48), .B(n512), .Y(n525) );
  OAI22XL U572 ( .A0(n550), .A1(n530), .B0(n970), .B1(n510), .Y(n540) );
  XOR2XL U573 ( .A(n48), .B(n512), .Y(n538) );
  OAI22XL U574 ( .A0(n8), .A1(n528), .B0(n1001), .B1(n511), .Y(n539) );
  NOR2XL U575 ( .A(n1176), .B(n1116), .Y(n1136) );
  OAI2BB1XL U576 ( .A0N(n10), .A1N(n1119), .B0(n1118), .Y(n1134) );
  XNOR2XL U577 ( .A(B[16]), .B(n1115), .Y(n1116) );
  CMPR32X1 U578 ( .A(n269), .B(n268), .C(n267), .CO(n688), .S(n704) );
  OAI22XL U579 ( .A0(n1119), .A1(n263), .B0(n10), .B1(n224), .Y(n267) );
  OAI22XL U580 ( .A0(n948), .A1(n260), .B0(n7), .B1(n222), .Y(n269) );
  OAI22XL U581 ( .A0(n1179), .A1(n259), .B0(n1180), .B1(n223), .Y(n268) );
  OAI21XL U582 ( .A0(n217), .A1(n1001), .B0(n65), .Y(n228) );
  OAI22XL U583 ( .A0(n948), .A1(n222), .B0(n7), .B1(n215), .Y(n230) );
  OAI22XL U584 ( .A0(n1179), .A1(n223), .B0(n1180), .B1(n216), .Y(n229) );
  CMPR32X1 U585 ( .A(n227), .B(n226), .C(n225), .CO(n249), .S(n687) );
  OAI2BB1XL U586 ( .A0N(n970), .A1N(n972), .B0(n208), .Y(n225) );
  NOR2XL U587 ( .A(n1176), .B(n205), .Y(n227) );
  INVXL U588 ( .A(n207), .Y(n208) );
  OAI22XL U589 ( .A0(n8), .A1(n758), .B0(n1001), .B1(n747), .Y(n774) );
  OAI22XL U590 ( .A0(n1155), .A1(n768), .B0(n9), .B1(n743), .Y(n769) );
  OAI22XL U591 ( .A0(n972), .A1(n754), .B0(n970), .B1(n741), .Y(n771) );
  OAI22XL U592 ( .A0(n972), .A1(n741), .B0(n970), .B1(n711), .Y(n727) );
  OAI22XL U593 ( .A0(n8), .A1(n747), .B0(n1001), .B1(n715), .Y(n731) );
  OR2XL U594 ( .A(n751), .B(n750), .Y(n729) );
  ADDFX2 U595 ( .A(n757), .B(n756), .CI(n755), .CO(n783), .S(n794) );
  OAI2BB1XL U596 ( .A0N(n1066), .A1N(n961), .B0(n725), .Y(n755) );
  OAI22XL U597 ( .A0(n1155), .A1(n807), .B0(n9), .B1(n768), .Y(n808) );
  OAI22XL U598 ( .A0(n8), .A1(n844), .B0(n1001), .B1(n811), .Y(n825) );
  ADDFX2 U599 ( .A(n795), .B(n794), .CI(n793), .CO(n801), .S(n833) );
  OAI22XL U600 ( .A0(n8), .A1(n877), .B0(n1001), .B1(n844), .Y(n857) );
  ADDFX2 U601 ( .A(n831), .B(n830), .CI(n829), .CO(n834), .S(n864) );
  OAI21XL U602 ( .A0(n840), .A1(n9), .B0(n43), .Y(n874) );
  OAI22XL U603 ( .A0(n8), .A1(n913), .B0(n1001), .B1(n877), .Y(n892) );
  OAI21XL U604 ( .A0(n873), .A1(n9), .B0(n44), .Y(n909) );
  OAI22XL U605 ( .A0(n8), .A1(n956), .B0(n1001), .B1(n913), .Y(n933) );
  OAI22XL U606 ( .A0(n1155), .A1(n387), .B0(n9), .B1(n997), .Y(n1028) );
  OAI22XL U607 ( .A0(n8), .A1(n385), .B0(n1001), .B1(n1002), .Y(n1030) );
  ADDFX2 U608 ( .A(n427), .B(n426), .CI(n425), .CO(n415), .S(n454) );
  ADDFX2 U609 ( .A(n403), .B(n402), .CI(n401), .CO(n417), .S(n444) );
  ADDFX2 U610 ( .A(n1038), .B(n1037), .CI(n1036), .CO(n1059), .S(n1054) );
  OAI22XL U611 ( .A0(n1155), .A1(n355), .B0(n9), .B1(n387), .Y(n376) );
  CMPR32X1 U612 ( .A(n381), .B(n380), .C(n379), .CO(n1052), .S(n393) );
  OAI22XL U613 ( .A0(n8), .A1(n353), .B0(n1001), .B1(n385), .Y(n380) );
  NOR2XL U614 ( .A(n1176), .B(n169), .Y(n1123) );
  OAI22XL U615 ( .A0(n1179), .A1(n168), .B0(n1180), .B1(n1121), .Y(n1124) );
  INVXL U616 ( .A(n1135), .Y(n1122) );
  OAI22XL U617 ( .A0(n1155), .A1(n171), .B0(n9), .B1(n1120), .Y(n1127) );
  NOR2XL U618 ( .A(n1176), .B(n146), .Y(n166) );
  OAI22XL U619 ( .A0(n1155), .A1(n161), .B0(n9), .B1(n157), .Y(n167) );
  XNOR2XL U620 ( .A(B[16]), .B(n922), .Y(n146) );
  OAI22XL U621 ( .A0(n1119), .A1(n186), .B0(n10), .B1(n181), .Y(n195) );
  OAI22XL U622 ( .A0(n961), .A1(n586), .B0(n591), .B1(n1066), .Y(n589) );
  NOR2BXL U623 ( .AN(n1067), .B(n966), .Y(n588) );
  OAI22XL U624 ( .A0(n41), .A1(n594), .B0(n966), .B1(n593), .Y(n595) );
  NAND2BXL U625 ( .AN(n1067), .B(n624), .Y(n593) );
  XNOR2XL U626 ( .A(n624), .B(n1067), .Y(n592) );
  XNOR2XL U627 ( .A(n1238), .B(n1267), .Y(PRODUCT[40]) );
  INVXL U628 ( .A(n1235), .Y(n1236) );
  NAND2XL U629 ( .A(n1222), .B(n1269), .Y(n1223) );
  OAI22XL U630 ( .A0(n1179), .A1(n1147), .B0(n1180), .B1(n1158), .Y(n1167) );
  NAND2X1 U631 ( .A(n93), .B(n92), .Y(n690) );
  OAI21XL U632 ( .A0(n693), .A1(n694), .B0(n692), .Y(n93) );
  NAND2XL U633 ( .A(n693), .B(n694), .Y(n92) );
  OAI2BB1XL U634 ( .A0N(n999), .A1N(n56), .B0(n52), .Y(n981) );
  NAND2BXL U635 ( .AN(n999), .B(n54), .Y(n53) );
  ADDFX2 U636 ( .A(n1041), .B(n1040), .CI(n1039), .CO(n1050), .S(n1058) );
  ADDFX2 U637 ( .A(n1053), .B(n1052), .CI(n1051), .CO(n1062), .S(n1065) );
  NAND2XL U638 ( .A(n589), .B(n588), .Y(n1247) );
  INVXL U639 ( .A(n1253), .Y(n1249) );
  NOR2XL U640 ( .A(n596), .B(n595), .Y(n1242) );
  NAND2XL U641 ( .A(n596), .B(n595), .Y(n1243) );
  AOI21XL U642 ( .A0(n1248), .A1(n1249), .B0(n590), .Y(n1245) );
  INVXL U643 ( .A(n1247), .Y(n590) );
  NAND2XL U644 ( .A(n605), .B(n604), .Y(n1239) );
  NOR2XL U645 ( .A(n1130), .B(n1129), .Y(mult_x_1_n136) );
  NAND2XL U646 ( .A(n680), .B(n679), .Y(n681) );
  NAND2XL U647 ( .A(n1187), .B(n1186), .Y(mult_x_1_n58) );
  NAND2XL U648 ( .A(n1185), .B(n1184), .Y(n1186) );
  NOR2XL U649 ( .A(n1169), .B(n1168), .Y(mult_x_1_n109) );
  NAND2XL U650 ( .A(n1169), .B(n1168), .Y(mult_x_1_n110) );
  NOR2XL U651 ( .A(n1171), .B(n1170), .Y(mult_x_1_n120) );
  NAND2XL U652 ( .A(n1171), .B(n1170), .Y(mult_x_1_n121) );
  NOR2XL U653 ( .A(n1146), .B(n1145), .Y(mult_x_1_n129) );
  NAND2XL U654 ( .A(n1146), .B(n1145), .Y(mult_x_1_n130) );
  NAND2XL U655 ( .A(n1130), .B(n1129), .Y(mult_x_1_n137) );
  OAI21XL U656 ( .A0(n51), .A1(n50), .B0(n49), .Y(mult_x_1_n617) );
  INVXL U657 ( .A(n1026), .Y(n50) );
  NOR2XL U658 ( .A(n1109), .B(n1108), .Y(mult_x_1_n151) );
  NOR2XL U659 ( .A(n1111), .B(n1110), .Y(mult_x_1_n160) );
  NOR2BXL U660 ( .AN(n1067), .B(n1066), .Y(n1345) );
  XNOR2XL U661 ( .A(n1250), .B(n1249), .Y(n1343) );
  NAND2XL U662 ( .A(n1248), .B(n1247), .Y(n1250) );
  XOR2XL U663 ( .A(n1246), .B(n1245), .Y(n1342) );
  NAND2XL U664 ( .A(n1244), .B(n1243), .Y(n1246) );
  INVXL U665 ( .A(n1242), .Y(n1244) );
  XNOR2XL U666 ( .A(n1241), .B(n1240), .Y(n1341) );
  NAND2XL U667 ( .A(n603), .B(n1239), .Y(n1241) );
  NAND2XL U668 ( .A(n1257), .B(n1256), .Y(n1259) );
  INVXL U669 ( .A(n1255), .Y(n1257) );
  XOR2XL U670 ( .A(n1211), .B(n1210), .Y(n1339) );
  NAND2XL U671 ( .A(n1209), .B(n1208), .Y(n1211) );
  INVXL U672 ( .A(n1207), .Y(n1209) );
  NAND2XL U673 ( .A(n1204), .B(n1203), .Y(n1205) );
  NAND2XL U674 ( .A(n1194), .B(n1193), .Y(n1195) );
  NOR2X1 U675 ( .A(n1068), .B(n109), .Y(n314) );
  INVX1 U676 ( .A(n117), .Y(n91) );
  INVX1 U677 ( .A(n1068), .Y(n86) );
  AND2X1 U678 ( .A(n96), .B(n320), .Y(n37) );
  CMPR22X1 U679 ( .A(n813), .B(n812), .CO(n790), .S(n824) );
  CMPR22X1 U680 ( .A(n879), .B(n878), .CO(n855), .S(n891) );
  CMPR22X1 U681 ( .A(n958), .B(n957), .CO(n931), .S(n977) );
  CMPR22X1 U682 ( .A(n1006), .B(n1005), .CO(n1013), .S(n1034) );
  INVXL U683 ( .A(n653), .Y(n39) );
  INVXL U684 ( .A(n39), .Y(n40) );
  NOR2X1 U685 ( .A(n1300), .B(n1299), .Y(n284) );
  OAI22X1 U686 ( .A0(n8), .A1(n159), .B0(n1001), .B1(n154), .Y(n173) );
  CMPR22X1 U687 ( .A(n760), .B(n759), .CO(n773), .S(n791) );
  CMPR22X1 U688 ( .A(n584), .B(n583), .CO(n578), .S(n607) );
  XOR2X1 U689 ( .A(n999), .B(n55), .Y(n1017) );
  OAI22X1 U690 ( .A0(n1155), .A1(n414), .B0(n9), .B1(n413), .Y(n465) );
  NAND2X1 U691 ( .A(n324), .B(n323), .Y(n325) );
  OAI21XL U692 ( .A0(n5), .A1(n1227), .B0(n1234), .Y(n204) );
  XOR2X1 U693 ( .A(n329), .B(n62), .Y(PRODUCT[19]) );
  OAI21XL U694 ( .A0(n499), .A1(n449), .B0(n448), .Y(n451) );
  NOR2X1 U695 ( .A(n448), .B(n1288), .Y(n88) );
  INVX4 U696 ( .A(n59), .Y(n58) );
  NAND2X1 U697 ( .A(n564), .B(n563), .Y(n1091) );
  INVX8 U698 ( .A(n42), .Y(n1155) );
  OAI22XL U699 ( .A0(n908), .A1(n9), .B0(n950), .B1(n1155), .Y(n951) );
  OAI22XL U700 ( .A0(n840), .A1(n1155), .B0(n807), .B1(n9), .Y(n841) );
  AND2X4 U701 ( .A(n145), .B(n337), .Y(n42) );
  OAI2BB1X4 U702 ( .A0N(n37), .A1N(n421), .B0(n97), .Y(n59) );
  NAND2X1 U703 ( .A(n47), .B(n46), .Y(n1093) );
  XOR3X2 U704 ( .A(n1027), .B(n1025), .C(n1026), .Y(mult_x_1_n618) );
  INVXL U705 ( .A(n1027), .Y(n51) );
  NAND2XL U706 ( .A(n53), .B(n998), .Y(n52) );
  XNOR2X4 U707 ( .A(B[13]), .B(B[14]), .Y(n335) );
  NAND3X1 U708 ( .A(n59), .B(n85), .C(n91), .Y(n90) );
  INVX1 U709 ( .A(n449), .Y(n60) );
  NAND3X2 U710 ( .A(n60), .B(n61), .C(n1294), .Y(n87) );
  INVX1 U711 ( .A(n1288), .Y(n61) );
  XOR2X1 U712 ( .A(n955), .B(n1138), .Y(n66) );
  OAI21XL U713 ( .A0(n1102), .A1(n1101), .B0(n1100), .Y(n1107) );
  CMPR22X1 U714 ( .A(n633), .B(n632), .CO(n669), .S(n665) );
  BUFX12 U715 ( .A(n719), .Y(n1179) );
  OR2X2 U716 ( .A(n1074), .B(n1079), .Y(n71) );
  AOI21X1 U717 ( .A0(n68), .A1(n86), .B0(n78), .Y(n77) );
  XOR2X2 U718 ( .A(n81), .B(n38), .Y(PRODUCT[26]) );
  NAND2X1 U719 ( .A(n303), .B(n82), .Y(n81) );
  NAND2X1 U720 ( .A(n315), .B(n98), .Y(n83) );
  OAI21X1 U721 ( .A0(n109), .A1(n1069), .B0(n110), .Y(n315) );
  OAI21XL U722 ( .A0(n1076), .A1(n1071), .B0(n1077), .Y(n84) );
  NAND2X1 U723 ( .A(n1312), .B(n1311), .Y(n1071) );
  NAND3BX4 U724 ( .AN(n88), .B(n87), .C(n1289), .Y(n421) );
  NAND2X1 U725 ( .A(n98), .B(n314), .Y(n117) );
  AOI21X2 U726 ( .A0(n1263), .A1(n1260), .B0(n1261), .Y(n448) );
  XOR2X1 U727 ( .A(n318), .B(n420), .Y(PRODUCT[17]) );
  XOR2X2 U728 ( .A(n116), .B(n35), .Y(PRODUCT[30]) );
  XNOR3X2 U729 ( .A(n694), .B(n692), .C(n94), .Y(n722) );
  OAI22X2 U730 ( .A0(n1179), .A1(n906), .B0(n994), .B1(n872), .Y(n910) );
  OAI22X2 U731 ( .A0(n1179), .A1(n872), .B0(n994), .B1(n839), .Y(n875) );
  OAI22X1 U732 ( .A0(n1179), .A1(n839), .B0(n994), .B1(n806), .Y(n842) );
  OAI22X1 U733 ( .A0(n1179), .A1(n806), .B0(n994), .B1(n767), .Y(n809) );
  CMPR22X1 U734 ( .A(n398), .B(n397), .CO(n403), .S(n432) );
  NOR2X1 U735 ( .A(n1087), .B(n1086), .Y(n1103) );
  NAND2X1 U736 ( .A(n150), .B(n152), .Y(n339) );
  NOR2X1 U737 ( .A(n674), .B(n673), .Y(n1101) );
  BUFX4 U738 ( .A(B[5]), .Y(n926) );
  BUFX8 U739 ( .A(B[13]), .Y(n1140) );
  INVX8 U740 ( .A(n151), .Y(n955) );
  XNOR2X1 U741 ( .A(n920), .B(A[3]), .Y(n461) );
  XNOR2XL U742 ( .A(B[1]), .B(A[19]), .Y(n959) );
  XNOR2X1 U743 ( .A(n955), .B(A[6]), .Y(n404) );
  XNOR2XL U744 ( .A(B[7]), .B(A[25]), .Y(n148) );
  OAI22X1 U745 ( .A0(n948), .A1(n638), .B0(n7), .B1(n637), .Y(n639) );
  OAI22X1 U746 ( .A0(n972), .A1(n711), .B0(n970), .B1(n258), .Y(n700) );
  XNOR2XL U747 ( .A(n955), .B(A[19]), .Y(n715) );
  XNOR2XL U748 ( .A(n920), .B(n1138), .Y(n186) );
  OAI22X1 U749 ( .A0(n972), .A1(n258), .B0(n970), .B1(n207), .Y(n226) );
  OAI22X1 U750 ( .A0(n1179), .A1(n347), .B0(n994), .B1(n342), .Y(n378) );
  NOR2X1 U751 ( .A(n1311), .B(n1312), .Y(n317) );
  NOR2X1 U752 ( .A(n1309), .B(n1310), .Y(n1076) );
  NOR2X1 U753 ( .A(n1307), .B(n1308), .Y(n301) );
  NOR2X1 U754 ( .A(n1305), .B(n1306), .Y(n305) );
  OAI21XL U755 ( .A0(n322), .A1(n327), .B0(n323), .Y(n95) );
  AOI21X1 U756 ( .A0(n96), .A1(n319), .B0(n95), .Y(n97) );
  NAND2XL U757 ( .A(n1309), .B(n1310), .Y(n1077) );
  NAND2X1 U758 ( .A(n1307), .B(n1308), .Y(n310) );
  OAI21XL U759 ( .A0(n305), .A1(n310), .B0(n306), .Y(n119) );
  NAND2X1 U760 ( .A(n1303), .B(n1304), .Y(n289) );
  NAND2XL U761 ( .A(n1301), .B(n1302), .Y(n297) );
  OAI21XL U762 ( .A0(n296), .A1(n289), .B0(n297), .Y(n99) );
  AOI21XL U763 ( .A0(n100), .A1(n119), .B0(n99), .Y(n101) );
  NOR2X1 U764 ( .A(n1298), .B(n1297), .Y(n113) );
  NOR2XL U765 ( .A(n284), .B(n113), .Y(n278) );
  NOR2XL U766 ( .A(n239), .B(n1282), .Y(n104) );
  NOR2XL U767 ( .A(n1227), .B(n1280), .Y(n136) );
  INVXL U768 ( .A(n136), .Y(n106) );
  NAND2XL U769 ( .A(n1298), .B(n1297), .Y(n114) );
  OAI21XL U770 ( .A0(n113), .A1(n285), .B0(n114), .Y(n240) );
  NAND2XL U771 ( .A(n1295), .B(n1296), .Y(n280) );
  OAI21XL U772 ( .A0(n1282), .A1(n280), .B0(n1283), .Y(n103) );
  AOI21X1 U773 ( .A0(n240), .A1(n104), .B0(n103), .Y(n1234) );
  INVXL U774 ( .A(n109), .Y(n111) );
  OAI21X1 U775 ( .A0(n5), .A1(n284), .B0(n285), .Y(n116) );
  INVXL U776 ( .A(n118), .Y(n288) );
  NAND2XL U777 ( .A(n91), .B(n118), .Y(n121) );
  INVXL U778 ( .A(n119), .Y(n291) );
  INVXL U779 ( .A(n290), .Y(n122) );
  NAND2XL U780 ( .A(n138), .B(n142), .Y(n127) );
  NOR2XL U781 ( .A(n127), .B(n1280), .Y(n1226) );
  INVXL U782 ( .A(n1226), .Y(n129) );
  NAND2XL U783 ( .A(n1213), .B(n1190), .Y(n132) );
  OAI21XL U784 ( .A0(n127), .A1(n1281), .B0(n126), .Y(n1231) );
  AOI21XL U785 ( .A0(n1219), .A1(n1190), .B0(n130), .Y(n131) );
  OAI21XL U786 ( .A0(n5), .A1(n132), .B0(n131), .Y(n135) );
  NAND2XL U787 ( .A(n136), .B(n138), .Y(n141) );
  AOI21XL U788 ( .A0(n139), .A1(n138), .B0(n137), .Y(n140) );
  OAI21XL U789 ( .A0(n5), .A1(n141), .B0(n140), .Y(n144) );
  XOR2X1 U790 ( .A(B[12]), .B(B[13]), .Y(n145) );
  XNOR2X1 U791 ( .A(n1140), .B(n1138), .Y(n157) );
  CLKINVX3 U792 ( .A(n566), .Y(n870) );
  XNOR2X1 U793 ( .A(n870), .B(A[24]), .Y(n215) );
  OAI22X1 U794 ( .A0(n948), .A1(n215), .B0(n7), .B1(n148), .Y(n191) );
  XNOR2X1 U795 ( .A(B[15]), .B(n883), .Y(n160) );
  XNOR2X1 U796 ( .A(B[15]), .B(A[19]), .Y(n156) );
  OAI22XL U797 ( .A0(n1179), .A1(n160), .B0(n1180), .B1(n156), .Y(n164) );
  XNOR2X1 U798 ( .A(n920), .B(n1156), .Y(n158) );
  OAI22XL U799 ( .A0(n1119), .A1(n181), .B0(n10), .B1(n158), .Y(n163) );
  XOR2X1 U800 ( .A(B[8]), .B(B[9]), .Y(n150) );
  XNOR2X1 U801 ( .A(B[8]), .B(B[7]), .Y(n152) );
  XNOR2X1 U802 ( .A(n955), .B(A[24]), .Y(n159) );
  BUFX8 U803 ( .A(n152), .Y(n1001) );
  XNOR2X1 U804 ( .A(n955), .B(A[25]), .Y(n154) );
  XNOR2X1 U805 ( .A(B[16]), .B(n883), .Y(n153) );
  XNOR2X1 U806 ( .A(B[15]), .B(n1115), .Y(n168) );
  XNOR2X1 U807 ( .A(n955), .B(n1156), .Y(n183) );
  XNOR2X1 U808 ( .A(B[15]), .B(n922), .Y(n185) );
  OAI22XL U809 ( .A0(n1179), .A1(n185), .B0(n1180), .B1(n160), .Y(n188) );
  CMPR32X1 U810 ( .A(n164), .B(n163), .C(n162), .CO(n180), .S(n197) );
  CMPR32X1 U811 ( .A(n167), .B(n166), .C(n165), .CO(n201), .S(n196) );
  XNOR2X1 U812 ( .A(B[15]), .B(n1138), .Y(n1121) );
  XNOR2XL U813 ( .A(n920), .B(A[25]), .Y(n1117) );
  OAI22X1 U814 ( .A0(n1119), .A1(n170), .B0(n10), .B1(n1117), .Y(n1135) );
  XNOR2X1 U815 ( .A(n1140), .B(n1156), .Y(n1120) );
  CMPR32X1 U816 ( .A(n174), .B(n173), .C(n172), .CO(n1126), .S(n179) );
  CMPR32X1 U817 ( .A(n177), .B(n176), .C(n175), .CO(n1125), .S(n178) );
  CMPR32X1 U818 ( .A(n180), .B(n179), .C(n178), .CO(n1112), .S(n200) );
  NAND2XL U819 ( .A(n1109), .B(n1108), .Y(mult_x_1_n152) );
  XNOR2X1 U820 ( .A(n955), .B(n1151), .Y(n217) );
  XNOR2X1 U821 ( .A(n949), .B(n885), .Y(n216) );
  CMPR32X1 U822 ( .A(n189), .B(n188), .C(n187), .CO(n198), .S(n233) );
  CMPR32X1 U823 ( .A(n192), .B(n191), .C(n190), .CO(n165), .S(n232) );
  ADDFHX1 U824 ( .A(n195), .B(n194), .CI(n193), .CO(n236), .S(n231) );
  CMPR32X1 U825 ( .A(n198), .B(n197), .C(n196), .CO(n199), .S(n234) );
  CMPR32X1 U826 ( .A(n201), .B(n200), .C(n199), .CO(n1109), .S(n1110) );
  NAND2XL U827 ( .A(n1111), .B(n1110), .Y(mult_x_1_n161) );
  XNOR2X1 U828 ( .A(n204), .B(n203), .Y(PRODUCT[33]) );
  XOR2X1 U829 ( .A(B[4]), .B(B[5]), .Y(n206) );
  XNOR2X1 U830 ( .A(B[4]), .B(B[3]), .Y(n360) );
  BUFX3 U831 ( .A(n360), .Y(n970) );
  CMPR32X1 U832 ( .A(n214), .B(n213), .C(n212), .CO(n194), .S(n247) );
  XNOR2X1 U833 ( .A(n870), .B(n1156), .Y(n222) );
  INVX8 U834 ( .A(n344), .Y(n949) );
  XNOR2X1 U835 ( .A(n949), .B(n925), .Y(n223) );
  INVXL U836 ( .A(n226), .Y(n264) );
  XNOR2X1 U837 ( .A(n870), .B(n1151), .Y(n260) );
  CMPR32X1 U838 ( .A(n230), .B(n229), .C(n228), .CO(n272), .S(n686) );
  CMPR32X1 U839 ( .A(n233), .B(n232), .C(n231), .CO(n235), .S(n273) );
  CMPR32X1 U840 ( .A(n236), .B(n235), .C(n234), .CO(n1111), .S(n237) );
  NOR2XL U841 ( .A(n238), .B(n237), .Y(mult_x_1_n169) );
  NAND2XL U842 ( .A(n238), .B(n237), .Y(mult_x_1_n170) );
  NAND2XL U843 ( .A(n278), .B(n281), .Y(n244) );
  INVXL U844 ( .A(n240), .Y(n241) );
  INVXL U845 ( .A(n280), .Y(n242) );
  AOI21XL U846 ( .A0(n240), .A1(n281), .B0(n242), .Y(n243) );
  OAI21XL U847 ( .A0(n5), .A1(n244), .B0(n243), .Y(n246) );
  CMPR32X1 U848 ( .A(n249), .B(n248), .C(n247), .CO(n275), .S(n685) );
  CMPR32X1 U849 ( .A(n252), .B(n251), .C(n250), .CO(n271), .S(n691) );
  XNOR2XL U850 ( .A(B[16]), .B(n912), .Y(n253) );
  XNOR2X1 U851 ( .A(B[2]), .B(B[1]), .Y(n255) );
  OAI22X1 U852 ( .A0(n968), .A1(n724), .B0(n255), .B1(n256), .Y(n713) );
  INVXL U853 ( .A(n256), .Y(n257) );
  XNOR2X1 U854 ( .A(n949), .B(n946), .Y(n697) );
  XNOR2X1 U855 ( .A(n870), .B(n1138), .Y(n695) );
  XNOR2X1 U856 ( .A(n920), .B(n922), .Y(n716) );
  OAI22XL U857 ( .A0(n1119), .A1(n716), .B0(n10), .B1(n263), .Y(n701) );
  CMPR32X1 U858 ( .A(n275), .B(n274), .C(n273), .CO(n238), .S(n276) );
  NOR2XL U859 ( .A(n277), .B(n276), .Y(mult_x_1_n176) );
  NAND2XL U860 ( .A(n277), .B(n276), .Y(mult_x_1_n177) );
  INVXL U861 ( .A(n278), .Y(n279) );
  NAND2X1 U862 ( .A(n281), .B(n280), .Y(n282) );
  NOR2XL U863 ( .A(n288), .B(n290), .Y(n293) );
  NAND2XL U864 ( .A(n293), .B(n91), .Y(n295) );
  OAI21XL U865 ( .A0(n291), .A1(n290), .B0(n289), .Y(n292) );
  AOI21XL U866 ( .A0(n308), .A1(n293), .B0(n292), .Y(n294) );
  OAI21X1 U867 ( .A0(n295), .A1(n58), .B0(n294), .Y(n300) );
  INVXL U868 ( .A(n296), .Y(n298) );
  XNOR2X2 U869 ( .A(n300), .B(n299), .Y(PRODUCT[28]) );
  NAND2XL U870 ( .A(n91), .B(n311), .Y(n304) );
  INVXL U871 ( .A(n310), .Y(n302) );
  AOI21XL U872 ( .A0(n308), .A1(n311), .B0(n302), .Y(n303) );
  INVXL U873 ( .A(n308), .Y(n309) );
  NAND2XL U874 ( .A(n311), .B(n310), .Y(n312) );
  INVXL U875 ( .A(n315), .Y(n316) );
  INVX1 U876 ( .A(n317), .Y(n1073) );
  INVXL U877 ( .A(n322), .Y(n324) );
  INVXL U878 ( .A(n321), .Y(n328) );
  NAND2XL U879 ( .A(n328), .B(n327), .Y(n329) );
  INVX1 U880 ( .A(n1286), .Y(n331) );
  INVXL U881 ( .A(n1284), .Y(n332) );
  NAND2X1 U882 ( .A(n332), .B(n1285), .Y(n333) );
  XOR2X1 U883 ( .A(n334), .B(n333), .Y(PRODUCT[18]) );
  XNOR2X1 U884 ( .A(n949), .B(n585), .Y(n347) );
  XNOR2X1 U885 ( .A(n949), .B(A[3]), .Y(n342) );
  XNOR2XL U886 ( .A(B[16]), .B(A[1]), .Y(n336) );
  NOR2XL U887 ( .A(n1176), .B(n336), .Y(n377) );
  XNOR2X1 U888 ( .A(B[7]), .B(A[10]), .Y(n368) );
  XNOR2X1 U889 ( .A(B[7]), .B(n954), .Y(n388) );
  OAI22XL U890 ( .A0(n948), .A1(n368), .B0(n7), .B1(n388), .Y(n381) );
  XNOR2X1 U891 ( .A(n955), .B(n907), .Y(n353) );
  BUFX3 U892 ( .A(n636), .Y(n961) );
  XNOR2X1 U893 ( .A(B[1]), .B(n885), .Y(n345) );
  XNOR2X1 U894 ( .A(B[1]), .B(n922), .Y(n389) );
  BUFX3 U895 ( .A(n814), .Y(n1066) );
  BUFX3 U896 ( .A(A[0]), .Y(n1067) );
  OAI22X1 U897 ( .A0(n1119), .A1(n357), .B0(n10), .B1(n964), .Y(n1009) );
  XNOR2X1 U898 ( .A(n949), .B(n917), .Y(n995) );
  XNOR2X1 U899 ( .A(B[1]), .B(A[14]), .Y(n399) );
  XNOR2X1 U900 ( .A(B[1]), .B(n925), .Y(n346) );
  OAI22X1 U901 ( .A0(n961), .A1(n399), .B0(n346), .B1(n1066), .Y(n398) );
  XNOR2X1 U902 ( .A(n949), .B(A[1]), .Y(n348) );
  XNOR2X1 U903 ( .A(n955), .B(A[7]), .Y(n354) );
  XNOR2X1 U904 ( .A(n949), .B(n1067), .Y(n349) );
  CMPR32X1 U905 ( .A(n352), .B(n351), .C(n350), .CO(n372), .S(n402) );
  OAI22X1 U906 ( .A0(n41), .A1(n361), .B0(n966), .B1(n359), .Y(n363) );
  OAI22XL U907 ( .A0(n1155), .A1(n356), .B0(n9), .B1(n355), .Y(n362) );
  XNOR2X1 U908 ( .A(n920), .B(A[6]), .Y(n366) );
  XNOR2X1 U909 ( .A(n920), .B(n917), .Y(n405) );
  XNOR2X1 U910 ( .A(n920), .B(A[5]), .Y(n367) );
  XNOR2X1 U911 ( .A(B[7]), .B(n907), .Y(n411) );
  XNOR2X1 U912 ( .A(B[7]), .B(n919), .Y(n369) );
  ADDFHX1 U913 ( .A(n372), .B(n371), .CI(n370), .CO(n1056), .S(n416) );
  CMPR32X1 U914 ( .A(n375), .B(n374), .C(n373), .CO(n395), .S(n425) );
  CMPR32X1 U915 ( .A(n378), .B(n377), .C(n376), .CO(n1053), .S(n394) );
  XNOR2X1 U916 ( .A(n955), .B(A[10]), .Y(n1002) );
  OAI22XL U917 ( .A0(n972), .A1(n386), .B0(n970), .B1(n971), .Y(n1029) );
  XNOR2X1 U918 ( .A(B[7]), .B(n912), .Y(n992) );
  OAI22XL U919 ( .A0(n948), .A1(n388), .B0(n7), .B1(n992), .Y(n1035) );
  XNOR2X1 U920 ( .A(B[1]), .B(n883), .Y(n960) );
  OAI22X1 U921 ( .A0(n961), .A1(n389), .B0(n960), .B1(n814), .Y(n1006) );
  XNOR2XL U922 ( .A(B[16]), .B(n585), .Y(n390) );
  ADDHXL U923 ( .A(n392), .B(n391), .CO(n1033), .S(n379) );
  XNOR2X1 U924 ( .A(B[1]), .B(n946), .Y(n412) );
  OAI22XL U925 ( .A0(n961), .A1(n412), .B0(n399), .B1(n1066), .Y(n435) );
  XNOR2X1 U926 ( .A(n955), .B(A[5]), .Y(n437) );
  XNOR2X1 U927 ( .A(n870), .B(A[7]), .Y(n458) );
  XNOR2X1 U928 ( .A(B[1]), .B(n912), .Y(n467) );
  NAND2XL U929 ( .A(n419), .B(n418), .Y(mult_x_1_n282) );
  NAND2X1 U930 ( .A(n331), .B(n1287), .Y(n420) );
  CMPR32X1 U931 ( .A(n430), .B(n429), .C(n428), .CO(n427), .S(n474) );
  CMPR32X1 U932 ( .A(n433), .B(n432), .C(n431), .CO(n445), .S(n473) );
  CMPR32X1 U933 ( .A(n436), .B(n435), .C(n434), .CO(n431), .S(n482) );
  NOR2XL U934 ( .A(n447), .B(n446), .Y(mult_x_1_n286) );
  NAND2XL U935 ( .A(n447), .B(n446), .Y(mult_x_1_n287) );
  NAND2XL U936 ( .A(n61), .B(n1289), .Y(n450) );
  XNOR2X1 U937 ( .A(n451), .B(n450), .Y(PRODUCT[16]) );
  CMPR32X1 U938 ( .A(n454), .B(n453), .C(n452), .CO(n446), .S(n476) );
  OAI22XL U939 ( .A0(n948), .A1(n469), .B0(n7), .B1(n458), .Y(n485) );
  XNOR2X1 U940 ( .A(n920), .B(n585), .Y(n468) );
  XNOR2X1 U941 ( .A(B[1]), .B(n954), .Y(n490) );
  XNOR2X1 U942 ( .A(n920), .B(A[1]), .Y(n507) );
  XNOR2X1 U943 ( .A(n870), .B(A[5]), .Y(n506) );
  OAI22XL U944 ( .A0(n948), .A1(n506), .B0(n7), .B1(n469), .Y(n515) );
  NOR2XL U945 ( .A(n476), .B(n475), .Y(mult_x_1_n292) );
  NAND2XL U946 ( .A(n476), .B(n475), .Y(mult_x_1_n293) );
  ADDFHX1 U947 ( .A(n482), .B(n481), .CI(n480), .CO(n472), .S(n502) );
  CMPR32X1 U948 ( .A(n485), .B(n484), .C(n483), .CO(n498), .S(n518) );
  XNOR2X1 U949 ( .A(n955), .B(A[3]), .Y(n511) );
  XNOR2XL U950 ( .A(B[1]), .B(A[10]), .Y(n527) );
  CMPR32X1 U951 ( .A(n498), .B(n497), .C(n496), .CO(n478), .S(n500) );
  NAND2XL U952 ( .A(n1098), .B(n1097), .Y(n1099) );
  INVXL U953 ( .A(n1099), .Y(mult_x_1_n298) );
  CMPR32X1 U954 ( .A(n502), .B(n501), .C(n500), .CO(n1097), .S(n521) );
  XNOR2X1 U955 ( .A(n870), .B(n917), .Y(n529) );
  OAI22XL U956 ( .A0(n948), .A1(n529), .B0(n7), .B1(n506), .Y(n534) );
  CMPR32X1 U957 ( .A(n515), .B(n514), .C(n513), .CO(n503), .S(n535) );
  NOR2XL U958 ( .A(n521), .B(n520), .Y(n519) );
  INVXL U959 ( .A(n519), .Y(mult_x_1_n304) );
  NAND2XL U960 ( .A(n521), .B(n520), .Y(n522) );
  INVXL U961 ( .A(n522), .Y(mult_x_1_n305) );
  NAND2XL U962 ( .A(mult_x_1_n304), .B(n522), .Y(mult_x_1_n84) );
  CMPR32X1 U963 ( .A(n526), .B(n525), .C(n524), .CO(n516), .S(n562) );
  OAI22XL U964 ( .A0(n636), .A1(n541), .B0(n527), .B1(n1066), .Y(n544) );
  XNOR2X1 U965 ( .A(n955), .B(A[1]), .Y(n547) );
  XNOR2X1 U966 ( .A(B[7]), .B(A[3]), .Y(n546) );
  OAI22X1 U967 ( .A0(n948), .A1(n546), .B0(n7), .B1(n529), .Y(n663) );
  CMPR32X1 U968 ( .A(n534), .B(n533), .C(n532), .CO(n537), .S(n551) );
  CMPR32X1 U969 ( .A(n540), .B(n539), .C(n538), .CO(n536), .S(n1082) );
  XNOR2XL U970 ( .A(B[1]), .B(n907), .Y(n634) );
  OAI22X1 U971 ( .A0(n948), .A1(n637), .B0(n7), .B1(n546), .Y(n623) );
  OAI22X1 U972 ( .A0(n8), .A1(n548), .B0(n1001), .B1(n547), .Y(n622) );
  OAI22X1 U973 ( .A0(n550), .A1(n626), .B0(n970), .B1(n549), .Y(n621) );
  ADDFHX1 U974 ( .A(n553), .B(n552), .CI(n551), .CO(n561), .S(n1080) );
  NOR2XL U975 ( .A(n556), .B(n555), .Y(n554) );
  INVXL U976 ( .A(n554), .Y(mult_x_1_n317) );
  INVXL U977 ( .A(n1128), .Y(mult_x_1_n318) );
  ADDFHX1 U978 ( .A(n559), .B(n558), .CI(n557), .CO(n520), .S(n564) );
  NAND2XL U979 ( .A(n1093), .B(n1091), .Y(mult_x_1_n85) );
  XNOR2X1 U980 ( .A(n1266), .B(n1293), .Y(PRODUCT[12]) );
  XNOR2X1 U981 ( .A(B[1]), .B(A[6]), .Y(n567) );
  XNOR2X1 U982 ( .A(B[1]), .B(A[7]), .Y(n635) );
  OAI22XL U983 ( .A0(n948), .A1(n566), .B0(n7), .B1(n565), .Y(n628) );
  NOR2BX1 U984 ( .AN(n1067), .B(n7), .Y(n576) );
  XNOR2X1 U985 ( .A(B[1]), .B(A[5]), .Y(n571) );
  OAI22X1 U986 ( .A0(n961), .A1(n571), .B0(n567), .B1(n1066), .Y(n575) );
  OAI22X1 U987 ( .A0(n968), .A1(n570), .B0(n966), .B1(n625), .Y(n644) );
  XNOR2X1 U988 ( .A(B[7]), .B(n1067), .Y(n568) );
  XNOR2X1 U989 ( .A(n870), .B(A[1]), .Y(n638) );
  OAI22X1 U990 ( .A0(n948), .A1(n568), .B0(n7), .B1(n638), .Y(n643) );
  XNOR2X1 U991 ( .A(B[1]), .B(n917), .Y(n597) );
  OAI22X1 U992 ( .A0(n961), .A1(n597), .B0(n571), .B1(n1066), .Y(n584) );
  OAI22X1 U993 ( .A0(n972), .A1(n573), .B0(n970), .B1(n572), .Y(n583) );
  CMPR32X1 U994 ( .A(n579), .B(n578), .C(n577), .CO(n617), .S(n616) );
  NOR2XL U995 ( .A(n1202), .B(n1207), .Y(n620) );
  XNOR2X1 U996 ( .A(B[1]), .B(A[1]), .Y(n586) );
  XNOR2X1 U997 ( .A(B[1]), .B(n585), .Y(n591) );
  XNOR2X1 U998 ( .A(B[1]), .B(A[3]), .Y(n598) );
  OAI22X1 U999 ( .A0(n961), .A1(n591), .B0(n598), .B1(n1066), .Y(n602) );
  OAI22X1 U1000 ( .A0(n41), .A1(n592), .B0(n966), .B1(n600), .Y(n601) );
  OAI21XL U1001 ( .A0(n1245), .A1(n1242), .B0(n1243), .Y(n1240) );
  CMPR22X1 U1002 ( .A(n602), .B(n601), .CO(n604), .S(n596) );
  CMPR32X1 U1003 ( .A(n609), .B(n608), .C(n607), .CO(n615), .S(n614) );
  CMPR32X1 U1004 ( .A(n612), .B(n611), .C(n610), .CO(n613), .S(n605) );
  OAI21XL U1005 ( .A0(n1258), .A1(n1255), .B0(n1256), .Y(n1201) );
  NAND2XL U1006 ( .A(n618), .B(n617), .Y(n1203) );
  OAI21XL U1007 ( .A0(n1202), .A1(n1208), .B0(n1203), .Y(n619) );
  AOI21XL U1008 ( .A0(n620), .A1(n1201), .B0(n619), .Y(n677) );
  ADDHXL U1009 ( .A(n629), .B(n628), .CO(n645), .S(n653) );
  OAI22XL U1010 ( .A0(n636), .A1(n635), .B0(n634), .B1(n1066), .Y(n640) );
  CMPR32X1 U1011 ( .A(n641), .B(n640), .C(n639), .CO(n664), .S(n650) );
  OR2X2 U1012 ( .A(n657), .B(n656), .Y(n680) );
  CMPR32X1 U1013 ( .A(n650), .B(n649), .C(n648), .CO(n656), .S(n655) );
  CMPR32X1 U1014 ( .A(n40), .B(n652), .C(n651), .CO(n654), .S(n618) );
  OR2X2 U1015 ( .A(n655), .B(n654), .Y(n1194) );
  NAND2X1 U1016 ( .A(n680), .B(n1194), .Y(n660) );
  NAND2XL U1017 ( .A(n655), .B(n654), .Y(n1193) );
  INVXL U1018 ( .A(n1193), .Y(n678) );
  NAND2XL U1019 ( .A(n657), .B(n656), .Y(n679) );
  INVXL U1020 ( .A(n679), .Y(n658) );
  AOI21X1 U1021 ( .A0(n680), .A1(n678), .B0(n658), .Y(n659) );
  OAI21X1 U1022 ( .A0(n677), .A1(n660), .B0(n659), .Y(n1090) );
  CMPR32X1 U1023 ( .A(n663), .B(n662), .C(n661), .CO(n552), .S(n1085) );
  CMPR32X1 U1024 ( .A(n666), .B(n665), .C(n664), .CO(n1084), .S(n670) );
  INVXL U1025 ( .A(n1101), .Y(n675) );
  NAND2XL U1026 ( .A(n675), .B(n1100), .Y(n676) );
  XOR2X1 U1027 ( .A(n1102), .B(n676), .Y(n1335) );
  INVXL U1028 ( .A(n677), .Y(n1196) );
  AOI21XL U1029 ( .A0(n1196), .A1(n1194), .B0(n678), .Y(n682) );
  ADDFHX1 U1030 ( .A(n685), .B(n684), .CI(n683), .CO(n277), .S(mult_x_1_n470)
         );
  CMPR32X1 U1031 ( .A(n691), .B(n690), .C(n689), .CO(n684), .S(n708) );
  XNOR2X1 U1032 ( .A(n870), .B(n1115), .Y(n717) );
  OAI22X1 U1033 ( .A0(n948), .A1(n717), .B0(n7), .B1(n695), .Y(n746) );
  XNOR2XL U1034 ( .A(B[16]), .B(n954), .Y(n696) );
  NOR2XL U1035 ( .A(n1176), .B(n696), .Y(n745) );
  XNOR2X1 U1036 ( .A(n949), .B(n912), .Y(n718) );
  OAI22XL U1037 ( .A0(n719), .A1(n718), .B0(n994), .B1(n697), .Y(n744) );
  CMPR32X1 U1038 ( .A(n703), .B(n702), .C(n701), .CO(n706), .S(n732) );
  CMPR32X1 U1039 ( .A(n706), .B(n705), .C(n704), .CO(n689), .S(n720) );
  CMPR32X1 U1040 ( .A(n709), .B(n708), .C(n707), .CO(mult_x_1_n481), .S(
        mult_x_1_n482) );
  OAI22XL U1041 ( .A0(n1155), .A1(n743), .B0(n9), .B1(n710), .Y(n728) );
  XNOR2X1 U1042 ( .A(n926), .B(n1151), .Y(n741) );
  INVXL U1043 ( .A(n713), .Y(n726) );
  CMPR32X1 U1044 ( .A(n714), .B(n713), .C(n712), .CO(n693), .S(n736) );
  XNOR2X1 U1045 ( .A(n955), .B(n883), .Y(n747) );
  XNOR2X1 U1046 ( .A(n920), .B(n885), .Y(n723) );
  OAI22XL U1047 ( .A0(n1119), .A1(n723), .B0(n10), .B1(n716), .Y(n730) );
  XNOR2X1 U1048 ( .A(n870), .B(A[19]), .Y(n766) );
  XNOR2X1 U1049 ( .A(n949), .B(n954), .Y(n767) );
  OAI22X1 U1050 ( .A0(n719), .A1(n767), .B0(n994), .B1(n718), .Y(n750) );
  ADDFHX1 U1051 ( .A(n722), .B(n721), .CI(n720), .CO(n707), .S(n739) );
  CMPR32X1 U1052 ( .A(n728), .B(n727), .C(n726), .CO(n737), .S(n782) );
  CMPR32X1 U1053 ( .A(n731), .B(n730), .C(n729), .CO(n735), .S(n781) );
  CMPR32X1 U1054 ( .A(n734), .B(n733), .C(n732), .CO(n721), .S(n776) );
  CMPR32X1 U1055 ( .A(n737), .B(n736), .C(n735), .CO(n740), .S(n775) );
  CMPR32X1 U1056 ( .A(n740), .B(n739), .C(n738), .CO(mult_x_1_n493), .S(
        mult_x_1_n494) );
  XNOR2XL U1057 ( .A(B[16]), .B(A[10]), .Y(n742) );
  NOR2XL U1058 ( .A(n1176), .B(n742), .Y(n770) );
  XNOR2X1 U1059 ( .A(n955), .B(n922), .Y(n758) );
  XNOR2X1 U1060 ( .A(B[1]), .B(A[24]), .Y(n761) );
  OAI22X1 U1061 ( .A0(n961), .A1(n761), .B0(n748), .B1(n1066), .Y(n760) );
  XNOR2XL U1062 ( .A(B[16]), .B(n919), .Y(n749) );
  XNOR2X1 U1063 ( .A(n955), .B(n885), .Y(n811) );
  XNOR2X1 U1064 ( .A(B[1]), .B(n1156), .Y(n815) );
  OAI22X1 U1065 ( .A0(n961), .A1(n815), .B0(n761), .B1(n814), .Y(n813) );
  XNOR2XL U1066 ( .A(B[16]), .B(n907), .Y(n762) );
  NOR2XL U1067 ( .A(n1176), .B(n762), .Y(n812) );
  CMPR32X1 U1068 ( .A(n765), .B(n764), .C(n763), .CO(n780), .S(n800) );
  XNOR2X1 U1069 ( .A(n870), .B(n883), .Y(n805) );
  OAI22X1 U1070 ( .A0(n948), .A1(n805), .B0(n7), .B1(n766), .Y(n810) );
  XNOR2X1 U1071 ( .A(n949), .B(A[10]), .Y(n806) );
  CMPR32X1 U1072 ( .A(n771), .B(n770), .C(n769), .CO(n765), .S(n797) );
  CMPR32X1 U1073 ( .A(n774), .B(n773), .C(n772), .CO(n763), .S(n796) );
  CMPR32X1 U1074 ( .A(n777), .B(n776), .C(n775), .CO(n738), .S(n778) );
  ADDFHX1 U1075 ( .A(n780), .B(n779), .CI(n778), .CO(mult_x_1_n507), .S(
        mult_x_1_n508) );
  CMPR32X1 U1076 ( .A(n783), .B(n782), .C(n781), .CO(n777), .S(n804) );
  CMPR32X1 U1077 ( .A(n792), .B(n791), .C(n790), .CO(n793), .S(n829) );
  CMPR32X1 U1078 ( .A(n798), .B(n797), .C(n796), .CO(n799), .S(n832) );
  XNOR2X1 U1079 ( .A(n870), .B(n922), .Y(n838) );
  OAI22X1 U1080 ( .A0(n948), .A1(n838), .B0(n7), .B1(n805), .Y(n843) );
  XNOR2X1 U1081 ( .A(n949), .B(n919), .Y(n839) );
  XNOR2X1 U1082 ( .A(B[1]), .B(n1151), .Y(n847) );
  XNOR2XL U1083 ( .A(B[16]), .B(A[7]), .Y(n816) );
  NOR2XL U1084 ( .A(n1176), .B(n816), .Y(n845) );
  CMPR32X1 U1085 ( .A(n825), .B(n824), .C(n823), .CO(n826), .S(n861) );
  CMPR32X1 U1086 ( .A(n828), .B(n827), .C(n826), .CO(n837), .S(n865) );
  XNOR2X1 U1087 ( .A(n870), .B(n885), .Y(n871) );
  OAI22X1 U1088 ( .A0(n948), .A1(n871), .B0(n7), .B1(n838), .Y(n876) );
  XNOR2X1 U1089 ( .A(n949), .B(n907), .Y(n872) );
  XNOR2X1 U1090 ( .A(n955), .B(A[14]), .Y(n877) );
  ADDHXL U1091 ( .A(n846), .B(n845), .CO(n823), .S(n856) );
  OAI22X1 U1092 ( .A0(n961), .A1(n880), .B0(n847), .B1(n1066), .Y(n879) );
  XNOR2XL U1093 ( .A(B[16]), .B(A[6]), .Y(n848) );
  CMPR32X1 U1094 ( .A(n857), .B(n855), .C(n856), .CO(n858), .S(n896) );
  CMPR32X1 U1095 ( .A(n860), .B(n859), .C(n858), .CO(n869), .S(n900) );
  XNOR2X1 U1096 ( .A(n870), .B(n925), .Y(n905) );
  OAI22X1 U1097 ( .A0(n948), .A1(n905), .B0(n7), .B1(n871), .Y(n911) );
  XNOR2X1 U1098 ( .A(n949), .B(A[7]), .Y(n906) );
  XNOR2X1 U1099 ( .A(B[1]), .B(n1115), .Y(n916) );
  XNOR2XL U1100 ( .A(B[16]), .B(A[5]), .Y(n881) );
  NOR2XL U1101 ( .A(n1176), .B(n881), .Y(n914) );
  CMPR32X1 U1102 ( .A(n892), .B(n891), .C(n890), .CO(n893), .S(n937) );
  CMPR32X1 U1103 ( .A(n895), .B(n894), .C(n893), .CO(n904), .S(n941) );
  OAI22X1 U1104 ( .A0(n948), .A1(n947), .B0(n7), .B1(n905), .Y(n953) );
  XNOR2X1 U1105 ( .A(n1140), .B(n907), .Y(n950) );
  XNOR2X1 U1106 ( .A(n955), .B(n912), .Y(n956) );
  ADDHXL U1107 ( .A(n915), .B(n914), .CO(n890), .S(n932) );
  OAI22X1 U1108 ( .A0(n961), .A1(n959), .B0(n916), .B1(n1066), .Y(n958) );
  XNOR2XL U1109 ( .A(B[16]), .B(n917), .Y(n918) );
  CMPR32X1 U1110 ( .A(n933), .B(n931), .C(n932), .CO(n934), .S(n982) );
  CMPR32X1 U1111 ( .A(n936), .B(n935), .C(n934), .CO(n945), .S(n986) );
  XNOR2X1 U1112 ( .A(B[7]), .B(n946), .Y(n991) );
  XNOR2X1 U1113 ( .A(n1140), .B(A[7]), .Y(n996) );
  OAI22X1 U1114 ( .A0(n1155), .A1(n996), .B0(n9), .B1(n950), .Y(n998) );
  XNOR2XL U1115 ( .A(B[16]), .B(A[3]), .Y(n962) );
  NOR2XL U1116 ( .A(n1176), .B(n962), .Y(n1003) );
  CMPR32X1 U1117 ( .A(n978), .B(n977), .C(n976), .CO(n979), .S(n1019) );
  CMPR32X1 U1118 ( .A(n981), .B(n980), .C(n979), .CO(n990), .S(n1023) );
  OAI22X1 U1119 ( .A0(n948), .A1(n992), .B0(n7), .B1(n991), .Y(n1032) );
  ADDHXL U1120 ( .A(n1004), .B(n1003), .CO(n976), .S(n1014) );
  CMPR32X1 U1121 ( .A(n1009), .B(n1008), .C(n1007), .CO(n1044), .S(n1051) );
  CMPR32X1 U1122 ( .A(n1015), .B(n1013), .C(n1014), .CO(n1016), .S(n1042) );
  CMPR32X1 U1123 ( .A(n1018), .B(n1017), .C(n1016), .CO(n1027), .S(n1046) );
  CMPR32X1 U1124 ( .A(n1030), .B(n1029), .C(n1028), .CO(n1041), .S(n1037) );
  CMPR32X1 U1125 ( .A(n1035), .B(n1034), .C(n1033), .CO(n1039), .S(n1036) );
  CMPR32X1 U1126 ( .A(n1062), .B(n1061), .C(n1060), .CO(mult_x_1_n649), .S(
        mult_x_1_n650) );
  NAND2XL U1127 ( .A(n86), .B(n1069), .Y(n1070) );
  INVXL U1128 ( .A(n1071), .Y(n1072) );
  AOI21XL U1129 ( .A0(n315), .A1(n1073), .B0(n1072), .Y(n1074) );
  INVXL U1130 ( .A(n1076), .Y(n1078) );
  NAND2XL U1131 ( .A(n1078), .B(n1077), .Y(n1079) );
  NOR2XL U1132 ( .A(n1103), .B(n1101), .Y(n1089) );
  OAI21XL U1133 ( .A0(n1103), .A1(n1100), .B0(n1104), .Y(n1088) );
  AOI21XL U1134 ( .A0(n1090), .A1(n1089), .B0(n1088), .Y(n1096) );
  NAND2XL U1135 ( .A(n1093), .B(mult_x_1_n317), .Y(n1095) );
  INVXL U1136 ( .A(n1091), .Y(n1092) );
  AOI21XL U1137 ( .A0(n1093), .A1(mult_x_1_n318), .B0(n1092), .Y(n1094) );
  OAI21XL U1138 ( .A0(n1096), .A1(n1095), .B0(n1094), .Y(mult_x_1_n309) );
  INVXL U1139 ( .A(n1096), .Y(mult_x_1_n321) );
  OR2X2 U1140 ( .A(n1098), .B(n1097), .Y(n1321) );
  NAND2XL U1141 ( .A(n1321), .B(n1099), .Y(mult_x_1_n83) );
  INVXL U1142 ( .A(n1103), .Y(n1105) );
  NAND2XL U1143 ( .A(n1105), .B(n1104), .Y(n1106) );
  XNOR2X1 U1144 ( .A(n1107), .B(n1106), .Y(n1334) );
  CMPR32X1 U1145 ( .A(n1114), .B(n1113), .C(n1112), .CO(n1130), .S(n1108) );
  CMPR32X1 U1146 ( .A(n1124), .B(n1123), .C(n1122), .CO(n1142), .S(n1114) );
  CMPR32X1 U1147 ( .A(n1127), .B(n1126), .C(n1125), .CO(n1131), .S(n1113) );
  NAND2XL U1148 ( .A(mult_x_1_n317), .B(n1128), .Y(mult_x_1_n86) );
  CMPR32X1 U1149 ( .A(n1133), .B(n1132), .C(n1131), .CO(n1146), .S(n1129) );
  CMPR32X1 U1150 ( .A(n1136), .B(n1135), .C(n1134), .CO(n1164), .S(n1133) );
  XNOR2X1 U1151 ( .A(B[15]), .B(n1156), .Y(n1147) );
  XNOR2XL U1152 ( .A(n1140), .B(A[25]), .Y(n1153) );
  OAI22X1 U1153 ( .A0(n1155), .A1(n1141), .B0(n9), .B1(n1153), .Y(n1161) );
  CMPR32X1 U1154 ( .A(n1144), .B(n1143), .C(n1142), .CO(n1162), .S(n1132) );
  CMPR32X1 U1155 ( .A(n1150), .B(n1149), .C(n1148), .CO(n1166), .S(n1163) );
  CMPR32X1 U1156 ( .A(n1161), .B(n1160), .C(n1159), .CO(n1172), .S(n1165) );
  CMPR32X1 U1157 ( .A(n1164), .B(n1163), .C(n1162), .CO(n1171), .S(n1145) );
  CMPR32X1 U1158 ( .A(n1167), .B(n1166), .C(n1165), .CO(n1169), .S(n1170) );
  CMPR32X1 U1159 ( .A(n1174), .B(n1173), .C(n1172), .CO(n1185), .S(n1168) );
  OAI2BB1X1 U1160 ( .A0N(n1180), .A1N(n1179), .B0(n1178), .Y(n1181) );
  XOR3X2 U1161 ( .A(n1183), .B(n1182), .C(n1181), .Y(n1184) );
  OAI21XL U1162 ( .A0(n5), .A1(n1189), .B0(n1188), .Y(n1192) );
  XNOR2X1 U1163 ( .A(n1192), .B(n1191), .Y(PRODUCT[36]) );
  OAI21XL U1164 ( .A0(n1272), .A1(n1275), .B0(n1273), .Y(n1216) );
  AOI21XL U1165 ( .A0(n1219), .A1(n1212), .B0(n1216), .Y(n1197) );
  OAI21XL U1166 ( .A0(n5), .A1(n1198), .B0(n1197), .Y(n1200) );
  OAI21XL U1167 ( .A0(n1210), .A1(n1207), .B0(n1208), .Y(n1206) );
  INVXL U1168 ( .A(n1202), .Y(n1204) );
  AOI21XL U1169 ( .A0(n1219), .A1(n1218), .B0(n1217), .Y(n1220) );
  OAI21XL U1170 ( .A0(n5), .A1(n1221), .B0(n1220), .Y(n1224) );
  OR2XL U1171 ( .A(n1227), .B(n1233), .Y(n1237) );
  OAI21XL U1172 ( .A0(n1228), .A1(n1268), .B0(n1269), .Y(n1229) );
  AOI21XL U1173 ( .A0(n1231), .A1(n1230), .B0(n1229), .Y(n1232) );
  OAI21XL U1174 ( .A0(n1234), .A1(n1233), .B0(n1232), .Y(n1235) );
  OAI21XL U1175 ( .A0(n5), .A1(n1237), .B0(n1236), .Y(n1238) );
  XOR2XL U1176 ( .A(n1259), .B(n1258), .Y(n1340) );
endmodule


module FFT2048_DW02_mult_2_stage_J1_4 ( A, B, TC, CLK, PRODUCT );
  input [25:0] A;
  input [16:0] B;
  output [42:0] PRODUCT;
  input TC, CLK;
  wire   n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, mult_x_1_n633, mult_x_1_n618, mult_x_1_n601,
         mult_x_1_n586, mult_x_1_n585, mult_x_1_n570, mult_x_1_n569,
         mult_x_1_n554, mult_x_1_n507, mult_x_1_n494, mult_x_1_n321,
         mult_x_1_n318, mult_x_1_n317, mult_x_1_n309, mult_x_1_n305,
         mult_x_1_n304, mult_x_1_n300, mult_x_1_n299, mult_x_1_n293,
         mult_x_1_n292, mult_x_1_n287, mult_x_1_n286, mult_x_1_n282,
         mult_x_1_n281, mult_x_1_n277, mult_x_1_n276, mult_x_1_n274,
         mult_x_1_n273, mult_x_1_n263, mult_x_1_n262, mult_x_1_n227,
         mult_x_1_n226, mult_x_1_n216, mult_x_1_n215, mult_x_1_n207,
         mult_x_1_n206, mult_x_1_n195, mult_x_1_n194, mult_x_1_n184,
         mult_x_1_n183, mult_x_1_n177, mult_x_1_n176, mult_x_1_n170,
         mult_x_1_n169, mult_x_1_n161, mult_x_1_n160, mult_x_1_n152,
         mult_x_1_n151, mult_x_1_n137, mult_x_1_n136, mult_x_1_n130,
         mult_x_1_n129, mult_x_1_n121, mult_x_1_n120, mult_x_1_n110,
         mult_x_1_n109, mult_x_1_n86, mult_x_1_n85, mult_x_1_n84, mult_x_1_n58,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354;

  DFFHQXL mult_x_1_clk_r_REG18_S1 ( .D(mult_x_1_n160), .CK(CLK), .Q(n1311) );
  DFFHQX4 mult_x_1_clk_r_REG38_S1 ( .D(mult_x_1_n633), .CK(CLK), .Q(n1354) );
  DFFHQX4 mult_x_1_clk_r_REG37_S1 ( .D(mult_x_1_n618), .CK(CLK), .Q(n1353) );
  DFFHQX4 mult_x_1_clk_r_REG34_S1 ( .D(mult_x_1_n601), .CK(CLK), .Q(n1352) );
  DFFHQX4 mult_x_1_clk_r_REG33_S1 ( .D(mult_x_1_n586), .CK(CLK), .Q(n1351) );
  DFFHQX4 mult_x_1_clk_r_REG32_S1 ( .D(mult_x_1_n585), .CK(CLK), .Q(n1350) );
  DFFHQX4 mult_x_1_clk_r_REG31_S1 ( .D(mult_x_1_n570), .CK(CLK), .Q(n1349) );
  DFFHQX4 mult_x_1_clk_r_REG55_S1 ( .D(mult_x_1_n309), .CK(CLK), .Q(n1344) );
  DFFHQX4 mult_x_1_clk_r_REG49_S1 ( .D(mult_x_1_n300), .CK(CLK), .Q(n1340) );
  DFFHQX4 mult_x_1_clk_r_REG50_S1 ( .D(mult_x_1_n299), .CK(CLK), .Q(n1339) );
  DFFHQX1 mult_x_1_clk_r_REG47_S1 ( .D(mult_x_1_n293), .CK(CLK), .Q(n1338) );
  DFFHQX4 mult_x_1_clk_r_REG45_S1 ( .D(mult_x_1_n287), .CK(CLK), .Q(n1336) );
  DFFHQX4 mult_x_1_clk_r_REG46_S1 ( .D(mult_x_1_n286), .CK(CLK), .Q(n1335) );
  DFFHQX4 mult_x_1_clk_r_REG44_S1 ( .D(mult_x_1_n281), .CK(CLK), .Q(n1333) );
  DFFHQX4 mult_x_1_clk_r_REG42_S1 ( .D(mult_x_1_n276), .CK(CLK), .Q(n1331) );
  DFFHQX1 mult_x_1_clk_r_REG39_S1 ( .D(mult_x_1_n274), .CK(CLK), .Q(n1330) );
  DFFHQXL mult_x_1_clk_r_REG5_S1 ( .D(mult_x_1_n207), .CK(CLK), .Q(n1322) );
  DFFHQXL mult_x_1_clk_r_REG6_S1 ( .D(mult_x_1_n206), .CK(CLK), .Q(n1321) );
  DFFHQX4 mult_x_1_clk_r_REG52_S1 ( .D(mult_x_1_n305), .CK(CLK), .Q(n1296) );
  DFFHQX2 mult_x_1_clk_r_REG53_S1 ( .D(mult_x_1_n304), .CK(CLK), .Q(n1295) );
  DFFHQXL clk_r_REG59_S1 ( .D(n1367), .CK(CLK), .Q(PRODUCT[11]) );
  DFFHQXL mult_x_1_clk_r_REG15_S1 ( .D(mult_x_1_n170), .CK(CLK), .Q(n1314) );
  DFFHQXL clk_r_REG61_S1 ( .D(n1368), .CK(CLK), .Q(PRODUCT[10]) );
  DFFHQXL mult_x_1_clk_r_REG51_S1 ( .D(mult_x_1_n84), .CK(CLK), .Q(n1341) );
  DFFHQXL mult_x_1_clk_r_REG17_S1 ( .D(mult_x_1_n161), .CK(CLK), .Q(n1312) );
  DFFHQXL clk_r_REG62_S1 ( .D(n1369), .CK(CLK), .Q(PRODUCT[9]) );
  DFFHQXL mult_x_1_clk_r_REG14_S1 ( .D(mult_x_1_n176), .CK(CLK), .Q(n1315) );
  DFFHQXL mult_x_1_clk_r_REG13_S1 ( .D(mult_x_1_n177), .CK(CLK), .Q(n1316) );
  DFFHQXL mult_x_1_clk_r_REG3_S1 ( .D(mult_x_1_n216), .CK(CLK), .Q(n1324) );
  DFFHQXL clk_r_REG69_S1 ( .D(n1376), .CK(CLK), .Q(PRODUCT[2]) );
  DFFHQXL mult_x_1_clk_r_REG1_S1 ( .D(mult_x_1_n227), .CK(CLK), .Q(n1326) );
  DFFHQXL mult_x_1_clk_r_REG29_S1 ( .D(mult_x_1_n58), .CK(CLK), .Q(n1300) );
  DFFHQXL mult_x_1_clk_r_REG16_S1 ( .D(mult_x_1_n169), .CK(CLK), .Q(n1313) );
  DFFHQX4 mult_x_1_clk_r_REG40_S1 ( .D(mult_x_1_n273), .CK(CLK), .Q(n1329) );
  DFFHQXL mult_x_1_clk_r_REG9_S1 ( .D(mult_x_1_n195), .CK(CLK), .Q(n1320) );
  DFFHQXL clk_r_REG63_S1 ( .D(n1370), .CK(CLK), .Q(PRODUCT[8]) );
  DFFHQXL clk_r_REG64_S1 ( .D(n1371), .CK(CLK), .Q(PRODUCT[7]) );
  DFFHQXL clk_r_REG65_S1 ( .D(n1372), .CK(CLK), .Q(PRODUCT[6]) );
  DFFHQXL clk_r_REG66_S1 ( .D(n1373), .CK(CLK), .Q(PRODUCT[5]) );
  DFFHQXL clk_r_REG67_S1 ( .D(n1374), .CK(CLK), .Q(PRODUCT[4]) );
  DFFHQXL clk_r_REG68_S1 ( .D(n1375), .CK(CLK), .Q(PRODUCT[3]) );
  DFFHQXL clk_r_REG70_S1 ( .D(n1377), .CK(CLK), .Q(PRODUCT[1]) );
  DFFHQXL clk_r_REG71_S1 ( .D(n1378), .CK(CLK), .Q(PRODUCT[0]) );
  DFFHQXL mult_x_1_clk_r_REG4_S1 ( .D(mult_x_1_n215), .CK(CLK), .Q(n1323) );
  DFFHQXL mult_x_1_clk_r_REG12_S1 ( .D(mult_x_1_n183), .CK(CLK), .Q(n1317) );
  DFFHQXL mult_x_1_clk_r_REG56_S1 ( .D(mult_x_1_n86), .CK(CLK), .Q(n1343) );
  DFFHQX1 mult_x_1_clk_r_REG54_S1 ( .D(mult_x_1_n85), .CK(CLK), .Q(n1342) );
  DFFHQXL mult_x_1_clk_r_REG10_S1 ( .D(mult_x_1_n194), .CK(CLK), .Q(n1319) );
  DFFHQXL mult_x_1_clk_r_REG11_S1 ( .D(mult_x_1_n184), .CK(CLK), .Q(n1318) );
  DFFHQXL mult_x_1_clk_r_REG19_S1 ( .D(mult_x_1_n152), .CK(CLK), .Q(n1310) );
  DFFHQXL mult_x_1_clk_r_REG21_S1 ( .D(mult_x_1_n137), .CK(CLK), .Q(n1308) );
  DFFHQXL mult_x_1_clk_r_REG23_S1 ( .D(mult_x_1_n130), .CK(CLK), .Q(n1306) );
  DFFHQXL mult_x_1_clk_r_REG24_S1 ( .D(mult_x_1_n129), .CK(CLK), .Q(n1305) );
  DFFHQXL mult_x_1_clk_r_REG25_S1 ( .D(mult_x_1_n121), .CK(CLK), .Q(n1304) );
  DFFHQXL mult_x_1_clk_r_REG26_S1 ( .D(mult_x_1_n120), .CK(CLK), .Q(n1303) );
  DFFHQXL mult_x_1_clk_r_REG27_S1 ( .D(mult_x_1_n110), .CK(CLK), .Q(n1302) );
  DFFHQXL mult_x_1_clk_r_REG28_S1 ( .D(mult_x_1_n109), .CK(CLK), .Q(n1301) );
  DFFHQX2 mult_x_1_clk_r_REG60_S1 ( .D(mult_x_1_n321), .CK(CLK), .Q(n1299) );
  DFFHQX1 mult_x_1_clk_r_REG57_S1 ( .D(mult_x_1_n318), .CK(CLK), .Q(n1298) );
  DFFHQX2 mult_x_1_clk_r_REG58_S1 ( .D(mult_x_1_n317), .CK(CLK), .Q(n1297) );
  DFFHQXL mult_x_1_clk_r_REG22_S1 ( .D(mult_x_1_n136), .CK(CLK), .Q(n1307) );
  DFFHQXL mult_x_1_clk_r_REG20_S1 ( .D(mult_x_1_n151), .CK(CLK), .Q(n1309) );
  DFFHQX4 mult_x_1_clk_r_REG2_S1 ( .D(mult_x_1_n226), .CK(CLK), .Q(n1325) );
  DFFHQX4 mult_x_1_clk_r_REG48_S1 ( .D(mult_x_1_n292), .CK(CLK), .Q(n1337) );
  DFFHQXL mult_x_1_clk_r_REG7_S1 ( .D(mult_x_1_n507), .CK(CLK), .Q(n1346) );
  DFFHQXL mult_x_1_clk_r_REG8_S1 ( .D(mult_x_1_n494), .CK(CLK), .Q(n1345) );
  DFFHQX1 mult_x_1_clk_r_REG43_S1 ( .D(mult_x_1_n282), .CK(CLK), .Q(n1334) );
  DFFHQX2 mult_x_1_clk_r_REG30_S1 ( .D(mult_x_1_n569), .CK(CLK), .Q(n1348) );
  DFFHQX2 mult_x_1_clk_r_REG0_S1 ( .D(mult_x_1_n554), .CK(CLK), .Q(n1347) );
  DFFHQX1 mult_x_1_clk_r_REG41_S1 ( .D(mult_x_1_n277), .CK(CLK), .Q(n1332) );
  DFFHQX1 mult_x_1_clk_r_REG35_S1 ( .D(mult_x_1_n263), .CK(CLK), .Q(n1328) );
  DFFHQX1 mult_x_1_clk_r_REG36_S1 ( .D(mult_x_1_n262), .CK(CLK), .Q(n1327) );
  ADDFX2 U1 ( .A(n805), .B(n804), .CI(n803), .CO(n796), .S(n829) );
  ADDFHX1 U2 ( .A(n745), .B(n744), .CI(n743), .CO(n736), .S(n771) );
  ADDFHX2 U3 ( .A(n429), .B(n428), .CI(n427), .CO(n1078), .S(n440) );
  ADDFHX1 U4 ( .A(n1112), .B(n1111), .CI(n1110), .CO(n1117), .S(n1119) );
  CMPR32X1 U5 ( .A(n1094), .B(n1093), .C(n1092), .CO(n1115), .S(n1110) );
  ADDFHX1 U6 ( .A(n511), .B(n510), .CI(n509), .CO(n514), .S(n1101) );
  ADDFX2 U7 ( .A(n394), .B(n393), .CI(n392), .CO(n1079), .S(n428) );
  ADDFHX2 U8 ( .A(n748), .B(n747), .CI(n746), .CO(n734), .S(n774) );
  ADDFX2 U9 ( .A(n559), .B(n558), .CI(n557), .CO(n574), .S(n624) );
  CMPR32X1 U10 ( .A(n282), .B(n281), .C(n280), .CO(n302), .S(n318) );
  ADDFX2 U11 ( .A(n592), .B(n591), .CI(n590), .CO(n1100), .S(n1093) );
  ADDFHX1 U12 ( .A(n663), .B(n662), .CI(n661), .CO(n666), .S(n700) );
  ADDFHX1 U13 ( .A(n1050), .B(n1049), .CI(n1048), .CO(n1051), .S(n918) );
  ADDFHX1 U14 ( .A(n605), .B(n604), .CI(n603), .CO(n556), .S(n621) );
  ADDFHX1 U15 ( .A(n577), .B(n576), .CI(n575), .CO(n1109), .S(n555) );
  ADDFHX1 U16 ( .A(n502), .B(n501), .CI(n500), .CO(n511), .S(n1099) );
  ADDFHX1 U17 ( .A(n1085), .B(n1084), .CI(n1083), .CO(n1097), .S(n1108) );
  ADDFHX2 U18 ( .A(n448), .B(n447), .CI(n446), .CO(n426), .S(n465) );
  ADDFHX2 U19 ( .A(n491), .B(n490), .CI(n489), .CO(n466), .S(n507) );
  OAI22X1 U20 ( .A0(n82), .A1(n497), .B0(n7), .B1(n455), .Y(n502) );
  ADDFHX1 U21 ( .A(n350), .B(n349), .CI(n348), .CO(n337), .S(n407) );
  ADDFHX1 U22 ( .A(n724), .B(n723), .CI(n722), .CO(n735), .S(n768) );
  ADDFHX1 U23 ( .A(n755), .B(n754), .CI(n753), .CO(n769), .S(n794) );
  ADDFHX1 U24 ( .A(n616), .B(n615), .CI(n614), .CO(n625), .S(n662) );
  ADDFHX1 U25 ( .A(n677), .B(n676), .CI(n675), .CO(n663), .S(n708) );
  ADDFHX1 U26 ( .A(n1032), .B(n1031), .CI(n1030), .CO(n1022), .S(n1033) );
  ADDFX2 U27 ( .A(n314), .B(n313), .CI(n312), .CO(n306), .S(n349) );
  ADDFX2 U28 ( .A(n1038), .B(n1037), .CI(n1036), .CO(n1039), .S(n1019) );
  XNOR2X1 U29 ( .A(n867), .B(A[9]), .Y(n547) );
  ADDFHX1 U30 ( .A(n687), .B(n686), .CI(n685), .CO(n699), .S(n722) );
  BUFX8 U31 ( .A(n681), .Y(n1199) );
  CLKBUFX8 U32 ( .A(n713), .Y(n1200) );
  BUFX3 U33 ( .A(B[16]), .Y(n1194) );
  NAND2X2 U34 ( .A(n157), .B(n713), .Y(n681) );
  XOR2X1 U35 ( .A(n867), .B(n118), .Y(n117) );
  ADDFHX1 U36 ( .A(n932), .B(n931), .CI(n930), .CO(n1014), .S(n933) );
  BUFX4 U37 ( .A(n906), .Y(n912) );
  BUFX4 U38 ( .A(B[13]), .Y(n1138) );
  BUFX3 U39 ( .A(n550), .Y(n986) );
  BUFX8 U40 ( .A(n454), .Y(n7) );
  BUFX3 U41 ( .A(n650), .Y(n9) );
  CLKBUFX8 U42 ( .A(B[9]), .Y(n331) );
  INVX4 U43 ( .A(n929), .Y(n8) );
  BUFX3 U44 ( .A(n869), .Y(n1137) );
  BUFX3 U45 ( .A(n599), .Y(n6) );
  BUFX4 U46 ( .A(n1000), .Y(n924) );
  CLKINVX3 U47 ( .A(B[11]), .Y(n850) );
  NAND2X2 U48 ( .A(n83), .B(n454), .Y(n869) );
  NAND2X1 U49 ( .A(n599), .B(n64), .Y(n1000) );
  NAND2X1 U50 ( .A(n13), .B(n950), .Y(n983) );
  CLKBUFX3 U51 ( .A(B[1]), .Y(n678) );
  INVX2 U52 ( .A(B[7]), .Y(n920) );
  OAI21XL U53 ( .A0(n635), .A1(n436), .B0(n435), .Y(n439) );
  XOR2X1 U54 ( .A(n130), .B(n137), .Y(PRODUCT[19]) );
  XOR2X1 U55 ( .A(n638), .B(n637), .Y(PRODUCT[20]) );
  NOR2XL U56 ( .A(n434), .B(n37), .Y(n435) );
  NAND2XL U57 ( .A(n477), .B(n38), .Y(n35) );
  NAND2X1 U58 ( .A(n532), .B(n142), .Y(n34) );
  NOR2X1 U59 ( .A(n1352), .B(n1351), .Y(n523) );
  OAI22X1 U60 ( .A0(n681), .A1(n396), .B0(n1200), .B1(n335), .Y(n380) );
  AOI21XL U61 ( .A0(n477), .A1(n519), .B0(n476), .Y(n478) );
  AND2X1 U62 ( .A(n636), .B(n1330), .Y(n637) );
  OAI21XL U63 ( .A0(n1290), .A1(n1219), .B0(n1218), .Y(n1258) );
  CLKINVX3 U64 ( .A(n55), .Y(n1293) );
  XNOR2X1 U65 ( .A(n296), .B(n295), .Y(PRODUCT[31]) );
  XNOR2XL U66 ( .A(n867), .B(A[0]), .Y(n868) );
  XNOR2XL U67 ( .A(n922), .B(A[1]), .Y(n999) );
  XNOR2XL U68 ( .A(n922), .B(A[4]), .Y(n890) );
  XNOR2XL U69 ( .A(n1138), .B(A[16]), .Y(n275) );
  XNOR2XL U70 ( .A(n1184), .B(A[14]), .Y(n272) );
  XNOR2XL U71 ( .A(n867), .B(A[19]), .Y(n238) );
  XNOR2XL U72 ( .A(n766), .B(n95), .Y(n721) );
  XNOR2XL U73 ( .A(n766), .B(n89), .Y(n445) );
  XNOR2XL U74 ( .A(n867), .B(A[11]), .Y(n560) );
  BUFX3 U75 ( .A(n869), .Y(n82) );
  XNOR2XL U76 ( .A(n867), .B(A[20]), .Y(n231) );
  XNOR2XL U77 ( .A(n766), .B(n99), .Y(n1174) );
  XNOR2XL U78 ( .A(B[2]), .B(B[1]), .Y(n950) );
  XNOR2XL U79 ( .A(n1184), .B(A[12]), .Y(n335) );
  XNOR2XL U80 ( .A(n766), .B(n88), .Y(n583) );
  XNOR2XL U81 ( .A(n922), .B(A[13]), .Y(n600) );
  ADDFX2 U82 ( .A(n732), .B(n731), .CI(n730), .CO(n748), .S(n775) );
  ADDFX2 U83 ( .A(n589), .B(n588), .CI(n587), .CO(n1094), .S(n573) );
  OAI2BB1X1 U84 ( .A0N(n30), .A1N(n767), .B0(n29), .Y(n744) );
  XNOR2XL U85 ( .A(n1236), .B(n1235), .Y(n1371) );
  XOR2XL U86 ( .A(n1073), .B(n1072), .Y(n1369) );
  XNOR2X1 U87 ( .A(n56), .B(n370), .Y(PRODUCT[28]) );
  INVX1 U88 ( .A(n477), .Y(n39) );
  NAND2XL U89 ( .A(n61), .B(n1065), .Y(n1062) );
  XOR2X1 U90 ( .A(n1068), .B(n1067), .Y(n1368) );
  NAND2XL U91 ( .A(n19), .B(n385), .Y(n18) );
  NAND2X1 U92 ( .A(n1041), .B(n1042), .Y(n1059) );
  NAND2X1 U93 ( .A(n1040), .B(n1039), .Y(n1065) );
  ADDFHX2 U94 ( .A(n1115), .B(n1114), .CI(n1113), .CO(n1105), .S(n1116) );
  INVX1 U95 ( .A(n22), .Y(n20) );
  NOR2X1 U96 ( .A(n1196), .B(n196), .Y(n224) );
  NOR2X1 U97 ( .A(n1196), .B(n648), .Y(n673) );
  NOR2X1 U98 ( .A(n1196), .B(n154), .Y(n204) );
  NOR2X1 U99 ( .A(n1196), .B(n153), .Y(n172) );
  NOR2X1 U100 ( .A(n1196), .B(n159), .Y(n180) );
  NOR2X1 U101 ( .A(n1196), .B(n175), .Y(n1142) );
  NOR2X1 U102 ( .A(n1196), .B(n218), .Y(n241) );
  NAND2X1 U103 ( .A(n973), .B(n972), .Y(n1242) );
  XNOR2X1 U104 ( .A(n1263), .B(n1262), .Y(PRODUCT[39]) );
  NAND2XL U105 ( .A(n54), .B(n255), .Y(n259) );
  OAI22X1 U106 ( .A0(n992), .A1(n562), .B0(n990), .B1(n498), .Y(n591) );
  OAI22XL U107 ( .A0(n942), .A1(n820), .B0(n765), .B1(n1128), .Y(n818) );
  NAND2XL U108 ( .A(n535), .B(n534), .Y(n536) );
  NAND2X1 U109 ( .A(n740), .B(n1334), .Y(n741) );
  NAND2X1 U110 ( .A(n126), .B(n1332), .Y(n137) );
  NAND2X1 U111 ( .A(n257), .B(n1316), .Y(n258) );
  NAND2X1 U112 ( .A(n480), .B(n1326), .Y(n481) );
  NAND2X1 U113 ( .A(n437), .B(n1324), .Y(n438) );
  NAND2X1 U114 ( .A(n1347), .B(n1348), .Y(n518) );
  INVX1 U115 ( .A(n1335), .Y(n138) );
  INVX1 U116 ( .A(A[5]), .Y(n28) );
  ADDFHX1 U117 ( .A(n1076), .B(n1075), .CI(n1074), .CO(n358), .S(mult_x_1_n494) );
  NAND2X1 U118 ( .A(n883), .B(n882), .Y(n884) );
  OAI2BB1X1 U119 ( .A0N(n386), .A1N(n22), .B0(n18), .Y(n411) );
  NAND2XL U120 ( .A(n701), .B(n702), .Y(n77) );
  XOR2X1 U121 ( .A(n702), .B(n700), .Y(n112) );
  XNOR2X1 U122 ( .A(n1211), .B(n1210), .Y(n1370) );
  NOR2X1 U123 ( .A(n1040), .B(n1039), .Y(n1064) );
  ADDFHX1 U124 ( .A(n1118), .B(n1117), .CI(n1116), .CO(mult_x_1_n585), .S(
        mult_x_1_n586) );
  ADDFHX1 U125 ( .A(n1106), .B(n1105), .CI(n1104), .CO(mult_x_1_n569), .S(
        mult_x_1_n570) );
  NAND2BX1 U126 ( .AN(n386), .B(n20), .Y(n19) );
  ADDFHX1 U127 ( .A(n628), .B(n627), .CI(n626), .CO(n1120), .S(n1122) );
  OR2X2 U128 ( .A(n768), .B(n769), .Y(n30) );
  INVX1 U129 ( .A(n407), .Y(n17) );
  ADDFHX1 U130 ( .A(n1103), .B(n1102), .CI(n1101), .CO(n1081), .S(n1104) );
  ADDFHX1 U131 ( .A(n1100), .B(n1099), .CI(n1098), .CO(n1103), .S(n1113) );
  NAND2X1 U132 ( .A(n25), .B(n23), .Y(n22) );
  NAND2BXL U133 ( .AN(n466), .B(n44), .Y(n43) );
  NAND2X1 U134 ( .A(n1017), .B(n1016), .Y(n1208) );
  INVXL U135 ( .A(n642), .Y(n73) );
  ADDHXL U136 ( .A(n818), .B(n817), .CO(n814), .S(n865) );
  NOR2X1 U137 ( .A(n975), .B(n974), .Y(n1232) );
  NOR2X1 U138 ( .A(n973), .B(n972), .Y(n1241) );
  OAI22XL U139 ( .A0(n912), .A1(n274), .B0(n904), .B1(n266), .Y(n308) );
  NOR2X1 U140 ( .A(n1196), .B(n1158), .Y(n1171) );
  NOR2X1 U141 ( .A(n1196), .B(n1134), .Y(n1156) );
  OAI22X1 U142 ( .A0(n1199), .A1(n1185), .B0(n1200), .B1(n1197), .Y(n1203) );
  OAI2BB1XL U143 ( .A0N(n1200), .A1N(n1199), .B0(n1198), .Y(n1201) );
  NOR2BX1 U144 ( .AN(A[0]), .B(n1200), .Y(n786) );
  XNOR2XL U145 ( .A(n1138), .B(A[23]), .Y(n1139) );
  XNOR2X1 U146 ( .A(n151), .B(n150), .Y(PRODUCT[35]) );
  XNOR2X1 U147 ( .A(n192), .B(n191), .Y(PRODUCT[34]) );
  XNOR2X1 U148 ( .A(n1240), .B(n1239), .Y(PRODUCT[38]) );
  XNOR2X1 U149 ( .A(n1230), .B(n1229), .Y(PRODUCT[37]) );
  CLKINVX3 U150 ( .A(n714), .Y(n1168) );
  OAI2BB1X1 U151 ( .A0N(n1128), .A1N(n942), .B0(n341), .Y(n385) );
  XOR2X1 U152 ( .A(n59), .B(n536), .Y(PRODUCT[23]) );
  OR2XL U153 ( .A(n1282), .B(n1289), .Y(n1283) );
  NOR2X1 U154 ( .A(n1282), .B(n1219), .Y(n1252) );
  XNOR2X1 U155 ( .A(n802), .B(n801), .Y(PRODUCT[16]) );
  INVX1 U156 ( .A(n523), .Y(n535) );
  NAND2X1 U157 ( .A(n538), .B(n1328), .Y(n539) );
  AND2X1 U158 ( .A(n216), .B(n1314), .Y(n69) );
  NOR2X1 U159 ( .A(n359), .B(n1319), .Y(n253) );
  INVX1 U160 ( .A(A[0]), .Y(n104) );
  INVX1 U161 ( .A(n1311), .Y(n1212) );
  NAND2XL U162 ( .A(n474), .B(n473), .Y(mult_x_1_n216) );
  OAI21XL U163 ( .A0(n15), .A1(n17), .B0(n14), .Y(n1074) );
  ADDFHX2 U164 ( .A(n1079), .B(n1078), .CI(n1077), .CO(mult_x_1_n507), .S(n431) );
  NAND2X1 U165 ( .A(n797), .B(n796), .Y(mult_x_1_n287) );
  INVXL U166 ( .A(n1057), .Y(n1068) );
  INVXL U167 ( .A(n1148), .Y(mult_x_1_n318) );
  XOR2X1 U168 ( .A(n112), .B(n701), .Y(n705) );
  NAND2XL U169 ( .A(n132), .B(n774), .Y(n133) );
  XOR2X1 U170 ( .A(n134), .B(n772), .Y(n797) );
  INVXL U171 ( .A(n1051), .Y(n123) );
  ADDFHX1 U172 ( .A(n862), .B(n861), .CI(n860), .CO(n857), .S(n883) );
  NAND2XL U173 ( .A(n630), .B(n629), .Y(mult_x_1_n263) );
  XOR2X1 U174 ( .A(n386), .B(n21), .Y(n422) );
  NAND2X1 U175 ( .A(n11), .B(n10), .Y(n706) );
  XOR2X1 U176 ( .A(n767), .B(n31), .Y(n772) );
  OAI21XL U177 ( .A0(n734), .A1(n735), .B0(n733), .Y(n11) );
  NAND2X1 U178 ( .A(n734), .B(n735), .Y(n10) );
  NAND2X1 U179 ( .A(n768), .B(n769), .Y(n29) );
  OAI2BB1XL U180 ( .A0N(n80), .A1N(n506), .B0(n79), .Y(n1082) );
  NAND2BXL U181 ( .AN(n826), .B(n115), .Y(n114) );
  INVXL U182 ( .A(n825), .Y(n85) );
  NAND2BXL U183 ( .AN(n698), .B(n108), .Y(n107) );
  ADDFHX2 U184 ( .A(n338), .B(n337), .CI(n336), .CO(n354), .S(n1075) );
  OR2XL U185 ( .A(n1205), .B(n1204), .Y(n1207) );
  INVXL U186 ( .A(n699), .Y(n108) );
  ADDFHX2 U187 ( .A(n622), .B(n621), .CI(n620), .CO(n1124), .S(n665) );
  NAND2XL U188 ( .A(n826), .B(n827), .Y(n113) );
  INVXL U189 ( .A(n827), .Y(n115) );
  ADDFHX1 U190 ( .A(n865), .B(n864), .CI(n863), .CO(n854), .S(n1047) );
  OAI21XL U191 ( .A0(n66), .A1(n67), .B0(n65), .Y(n1018) );
  NAND2BX1 U192 ( .AN(n382), .B(n26), .Y(n25) );
  INVXL U193 ( .A(n465), .Y(n44) );
  NAND2XL U194 ( .A(n466), .B(n465), .Y(n42) );
  ADDFHX1 U195 ( .A(n308), .B(n307), .CI(n306), .CO(n304), .S(n338) );
  XNOR3X2 U196 ( .A(n67), .B(n1011), .C(n1010), .Y(n1017) );
  ADDFHX1 U197 ( .A(n761), .B(n760), .CI(n759), .CO(n753), .S(n807) );
  NAND2BX1 U198 ( .AN(n339), .B(n24), .Y(n23) );
  INVXL U199 ( .A(n1011), .Y(n66) );
  OAI22X1 U200 ( .A0(n812), .A1(n543), .B0(n819), .B1(n583), .Y(n575) );
  OR2X2 U201 ( .A(n962), .B(n961), .Y(n960) );
  OAI21XL U202 ( .A0(n1293), .A1(n190), .B0(n189), .Y(n192) );
  AND2XL U203 ( .A(n1279), .B(n1278), .Y(n1377) );
  NAND3X2 U204 ( .A(n145), .B(n36), .C(n35), .Y(n55) );
  OR2XL U205 ( .A(n1277), .B(n1276), .Y(n1279) );
  XOR2X1 U206 ( .A(n521), .B(n520), .Y(PRODUCT[25]) );
  INVXL U207 ( .A(B[4]), .Y(n111) );
  XOR2X1 U208 ( .A(n70), .B(n739), .Y(PRODUCT[17]) );
  NAND2X1 U209 ( .A(B[1]), .B(n953), .Y(n764) );
  NOR2XL U210 ( .A(n129), .B(n1331), .Y(n128) );
  AND2X2 U211 ( .A(n519), .B(n518), .Y(n520) );
  NOR2X1 U212 ( .A(n631), .B(n1327), .Y(n522) );
  INVX1 U213 ( .A(B[0]), .Y(n953) );
  AND2X2 U214 ( .A(n369), .B(n1322), .Y(n370) );
  INVXL U215 ( .A(A[2]), .Y(n97) );
  INVXL U216 ( .A(A[14]), .Y(n98) );
  INVXL U217 ( .A(A[19]), .Y(n96) );
  INVXL U218 ( .A(A[12]), .Y(n89) );
  INVXL U219 ( .A(A[11]), .Y(n91) );
  INVXL U220 ( .A(A[10]), .Y(n90) );
  INVXL U221 ( .A(A[25]), .Y(n99) );
  INVXL U222 ( .A(A[6]), .Y(n93) );
  INVXL U223 ( .A(A[8]), .Y(n92) );
  INVXL U224 ( .A(A[9]), .Y(n88) );
  INVXL U225 ( .A(A[3]), .Y(n95) );
  INVXL U226 ( .A(A[4]), .Y(n94) );
  OAI21XL U227 ( .A0(n1329), .A1(n1332), .B0(n1330), .Y(n47) );
  INVXL U228 ( .A(n1331), .Y(n126) );
  INVXL U229 ( .A(n1332), .Y(n125) );
  NAND2X1 U230 ( .A(n1052), .B(n1051), .Y(n1055) );
  OAI21XL U231 ( .A0(n897), .A1(n898), .B0(n896), .Y(n120) );
  NAND2X1 U232 ( .A(n122), .B(n1056), .Y(n1053) );
  XNOR2X1 U233 ( .A(n381), .B(n380), .Y(n403) );
  AOI2BB1X1 U234 ( .A0N(n368), .A1N(n635), .B0(n57), .Y(n56) );
  NAND2X2 U235 ( .A(n34), .B(n32), .Y(n477) );
  XNOR2X1 U236 ( .A(n907), .B(n102), .Y(n1031) );
  NOR2X2 U237 ( .A(n7), .B(n104), .Y(n103) );
  NOR2X1 U238 ( .A(n1042), .B(n1041), .Y(n1058) );
  AOI21X1 U239 ( .A0(n1057), .A1(n1044), .B0(n1043), .Y(n1063) );
  XOR2X2 U240 ( .A(n466), .B(n465), .Y(n45) );
  OAI2BB1X1 U241 ( .A0N(n107), .A1N(n697), .B0(n106), .Y(n702) );
  XNOR2X1 U242 ( .A(B[4]), .B(B[3]), .Y(n650) );
  OAI22X1 U243 ( .A0(n986), .A1(n651), .B0(n9), .B1(n640), .Y(n653) );
  XNOR2X1 U244 ( .A(n12), .B(n733), .Y(n743) );
  XNOR2X1 U245 ( .A(n734), .B(n735), .Y(n12) );
  XOR2X1 U246 ( .A(B[3]), .B(B[2]), .Y(n13) );
  INVX1 U247 ( .A(n1052), .Y(n121) );
  NAND2X1 U248 ( .A(n431), .B(n430), .Y(mult_x_1_n207) );
  OAI21XL U249 ( .A0(n408), .A1(n407), .B0(n406), .Y(n14) );
  INVX1 U250 ( .A(n408), .Y(n15) );
  XOR2X2 U251 ( .A(n16), .B(n408), .Y(n1077) );
  XNOR2X2 U252 ( .A(n406), .B(n17), .Y(n16) );
  XOR2X1 U253 ( .A(n22), .B(n385), .Y(n21) );
  INVX1 U254 ( .A(n7), .Y(n24) );
  INVX1 U255 ( .A(n1137), .Y(n26) );
  OAI22X1 U256 ( .A0(n82), .A1(n757), .B0(n7), .B1(n27), .Y(n779) );
  OAI22X1 U257 ( .A0(n82), .A1(n27), .B0(n689), .B1(n7), .Y(n731) );
  XOR2X1 U258 ( .A(n867), .B(n28), .Y(n27) );
  XOR2X1 U259 ( .A(n768), .B(n769), .Y(n31) );
  NAND2BX2 U260 ( .AN(n1337), .B(n1344), .Y(n52) );
  AOI21X1 U261 ( .A0(n537), .A1(n522), .B0(n60), .Y(n59) );
  NOR2BX1 U262 ( .AN(n528), .B(n33), .Y(n32) );
  NOR2X1 U263 ( .A(n534), .B(n527), .Y(n33) );
  NAND2X1 U264 ( .A(n1351), .B(n1352), .Y(n534) );
  OAI21X2 U265 ( .A0(n1327), .A1(n632), .B0(n1328), .Y(n532) );
  NAND2X2 U266 ( .A(n1354), .B(n1353), .Y(n632) );
  NAND2X1 U267 ( .A(n40), .B(n537), .Y(n36) );
  AND2X4 U268 ( .A(n477), .B(n363), .Y(n37) );
  INVX1 U269 ( .A(n41), .Y(n38) );
  NAND2X1 U270 ( .A(n144), .B(n363), .Y(n41) );
  NOR2X2 U271 ( .A(n1321), .B(n1323), .Y(n144) );
  NOR2X1 U272 ( .A(n364), .B(n41), .Y(n40) );
  NOR2X2 U273 ( .A(n1325), .B(n475), .Y(n363) );
  NAND2X1 U274 ( .A(n142), .B(n522), .Y(n364) );
  OAI21X4 U275 ( .A0(n141), .A1(n48), .B0(n46), .Y(n537) );
  NOR2X4 U276 ( .A(n51), .B(n50), .Y(n141) );
  OAI2BB1XL U277 ( .A0N(n43), .A1N(n464), .B0(n42), .Y(n485) );
  XOR2X2 U278 ( .A(n464), .B(n45), .Y(n513) );
  INVX4 U279 ( .A(n537), .Y(n635) );
  AOI21X2 U280 ( .A0(n140), .A1(n49), .B0(n47), .Y(n46) );
  OAI21X2 U281 ( .A0(n1333), .A1(n1336), .B0(n1334), .Y(n140) );
  NAND2X1 U282 ( .A(n139), .B(n49), .Y(n48) );
  NOR2X1 U283 ( .A(n1329), .B(n1331), .Y(n49) );
  NOR2X1 U284 ( .A(n1333), .B(n1335), .Y(n139) );
  NOR2X2 U285 ( .A(n798), .B(n1337), .Y(n50) );
  OAI21X4 U286 ( .A0(n52), .A1(n799), .B0(n1338), .Y(n51) );
  XOR2X1 U287 ( .A(n53), .B(n1342), .Y(PRODUCT[13]) );
  AOI21X1 U288 ( .A0(n1299), .A1(n1297), .B0(n1298), .Y(n53) );
  NAND2BX1 U289 ( .AN(n256), .B(n55), .Y(n54) );
  OR2X2 U290 ( .A(n58), .B(n366), .Y(n57) );
  NOR2BX1 U291 ( .AN(n367), .B(n39), .Y(n58) );
  NOR2X2 U292 ( .A(n1350), .B(n1349), .Y(n527) );
  INVXL U293 ( .A(n533), .Y(n60) );
  NAND2BX1 U294 ( .AN(n1064), .B(n1057), .Y(n61) );
  NAND2X1 U295 ( .A(n63), .B(n62), .Y(n1057) );
  NAND3BX1 U296 ( .AN(n1069), .B(n1209), .C(n135), .Y(n62) );
  AOI21X1 U297 ( .A0(n1070), .A1(n135), .B0(n1020), .Y(n63) );
  XOR2X1 U298 ( .A(B[6]), .B(B[7]), .Y(n64) );
  OAI21XL U299 ( .A0(n1011), .A1(n1012), .B0(n1010), .Y(n65) );
  INVX1 U300 ( .A(n1012), .Y(n67) );
  XNOR2XL U301 ( .A(n678), .B(A[14]), .Y(n751) );
  NAND2XL U302 ( .A(n1228), .B(n1306), .Y(n1229) );
  XNOR2X1 U303 ( .A(B[6]), .B(B[5]), .Y(n599) );
  BUFX4 U304 ( .A(B[16]), .Y(n668) );
  NAND2XL U305 ( .A(n1212), .B(n1214), .Y(n1217) );
  NAND2XL U306 ( .A(n1225), .B(n1308), .Y(n1222) );
  XNOR2XL U307 ( .A(n678), .B(A[25]), .Y(n378) );
  XNOR2XL U308 ( .A(n678), .B(A[24]), .Y(n390) );
  INVX1 U309 ( .A(A[1]), .Y(n118) );
  XNOR2XL U310 ( .A(n678), .B(A[11]), .Y(n848) );
  XNOR2XL U311 ( .A(n331), .B(A[1]), .Y(n910) );
  XNOR2XL U312 ( .A(n8), .B(A[5]), .Y(n913) );
  XNOR2XL U313 ( .A(n8), .B(A[24]), .Y(n271) );
  XNOR2XL U314 ( .A(n8), .B(A[25]), .Y(n220) );
  XNOR2XL U315 ( .A(n1168), .B(A[16]), .Y(n229) );
  XNOR2XL U316 ( .A(n1168), .B(A[19]), .Y(n162) );
  XNOR2XL U317 ( .A(n1168), .B(A[17]), .Y(n197) );
  XNOR2XL U318 ( .A(n331), .B(A[23]), .Y(n195) );
  XNOR2XL U319 ( .A(n331), .B(A[24]), .Y(n165) );
  AOI21XL U320 ( .A0(n1258), .A1(n1251), .B0(n1255), .Y(n1237) );
  NAND2X1 U321 ( .A(n127), .B(n124), .Y(n638) );
  XNOR2XL U322 ( .A(n1168), .B(A[21]), .Y(n1140) );
  XNOR2XL U323 ( .A(n1168), .B(A[20]), .Y(n174) );
  AND2X1 U324 ( .A(n750), .B(n116), .Y(n755) );
  NAND2X1 U325 ( .A(n219), .B(n650), .Y(n550) );
  XNOR2X1 U326 ( .A(B[5]), .B(n111), .Y(n219) );
  XNOR2XL U327 ( .A(n922), .B(A[14]), .Y(n541) );
  XNOR2XL U328 ( .A(n1184), .B(A[5]), .Y(n601) );
  XNOR2XL U329 ( .A(n1184), .B(A[4]), .Y(n612) );
  XNOR2XL U330 ( .A(n8), .B(A[14]), .Y(n640) );
  BUFX3 U331 ( .A(n983), .Y(n992) );
  BUFX3 U332 ( .A(n950), .Y(n990) );
  XNOR2XL U333 ( .A(n1184), .B(A[25]), .Y(n1197) );
  XNOR2XL U334 ( .A(n1168), .B(A[24]), .Y(n1185) );
  OAI2BB1XL U335 ( .A0N(n1177), .A1N(n1176), .B0(n1175), .Y(n1186) );
  NOR2XL U336 ( .A(n1196), .B(n1173), .Y(n1187) );
  INVXL U337 ( .A(n1174), .Y(n1175) );
  XNOR2XL U338 ( .A(n1168), .B(A[23]), .Y(n1169) );
  OAI22XL U339 ( .A0(n942), .A1(n567), .B0(n495), .B1(n1128), .Y(n596) );
  OAI22XL U340 ( .A0(n924), .A1(n578), .B0(n6), .B1(n486), .Y(n1088) );
  OAI22X1 U341 ( .A0(n1199), .A1(n580), .B0(n1200), .B1(n487), .Y(n1087) );
  INVXL U342 ( .A(n1312), .Y(n1215) );
  NOR2XL U343 ( .A(n1307), .B(n1305), .Y(n1251) );
  AOI21XL U344 ( .A0(n188), .A1(n1212), .B0(n1215), .Y(n148) );
  INVXL U345 ( .A(n1309), .Y(n1214) );
  NAND2XL U346 ( .A(n253), .B(n294), .Y(n256) );
  INVXL U347 ( .A(n1318), .Y(n254) );
  INVXL U348 ( .A(n1315), .Y(n257) );
  INVXL U349 ( .A(n1313), .Y(n216) );
  INVXL U350 ( .A(n1317), .Y(n294) );
  INVXL U351 ( .A(n475), .Y(n519) );
  XNOR2XL U352 ( .A(n678), .B(A[12]), .Y(n820) );
  XNOR2XL U353 ( .A(n981), .B(A[7]), .Y(n989) );
  ADDFX2 U354 ( .A(n717), .B(n716), .CI(n715), .CO(n724), .S(n754) );
  OAI22X1 U355 ( .A0(n942), .A1(n711), .B0(n679), .B1(n1128), .Y(n716) );
  NOR2BXL U356 ( .AN(A[0]), .B(n234), .Y(n717) );
  OAI22X1 U357 ( .A0(n681), .A1(n719), .B0(n1200), .B1(n680), .Y(n715) );
  XNOR2XL U358 ( .A(n331), .B(A[7]), .Y(n718) );
  XNOR2XL U359 ( .A(n678), .B(A[15]), .Y(n711) );
  XNOR2XL U360 ( .A(n331), .B(A[6]), .Y(n756) );
  XNOR2XL U361 ( .A(n331), .B(A[5]), .Y(n787) );
  XNOR2XL U362 ( .A(n8), .B(A[9]), .Y(n789) );
  XNOR2XL U363 ( .A(n981), .B(A[22]), .Y(n413) );
  XNOR2XL U364 ( .A(n8), .B(A[20]), .Y(n414) );
  XNOR2XL U365 ( .A(n981), .B(A[21]), .Y(n456) );
  XNOR2XL U366 ( .A(n8), .B(A[19]), .Y(n457) );
  XNOR2XL U367 ( .A(n981), .B(A[19]), .Y(n562) );
  XNOR2XL U368 ( .A(n8), .B(A[17]), .Y(n564) );
  XNOR2XL U369 ( .A(n678), .B(A[18]), .Y(n609) );
  XNOR2XL U370 ( .A(n678), .B(A[19]), .Y(n545) );
  XNOR2XL U371 ( .A(n981), .B(A[18]), .Y(n563) );
  XNOR2XL U372 ( .A(n8), .B(A[16]), .Y(n565) );
  XNOR2XL U373 ( .A(n1194), .B(A[14]), .Y(n218) );
  XNOR2XL U374 ( .A(n1168), .B(A[15]), .Y(n237) );
  XNOR2XL U375 ( .A(n981), .B(A[24]), .Y(n340) );
  INVXL U376 ( .A(n378), .Y(n341) );
  XNOR2XL U377 ( .A(n981), .B(A[23]), .Y(n383) );
  XNOR2XL U378 ( .A(n678), .B(A[6]), .Y(n921) );
  XNOR2XL U379 ( .A(n8), .B(A[2]), .Y(n925) );
  XNOR2XL U380 ( .A(n981), .B(A[5]), .Y(n982) );
  XNOR2X1 U381 ( .A(n8), .B(A[3]), .Y(n985) );
  XNOR2XL U382 ( .A(n678), .B(A[7]), .Y(n997) );
  NAND2XL U383 ( .A(n1281), .B(n1286), .Y(n1289) );
  NAND2XL U384 ( .A(n1252), .B(n1251), .Y(n1238) );
  INVXL U385 ( .A(n1303), .Y(n1254) );
  INVXL U386 ( .A(n1287), .Y(n1218) );
  INVXL U387 ( .A(n1280), .Y(n1257) );
  XNOR2XL U388 ( .A(n668), .B(A[11]), .Y(n310) );
  XNOR2XL U389 ( .A(B[9]), .B(A[17]), .Y(n387) );
  XNOR2XL U390 ( .A(n668), .B(A[9]), .Y(n379) );
  XNOR2XL U391 ( .A(n668), .B(A[10]), .Y(n372) );
  XNOR2X1 U392 ( .A(n766), .B(n87), .Y(n399) );
  INVXL U393 ( .A(A[13]), .Y(n87) );
  XNOR2XL U394 ( .A(n8), .B(A[21]), .Y(n384) );
  XNOR2XL U395 ( .A(n981), .B(A[10]), .Y(n823) );
  XNOR2XL U396 ( .A(n8), .B(A[8]), .Y(n824) );
  XNOR2XL U397 ( .A(n981), .B(A[9]), .Y(n870) );
  XNOR2XL U398 ( .A(n981), .B(A[8]), .Y(n892) );
  XNOR2XL U399 ( .A(n331), .B(A[2]), .Y(n889) );
  XNOR2X1 U400 ( .A(n8), .B(A[7]), .Y(n871) );
  XNOR2XL U401 ( .A(n331), .B(A[3]), .Y(n872) );
  OAI22XL U402 ( .A0(n764), .A1(n888), .B0(n848), .B1(n1128), .Y(n874) );
  NAND2BXL U403 ( .AN(A[0]), .B(n867), .Y(n849) );
  OAI22XL U404 ( .A0(n942), .A1(n902), .B0(n888), .B1(n1128), .Y(n908) );
  INVXL U405 ( .A(n908), .Y(n105) );
  ADDFX2 U406 ( .A(n980), .B(n979), .CI(n978), .CO(n1030), .S(n1038) );
  OAI22X1 U407 ( .A0(n912), .A1(n911), .B0(n995), .B1(n910), .Y(n979) );
  OAI22X1 U408 ( .A0(n924), .A1(n998), .B0(n6), .B1(n909), .Y(n980) );
  INVXL U409 ( .A(n331), .Y(n905) );
  XNOR2XL U410 ( .A(n1194), .B(A[20]), .Y(n1134) );
  XNOR2XL U411 ( .A(n1194), .B(A[19]), .Y(n175) );
  XNOR2XL U412 ( .A(n981), .B(A[13]), .Y(n725) );
  XNOR2XL U413 ( .A(n981), .B(A[12]), .Y(n758) );
  XNOR2XL U414 ( .A(n8), .B(A[10]), .Y(n762) );
  NAND2BXL U415 ( .AN(A[0]), .B(n1184), .Y(n712) );
  XNOR2XL U416 ( .A(n8), .B(A[11]), .Y(n749) );
  OAI22XL U417 ( .A0(n942), .A1(n765), .B0(n751), .B1(n1128), .Y(n785) );
  OAI22XL U418 ( .A0(n812), .A1(n810), .B0(n819), .B1(n752), .Y(n784) );
  XNOR2XL U419 ( .A(n981), .B(A[25]), .Y(n269) );
  XNOR2XL U420 ( .A(n8), .B(A[22]), .Y(n371) );
  OAI22X1 U421 ( .A0(n992), .A1(n340), .B0(n990), .B1(n269), .Y(n329) );
  OAI22XL U422 ( .A0(n924), .A1(n395), .B0(n6), .B1(n334), .Y(n381) );
  XNOR2XL U423 ( .A(n331), .B(A[18]), .Y(n377) );
  ADDFX2 U424 ( .A(n279), .B(n278), .CI(n277), .CO(n263), .S(n319) );
  OAI22XL U425 ( .A0(n1176), .A1(n275), .B0(n1177), .B1(n233), .Y(n279) );
  XNOR2XL U426 ( .A(B[9]), .B(A[21]), .Y(n266) );
  XNOR2XL U427 ( .A(n331), .B(A[20]), .Y(n274) );
  XNOR2X1 U428 ( .A(n1184), .B(A[7]), .Y(n581) );
  OAI22XL U429 ( .A0(n942), .A1(n679), .B0(n647), .B1(n1128), .Y(n674) );
  NAND2BXL U430 ( .AN(A[0]), .B(n668), .Y(n648) );
  XNOR2XL U431 ( .A(n981), .B(A[17]), .Y(n548) );
  XNOR2XL U432 ( .A(n8), .B(A[15]), .Y(n549) );
  CMPR32X1 U433 ( .A(n227), .B(n226), .C(n225), .CO(n206), .S(n260) );
  OAI22XL U434 ( .A0(n912), .A1(n230), .B0(n904), .B1(n195), .Y(n226) );
  OAI22XL U435 ( .A0(n1176), .A1(n232), .B0(n1177), .B1(n194), .Y(n227) );
  OAI22XL U436 ( .A0(n1137), .A1(n231), .B0(n7), .B1(n198), .Y(n222) );
  OAI22XL U437 ( .A0(n1199), .A1(n229), .B0(n1200), .B1(n197), .Y(n223) );
  OAI2BB1XL U438 ( .A0N(n6), .A1N(n924), .B0(n156), .Y(n202) );
  INVXL U439 ( .A(n155), .Y(n156) );
  OAI2BB1XL U440 ( .A0N(n904), .A1N(n912), .B0(n161), .Y(n178) );
  INVXL U441 ( .A(n160), .Y(n161) );
  OAI22XL U442 ( .A0(n1137), .A1(n164), .B0(n7), .B1(n176), .Y(n181) );
  OAI22XL U443 ( .A0(n1199), .A1(n162), .B0(n1200), .B1(n174), .Y(n183) );
  OAI22XL U444 ( .A0(n1176), .A1(n163), .B0(n1177), .B1(n177), .Y(n182) );
  XNOR2XL U445 ( .A(n678), .B(A[2]), .Y(n947) );
  XNOR2XL U446 ( .A(n981), .B(A[1]), .Y(n957) );
  XNOR2XL U447 ( .A(n678), .B(A[3]), .Y(n955) );
  XNOR2XL U448 ( .A(n981), .B(A[4]), .Y(n926) );
  NAND2XL U449 ( .A(n1252), .B(n1257), .Y(n1260) );
  AOI21XL U450 ( .A0(n1258), .A1(n1257), .B0(n1256), .Y(n1259) );
  INVXL U451 ( .A(n1284), .Y(n1256) );
  INVXL U452 ( .A(n1301), .Y(n1261) );
  INVXL U453 ( .A(n1188), .Y(n1170) );
  OAI22XL U454 ( .A0(n1199), .A1(n1157), .B0(n1200), .B1(n1169), .Y(n1172) );
  OAI22XL U455 ( .A0(n1176), .A1(n1139), .B0(n1177), .B1(n1159), .Y(n1162) );
  OAI22XL U456 ( .A0(n1199), .A1(n1140), .B0(n1200), .B1(n1157), .Y(n1161) );
  ADDFX2 U457 ( .A(n880), .B(n879), .CI(n878), .CO(n861), .S(n1045) );
  OAI22X1 U458 ( .A0(n924), .A1(n600), .B0(n6), .B1(n541), .Y(n605) );
  OAI22X1 U459 ( .A0(n924), .A1(n644), .B0(n6), .B1(n600), .Y(n643) );
  OAI22XL U460 ( .A0(n912), .A1(n672), .B0(n995), .B1(n639), .Y(n654) );
  OAI22XL U461 ( .A0(n992), .A1(n649), .B0(n950), .B1(n613), .Y(n675) );
  XNOR2XL U462 ( .A(n678), .B(A[1]), .Y(n941) );
  OAI22XL U463 ( .A0(n992), .A1(n956), .B0(n990), .B1(n936), .Y(n966) );
  XNOR2XL U464 ( .A(n8), .B(A[0]), .Y(n938) );
  ADDFX2 U465 ( .A(n935), .B(n933), .CI(n934), .CO(n974), .S(n973) );
  OAI22XL U466 ( .A0(n992), .A1(n936), .B0(n990), .B1(n926), .Y(n935) );
  NOR2XL U467 ( .A(n1196), .B(n1195), .Y(n1202) );
  XNOR2XL U468 ( .A(n1194), .B(A[24]), .Y(n1195) );
  INVXL U469 ( .A(n1197), .Y(n1198) );
  ADDFX2 U470 ( .A(n1047), .B(n1046), .CI(n1045), .CO(n882), .S(n1052) );
  NAND2X1 U471 ( .A(n120), .B(n119), .Y(n1046) );
  NAND2XL U472 ( .A(n897), .B(n898), .Y(n119) );
  XOR3X2 U473 ( .A(n897), .B(n896), .C(n898), .Y(n1048) );
  NOR2XL U474 ( .A(n1196), .B(n1183), .Y(n1193) );
  INVXL U475 ( .A(n1203), .Y(n1192) );
  XNOR2XL U476 ( .A(n1194), .B(A[23]), .Y(n1183) );
  NAND2X1 U477 ( .A(n121), .B(n123), .Y(n1056) );
  NAND2X1 U478 ( .A(n918), .B(n917), .Y(n1148) );
  OAI22X1 U479 ( .A0(n924), .A1(n486), .B0(n6), .B1(n443), .Y(n491) );
  OAI22X2 U480 ( .A0(n1199), .A1(n487), .B0(n1200), .B1(n444), .Y(n490) );
  OAI22XL U481 ( .A0(n812), .A1(n488), .B0(n819), .B1(n445), .Y(n489) );
  XNOR3X2 U482 ( .A(n508), .B(n81), .C(n506), .Y(n1102) );
  NAND2X1 U483 ( .A(n698), .B(n699), .Y(n106) );
  OAI22XL U484 ( .A0(n942), .A1(A[0]), .B0(n941), .B1(n1128), .Y(n1277) );
  NAND2XL U485 ( .A(n943), .B(n942), .Y(n1276) );
  NAND2BXL U486 ( .AN(A[0]), .B(n678), .Y(n943) );
  NAND2XL U487 ( .A(n1277), .B(n1276), .Y(n1278) );
  INVXL U488 ( .A(n1231), .Y(n1244) );
  INVXL U489 ( .A(n1252), .Y(n1221) );
  INVXL U490 ( .A(n1258), .Y(n1220) );
  INVXL U491 ( .A(n1307), .Y(n1225) );
  NOR2XL U492 ( .A(n1217), .B(n1313), .Y(n1281) );
  INVXL U493 ( .A(n1281), .Y(n1219) );
  NAND2XL U494 ( .A(n1251), .B(n1254), .Y(n1280) );
  NAND2XL U495 ( .A(n1252), .B(n1225), .Y(n1227) );
  AOI21XL U496 ( .A0(n1258), .A1(n1225), .B0(n1224), .Y(n1226) );
  INVXL U497 ( .A(n1308), .Y(n1224) );
  INVXL U498 ( .A(n1305), .Y(n1228) );
  INVXL U499 ( .A(n253), .Y(n293) );
  INVXL U500 ( .A(n291), .Y(n292) );
  INVXL U501 ( .A(n1319), .Y(n323) );
  INVXL U502 ( .A(n1323), .Y(n437) );
  AOI21XL U503 ( .A0(n532), .A1(n535), .B0(n524), .Y(n525) );
  INVXL U504 ( .A(n534), .Y(n524) );
  NAND2XL U505 ( .A(n1349), .B(n1350), .Y(n528) );
  INVXL U506 ( .A(n527), .Y(n529) );
  INVXL U507 ( .A(n532), .Y(n533) );
  INVXL U508 ( .A(n139), .Y(n129) );
  AOI21XL U509 ( .A0(n140), .A1(n126), .B0(n125), .Y(n124) );
  XNOR2XL U510 ( .A(n678), .B(A[10]), .Y(n888) );
  XNOR2XL U511 ( .A(n331), .B(A[0]), .Y(n911) );
  XNOR2XL U512 ( .A(n678), .B(A[9]), .Y(n902) );
  NAND2BXL U513 ( .AN(A[0]), .B(n331), .Y(n903) );
  XNOR2X1 U514 ( .A(n668), .B(A[1]), .Y(n669) );
  XNOR2XL U515 ( .A(n331), .B(A[8]), .Y(n682) );
  XNOR2XL U516 ( .A(n678), .B(A[13]), .Y(n765) );
  XNOR2XL U517 ( .A(n981), .B(A[20]), .Y(n498) );
  XNOR2XL U518 ( .A(n8), .B(A[18]), .Y(n499) );
  XNOR2XL U519 ( .A(n678), .B(A[16]), .Y(n679) );
  XNOR2XL U520 ( .A(n1194), .B(A[15]), .Y(n196) );
  XNOR2XL U521 ( .A(n1194), .B(A[16]), .Y(n154) );
  XNOR2XL U522 ( .A(n1194), .B(A[18]), .Y(n159) );
  OAI22XL U523 ( .A0(n942), .A1(n452), .B0(n390), .B1(n1128), .Y(n451) );
  XNOR2XL U524 ( .A(n981), .B(A[6]), .Y(n991) );
  XNOR2XL U525 ( .A(n8), .B(A[4]), .Y(n984) );
  XNOR2XL U526 ( .A(n922), .B(A[2]), .Y(n998) );
  XNOR2XL U527 ( .A(n678), .B(A[8]), .Y(n996) );
  AOI21XL U528 ( .A0(n1215), .A1(n1214), .B0(n1213), .Y(n1216) );
  INVXL U529 ( .A(n1310), .Y(n1213) );
  NOR2XL U530 ( .A(n1280), .B(n1301), .Y(n1286) );
  AOI21XL U531 ( .A0(n1255), .A1(n1254), .B0(n1253), .Y(n1284) );
  INVXL U532 ( .A(n1304), .Y(n1253) );
  NAND2XL U533 ( .A(n1212), .B(n1312), .Y(n191) );
  NAND2XL U534 ( .A(n1214), .B(n1310), .Y(n150) );
  INVXL U535 ( .A(n359), .Y(n361) );
  OAI2BB1X1 U536 ( .A0N(n537), .A1N(n633), .B0(n632), .Y(n540) );
  AND2XL U537 ( .A(n138), .B(n1336), .Y(n70) );
  ADDFX2 U538 ( .A(n1029), .B(n1028), .CI(n1027), .CO(n1034), .S(n1036) );
  OAI22XL U539 ( .A0(n992), .A1(n991), .B0(n990), .B1(n989), .Y(n1029) );
  OAI22XL U540 ( .A0(n942), .A1(n848), .B0(n820), .B1(n953), .Y(n852) );
  OAI22X1 U541 ( .A0(n821), .A1(n7), .B0(n82), .B1(n117), .Y(n851) );
  NOR2BX1 U542 ( .AN(A[0]), .B(n819), .Y(n853) );
  OAI22XL U543 ( .A0(n992), .A1(n989), .B0(n990), .B1(n892), .Y(n1024) );
  OAI22XL U544 ( .A0(n924), .A1(n909), .B0(n6), .B1(n890), .Y(n1026) );
  XNOR2XL U545 ( .A(n1194), .B(A[22]), .Y(n1173) );
  XNOR2XL U546 ( .A(n1194), .B(A[21]), .Y(n1158) );
  XNOR2XL U547 ( .A(n1138), .B(A[24]), .Y(n1159) );
  OAI22X1 U548 ( .A0(n912), .A1(n756), .B0(n995), .B1(n718), .Y(n761) );
  OAI22X1 U549 ( .A0(n1199), .A1(n720), .B0(n1200), .B1(n719), .Y(n760) );
  OAI22XL U550 ( .A0(n812), .A1(n752), .B0(n819), .B1(n721), .Y(n759) );
  OAI22XL U551 ( .A0(n992), .A1(n788), .B0(n990), .B1(n758), .Y(n790) );
  OAI22XL U552 ( .A0(n912), .A1(n787), .B0(n995), .B1(n756), .Y(n792) );
  OAI22XL U553 ( .A0(n986), .A1(n824), .B0(n9), .B1(n789), .Y(n844) );
  OAI22XL U554 ( .A0(n986), .A1(n789), .B0(n9), .B1(n762), .Y(n816) );
  OAI22XL U555 ( .A0(n869), .A1(n821), .B0(n7), .B1(n813), .Y(n841) );
  XNOR2XL U556 ( .A(n8), .B(A[23]), .Y(n327) );
  ADDFX2 U557 ( .A(n317), .B(n316), .CI(n315), .CO(n320), .S(n348) );
  OAI22XL U558 ( .A0(n1176), .A1(n326), .B0(n1177), .B1(n275), .Y(n316) );
  XNOR2XL U559 ( .A(n678), .B(A[23]), .Y(n452) );
  XNOR2XL U560 ( .A(n678), .B(A[22]), .Y(n495) );
  XNOR2XL U561 ( .A(n678), .B(A[21]), .Y(n567) );
  ADDFX2 U562 ( .A(n417), .B(n416), .CI(n415), .CO(n423), .S(n468) );
  OAI22XL U563 ( .A0(n986), .A1(n414), .B0(n9), .B1(n384), .Y(n415) );
  OAI22XL U564 ( .A0(n992), .A1(n413), .B0(n990), .B1(n383), .Y(n416) );
  OAI22XL U565 ( .A0(n1137), .A1(n412), .B0(n7), .B1(n382), .Y(n417) );
  ADDFX2 U566 ( .A(n420), .B(n419), .CI(n418), .CO(n421), .S(n467) );
  OAI22XL U567 ( .A0(n912), .A1(n449), .B0(n904), .B1(n387), .Y(n420) );
  CMPR32X1 U568 ( .A(n460), .B(n459), .C(n458), .CO(n469), .S(n510) );
  OAI22XL U569 ( .A0(n986), .A1(n457), .B0(n9), .B1(n414), .Y(n458) );
  OAI22XL U570 ( .A0(n992), .A1(n456), .B0(n990), .B1(n413), .Y(n459) );
  OAI22XL U571 ( .A0(n942), .A1(n545), .B0(n568), .B1(n1128), .Y(n571) );
  OAI22XL U572 ( .A0(n986), .A1(n565), .B0(n9), .B1(n564), .Y(n587) );
  XNOR2X1 U573 ( .A(n867), .B(A[6]), .Y(n689) );
  XNOR2XL U574 ( .A(n8), .B(A[12]), .Y(n688) );
  XNOR2X1 U575 ( .A(n766), .B(n28), .Y(n670) );
  XNOR2XL U576 ( .A(n8), .B(A[13]), .Y(n651) );
  XNOR2XL U577 ( .A(n922), .B(A[11]), .Y(n671) );
  XNOR2XL U578 ( .A(n981), .B(A[15]), .Y(n649) );
  XNOR2XL U579 ( .A(n331), .B(A[10]), .Y(n639) );
  XNOR2XL U580 ( .A(n331), .B(A[11]), .Y(n606) );
  NOR2XL U581 ( .A(n234), .B(n546), .Y(n607) );
  OAI2BB1XL U582 ( .A0N(n9), .A1N(n550), .B0(n221), .Y(n239) );
  INVXL U583 ( .A(n220), .Y(n221) );
  OAI22XL U584 ( .A0(n912), .A1(n266), .B0(n904), .B1(n230), .Y(n242) );
  OAI22XL U585 ( .A0(n1199), .A1(n237), .B0(n1200), .B1(n229), .Y(n243) );
  OAI22XL U586 ( .A0(n1137), .A1(n276), .B0(n7), .B1(n238), .Y(n280) );
  OAI22XL U587 ( .A0(n1137), .A1(n238), .B0(n7), .B1(n231), .Y(n265) );
  OAI22XL U588 ( .A0(n1176), .A1(n233), .B0(n1177), .B1(n232), .Y(n264) );
  INVXL U589 ( .A(n179), .Y(n168) );
  OAI22XL U590 ( .A0(n1199), .A1(n166), .B0(n1200), .B1(n162), .Y(n170) );
  OAI22XL U591 ( .A0(n912), .A1(n195), .B0(n904), .B1(n165), .Y(n201) );
  OAI22XL U592 ( .A0(n1176), .A1(n194), .B0(n1177), .B1(n167), .Y(n199) );
  OAI22XL U593 ( .A0(n992), .A1(n383), .B0(n950), .B1(n340), .Y(n386) );
  OAI22X1 U594 ( .A0(n924), .A1(n443), .B0(n6), .B1(n395), .Y(n448) );
  XNOR2X1 U595 ( .A(n8), .B(A[1]), .Y(n937) );
  XNOR2XL U596 ( .A(n981), .B(A[3]), .Y(n936) );
  OAI22XL U597 ( .A0(n942), .A1(n954), .B0(n927), .B1(n1128), .Y(n940) );
  NAND2BXL U598 ( .AN(A[0]), .B(n8), .Y(n928) );
  NAND2BXL U599 ( .AN(A[0]), .B(n922), .Y(n919) );
  ADDFX2 U600 ( .A(n1006), .B(n1005), .CI(n1004), .CO(n1011), .S(n1013) );
  OAI22X1 U601 ( .A0(n924), .A1(n923), .B0(n6), .B1(n999), .Y(n1005) );
  OAI22XL U602 ( .A0(n992), .A1(n926), .B0(n990), .B1(n982), .Y(n1006) );
  ADDFX2 U603 ( .A(n1009), .B(n1008), .CI(n1007), .CO(n1037), .S(n1010) );
  OAI22X1 U604 ( .A0(n986), .A1(n985), .B0(n9), .B1(n984), .Y(n1008) );
  OAI22XL U605 ( .A0(n983), .A1(n982), .B0(n990), .B1(n991), .Y(n1009) );
  ADDFX2 U606 ( .A(n1003), .B(n1002), .CI(n1001), .CO(n1027), .S(n1012) );
  OAI22XL U607 ( .A0(n764), .A1(n997), .B0(n996), .B1(n1128), .Y(n1002) );
  OAI22XL U608 ( .A0(n1000), .A1(n999), .B0(n6), .B1(n998), .Y(n1001) );
  NOR2BXL U609 ( .AN(A[0]), .B(n995), .Y(n1003) );
  NAND2XL U610 ( .A(n1254), .B(n1304), .Y(n1239) );
  NOR2BXL U611 ( .AN(A[0]), .B(n990), .Y(n944) );
  OAI22XL U612 ( .A0(n942), .A1(n941), .B0(n947), .B1(n1128), .Y(n945) );
  CMPR32X1 U613 ( .A(n376), .B(n375), .C(n374), .CO(n350), .S(n393) );
  OAI22X1 U614 ( .A0(n924), .A1(n334), .B0(n6), .B1(n309), .Y(n376) );
  OAI22XL U615 ( .A0(n681), .A1(n335), .B0(n1200), .B1(n311), .Y(n374) );
  ADDFX2 U616 ( .A(n405), .B(n404), .CI(n403), .CO(n392), .S(n424) );
  OAI22XL U617 ( .A0(n912), .A1(n387), .B0(n904), .B1(n377), .Y(n405) );
  OAI22XL U618 ( .A0(n550), .A1(n384), .B0(n9), .B1(n371), .Y(n402) );
  OAI22XL U619 ( .A0(n1176), .A1(n399), .B0(n1177), .B1(n373), .Y(n400) );
  NOR2XL U620 ( .A(n1196), .B(n372), .Y(n401) );
  OAI22XL U621 ( .A0(n986), .A1(n871), .B0(n9), .B1(n824), .Y(n875) );
  OAI22XL U622 ( .A0(n983), .A1(n870), .B0(n990), .B1(n823), .Y(n876) );
  OAI22XL U623 ( .A0(n992), .A1(n892), .B0(n990), .B1(n870), .Y(n893) );
  OAI22XL U624 ( .A0(n1000), .A1(n890), .B0(n6), .B1(n866), .Y(n895) );
  OAI22X1 U625 ( .A0(n868), .A1(n82), .B0(n7), .B1(n117), .Y(n894) );
  ADDFX2 U626 ( .A(n887), .B(n71), .CI(n885), .CO(n878), .S(n1050) );
  OAI22XL U627 ( .A0(n912), .A1(n872), .B0(n995), .B1(n847), .Y(n887) );
  BUFX1 U628 ( .A(n886), .Y(n71) );
  OAI22XL U629 ( .A0(n986), .A1(n891), .B0(n9), .B1(n871), .Y(n901) );
  OAI22XL U630 ( .A0(n912), .A1(n889), .B0(n995), .B1(n872), .Y(n900) );
  ADDFX2 U631 ( .A(n916), .B(n915), .CI(n914), .CO(n1049), .S(n1021) );
  OAI2BB1XL U632 ( .A0N(n101), .A1N(n907), .B0(n100), .Y(n916) );
  NAND2XL U633 ( .A(n103), .B(n908), .Y(n100) );
  NAND2BXL U634 ( .AN(n103), .B(n105), .Y(n101) );
  XOR2X1 U635 ( .A(n105), .B(n103), .Y(n102) );
  OAI2BB1XL U636 ( .A0N(n7), .A1N(n1137), .B0(n1136), .Y(n1154) );
  INVXL U637 ( .A(n1135), .Y(n1136) );
  INVXL U638 ( .A(n1155), .Y(n1141) );
  OAI22XL U639 ( .A0(n1199), .A1(n174), .B0(n1200), .B1(n1140), .Y(n1143) );
  OAI22XL U640 ( .A0(n1176), .A1(n177), .B0(n1177), .B1(n1139), .Y(n1146) );
  XOR3X2 U641 ( .A(n699), .B(n698), .C(n697), .Y(n733) );
  OAI22XL U642 ( .A0(n924), .A1(n763), .B0(n6), .B1(n726), .Y(n778) );
  OAI22XL U643 ( .A0(n992), .A1(n758), .B0(n990), .B1(n725), .Y(n780) );
  OAI22XL U644 ( .A0(n986), .A1(n762), .B0(n9), .B1(n749), .Y(n783) );
  CMPR32X1 U645 ( .A(n330), .B(n329), .C(n328), .CO(n307), .S(n352) );
  OAI2BB1XL U646 ( .A0N(n990), .A1N(n992), .B0(n270), .Y(n328) );
  INVXL U647 ( .A(n269), .Y(n270) );
  CMPR32X1 U648 ( .A(n344), .B(n343), .C(n342), .CO(n353), .S(n410) );
  INVXL U649 ( .A(n329), .Y(n342) );
  OAI22XL U650 ( .A0(n550), .A1(n371), .B0(n9), .B1(n327), .Y(n343) );
  OAI22XL U651 ( .A0(n1176), .A1(n373), .B0(n1177), .B1(n326), .Y(n344) );
  OAI22XL U652 ( .A0(n912), .A1(n377), .B0(n904), .B1(n332), .Y(n347) );
  ADDFX2 U653 ( .A(n320), .B(n319), .CI(n318), .CO(n303), .S(n336) );
  XNOR2XL U654 ( .A(n922), .B(A[18]), .Y(n443) );
  XNOR2X1 U655 ( .A(n766), .B(n91), .Y(n488) );
  XNOR2XL U656 ( .A(n922), .B(A[17]), .Y(n486) );
  OAI22XL U657 ( .A0(n986), .A1(n640), .B0(n9), .B1(n549), .Y(n614) );
  OAI22XL U658 ( .A0(n1137), .A1(n198), .B0(n7), .B1(n193), .Y(n207) );
  OAI22XL U659 ( .A0(n1176), .A1(n167), .B0(n1177), .B1(n163), .Y(n173) );
  XNOR2XL U660 ( .A(n1194), .B(A[17]), .Y(n153) );
  ADDFX2 U661 ( .A(n411), .B(n410), .CI(n409), .CO(n408), .S(n442) );
  OAI22XL U662 ( .A0(n992), .A1(n268), .B0(n950), .B1(n949), .Y(n951) );
  NAND2BXL U663 ( .AN(A[0]), .B(n981), .Y(n949) );
  XNOR2XL U664 ( .A(n981), .B(A[0]), .Y(n948) );
  OAI22XL U665 ( .A0(n942), .A1(n955), .B0(n954), .B1(n953), .Y(n968) );
  NOR2BXL U666 ( .AN(A[0]), .B(n9), .Y(n969) );
  INVXL U667 ( .A(n1291), .Y(n1292) );
  NAND2XL U668 ( .A(n1261), .B(n1302), .Y(n1262) );
  NAND2XL U669 ( .A(n945), .B(n944), .Y(n1272) );
  INVXL U670 ( .A(n1278), .Y(n1274) );
  OAI22XL U671 ( .A0(n1199), .A1(n1169), .B0(n1200), .B1(n1185), .Y(n1182) );
  NAND2X1 U672 ( .A(n131), .B(n133), .Y(n770) );
  OAI21XL U673 ( .A0(n132), .A1(n774), .B0(n772), .Y(n131) );
  BUFX1 U674 ( .A(n773), .Y(n132) );
  OAI2BB1X1 U675 ( .A0N(n825), .A1N(n114), .B0(n113), .Y(n804) );
  ADDFX2 U676 ( .A(n837), .B(n836), .CI(n835), .CO(n828), .S(n858) );
  XOR2X1 U677 ( .A(n86), .B(n85), .Y(n835) );
  XOR2X1 U678 ( .A(n826), .B(n115), .Y(n86) );
  ADDFX2 U679 ( .A(n1097), .B(n1096), .CI(n1095), .CO(n1106), .S(n1114) );
  INVXL U680 ( .A(n643), .Y(n72) );
  NOR2XL U681 ( .A(n952), .B(n951), .Y(n1267) );
  NAND2XL U682 ( .A(n952), .B(n951), .Y(n1268) );
  AOI21XL U683 ( .A0(n1273), .A1(n1274), .B0(n946), .Y(n1270) );
  INVXL U684 ( .A(n1272), .Y(n946) );
  NAND2XL U685 ( .A(n962), .B(n961), .Y(n1264) );
  AOI21XL U686 ( .A0(n1265), .A1(n960), .B0(n963), .Y(n1249) );
  INVXL U687 ( .A(n1264), .Y(n963) );
  NOR2XL U688 ( .A(n971), .B(n970), .Y(n1246) );
  NAND2XL U689 ( .A(n971), .B(n970), .Y(n1247) );
  NAND2XL U690 ( .A(n1207), .B(n1206), .Y(mult_x_1_n58) );
  NAND2XL U691 ( .A(n1205), .B(n1204), .Y(n1206) );
  XNOR2XL U692 ( .A(n1275), .B(n1274), .Y(n1376) );
  NAND2XL U693 ( .A(n1273), .B(n1272), .Y(n1275) );
  NAND2XL U694 ( .A(n135), .B(n1071), .Y(n1072) );
  NOR2XL U695 ( .A(n1130), .B(n1129), .Y(mult_x_1_n151) );
  NOR2XL U696 ( .A(n1150), .B(n1149), .Y(mult_x_1_n136) );
  NOR2XL U697 ( .A(n883), .B(n882), .Y(n881) );
  NOR2XL U698 ( .A(n1190), .B(n1189), .Y(mult_x_1_n109) );
  NAND2XL U699 ( .A(n1190), .B(n1189), .Y(mult_x_1_n110) );
  NOR2XL U700 ( .A(n1179), .B(n1178), .Y(mult_x_1_n120) );
  NAND2XL U701 ( .A(n1179), .B(n1178), .Y(mult_x_1_n121) );
  NOR2XL U702 ( .A(n1164), .B(n1163), .Y(mult_x_1_n129) );
  NAND2XL U703 ( .A(n1164), .B(n1163), .Y(mult_x_1_n130) );
  NAND2XL U704 ( .A(n1150), .B(n1149), .Y(mult_x_1_n137) );
  NOR2XL U705 ( .A(n431), .B(n430), .Y(mult_x_1_n206) );
  NAND2XL U706 ( .A(n858), .B(n857), .Y(mult_x_1_n300) );
  NAND2X1 U707 ( .A(n1055), .B(n1148), .Y(n122) );
  NAND2XL U708 ( .A(n508), .B(n507), .Y(n79) );
  NAND2BXL U709 ( .AN(n508), .B(n81), .Y(n80) );
  OAI21XL U710 ( .A0(n701), .A1(n702), .B0(n700), .Y(n78) );
  NOR2BXL U711 ( .AN(A[0]), .B(n1128), .Y(n1378) );
  XOR2XL U712 ( .A(n1271), .B(n1270), .Y(n1375) );
  NAND2XL U713 ( .A(n1269), .B(n1268), .Y(n1271) );
  INVXL U714 ( .A(n1267), .Y(n1269) );
  XNOR2XL U715 ( .A(n1266), .B(n1265), .Y(n1374) );
  NAND2XL U716 ( .A(n960), .B(n1264), .Y(n1266) );
  XOR2XL U717 ( .A(n1250), .B(n1249), .Y(n1373) );
  NAND2XL U718 ( .A(n1248), .B(n1247), .Y(n1250) );
  INVXL U719 ( .A(n1246), .Y(n1248) );
  XOR2XL U720 ( .A(n1245), .B(n1244), .Y(n1372) );
  NAND2XL U721 ( .A(n1243), .B(n1242), .Y(n1245) );
  INVXL U722 ( .A(n1241), .Y(n1243) );
  NAND2XL U723 ( .A(n1234), .B(n1233), .Y(n1235) );
  NAND2XL U724 ( .A(n1209), .B(n1208), .Y(n1210) );
  OR2X2 U725 ( .A(n766), .B(A[0]), .Y(n68) );
  NOR2X1 U726 ( .A(n1353), .B(n1354), .Y(n631) );
  BUFX3 U727 ( .A(B[3]), .Y(n981) );
  INVX1 U728 ( .A(A[7]), .Y(n110) );
  OAI21XL U729 ( .A0(n433), .A1(n1323), .B0(n1324), .Y(n366) );
  INVX4 U730 ( .A(B[15]), .Y(n714) );
  AOI21X1 U731 ( .A0(n739), .A1(n138), .B0(n738), .Y(n742) );
  OAI21XL U732 ( .A0(n1293), .A1(n1282), .B0(n1290), .Y(n217) );
  CMPR22X1 U733 ( .A(n494), .B(n493), .CO(n461), .S(n504) );
  CMPR22X1 U734 ( .A(n598), .B(n597), .CO(n1089), .S(n585) );
  CMPR22X1 U735 ( .A(n608), .B(n607), .CO(n551), .S(n618) );
  CMPR22X1 U736 ( .A(n646), .B(n645), .CO(n617), .S(n656) );
  OAI22X1 U737 ( .A0(n912), .A1(n165), .B0(n904), .B1(n160), .Y(n179) );
  XNOR2XL U738 ( .A(n1184), .B(A[13]), .Y(n311) );
  OAI22X1 U739 ( .A0(n1176), .A1(n766), .B0(n1177), .B1(n68), .Y(n817) );
  OAI22X1 U740 ( .A0(n924), .A1(n228), .B0(n6), .B1(n155), .Y(n203) );
  CMPR22X1 U741 ( .A(n988), .B(n987), .CO(n1007), .S(n1015) );
  OAI22X1 U742 ( .A0(n924), .A1(n920), .B0(n6), .B1(n919), .Y(n987) );
  NAND2X1 U743 ( .A(n253), .B(n147), .Y(n1282) );
  OAI22X1 U744 ( .A0(n942), .A1(n751), .B0(n711), .B1(n1128), .Y(n750) );
  CMPR22X1 U745 ( .A(n389), .B(n388), .CO(n404), .S(n419) );
  AOI21X1 U746 ( .A0(n739), .A1(n139), .B0(n140), .Y(n130) );
  XOR2X1 U747 ( .A(n742), .B(n741), .Y(PRODUCT[18]) );
  XNOR2X1 U748 ( .A(n540), .B(n539), .Y(PRODUCT[22]) );
  XNOR3X2 U749 ( .A(n643), .B(n642), .C(n75), .Y(n659) );
  INVX8 U750 ( .A(n1138), .Y(n766) );
  OAI22X1 U751 ( .A0(n75), .A1(n74), .B0(n73), .B1(n72), .Y(n622) );
  NOR2XL U752 ( .A(n642), .B(n643), .Y(n74) );
  AOI2BB1X1 U753 ( .A0N(n819), .A1N(n602), .B0(n76), .Y(n75) );
  NOR2X1 U754 ( .A(n641), .B(n812), .Y(n76) );
  NAND2X1 U755 ( .A(n78), .B(n77), .Y(n1126) );
  INVX1 U756 ( .A(n507), .Y(n81) );
  XOR2X2 U757 ( .A(B[10]), .B(B[11]), .Y(n83) );
  XOR2X4 U758 ( .A(B[10]), .B(n84), .Y(n454) );
  CLKINVX3 U759 ( .A(B[9]), .Y(n84) );
  XNOR2X1 U760 ( .A(n766), .B(n90), .Y(n582) );
  XNOR2X1 U761 ( .A(n766), .B(n92), .Y(n543) );
  XNOR2X1 U762 ( .A(n766), .B(n110), .Y(n602) );
  XNOR2X1 U763 ( .A(n766), .B(n93), .Y(n641) );
  XNOR2X1 U764 ( .A(n766), .B(n94), .Y(n684) );
  XNOR2X1 U765 ( .A(n766), .B(n118), .Y(n810) );
  XNOR2X1 U766 ( .A(n766), .B(n96), .Y(n194) );
  XNOR2X1 U767 ( .A(n766), .B(n104), .Y(n811) );
  XNOR2X1 U768 ( .A(n766), .B(n97), .Y(n752) );
  XNOR2X1 U769 ( .A(n766), .B(n98), .Y(n373) );
  OAI22X1 U770 ( .A0(n82), .A1(n689), .B0(n7), .B1(n109), .Y(n687) );
  OAI22X2 U771 ( .A0(n7), .A1(n611), .B0(n82), .B1(n109), .Y(n677) );
  XOR2X1 U772 ( .A(n867), .B(n110), .Y(n109) );
  XOR2X1 U773 ( .A(n116), .B(n750), .Y(n782) );
  OAI22X1 U774 ( .A0(n1199), .A1(n714), .B0(n713), .B1(n712), .Y(n116) );
  NAND2X1 U775 ( .A(n739), .B(n128), .Y(n127) );
  XOR2X1 U776 ( .A(n773), .B(n774), .Y(n134) );
  OAI22X4 U777 ( .A0(n1199), .A1(n612), .B0(n1200), .B1(n601), .Y(n642) );
  XNOR2X1 U778 ( .A(n1062), .B(n1061), .Y(n1367) );
  XNOR2X1 U779 ( .A(n439), .B(n438), .Y(PRODUCT[27]) );
  XOR2X1 U780 ( .A(n217), .B(n69), .Y(PRODUCT[33]) );
  XNOR2X2 U781 ( .A(B[16]), .B(B[15]), .Y(n234) );
  XOR2X2 U782 ( .A(n1293), .B(n362), .Y(PRODUCT[29]) );
  NAND2X1 U783 ( .A(n152), .B(n398), .Y(n397) );
  XNOR2X2 U784 ( .A(B[12]), .B(B[11]), .Y(n398) );
  OAI22X1 U785 ( .A0(n82), .A1(n611), .B0(n7), .B1(n547), .Y(n616) );
  OAI22X1 U786 ( .A0(n82), .A1(n560), .B0(n7), .B1(n497), .Y(n592) );
  OAI2BB1X1 U787 ( .A0N(n537), .A1N(n517), .B0(n39), .Y(n521) );
  OR2X2 U788 ( .A(n1019), .B(n1018), .Y(n135) );
  AOI21XL U789 ( .A0(n1287), .A1(n1286), .B0(n1285), .Y(n1288) );
  INVX1 U790 ( .A(n1344), .Y(n859) );
  XNOR2XL U791 ( .A(n678), .B(A[5]), .Y(n927) );
  XNOR2XL U792 ( .A(n678), .B(A[20]), .Y(n568) );
  XNOR2XL U793 ( .A(n678), .B(A[17]), .Y(n647) );
  XNOR2XL U794 ( .A(n678), .B(A[4]), .Y(n954) );
  XNOR2XL U795 ( .A(n1168), .B(A[22]), .Y(n1157) );
  OAI22X1 U796 ( .A0(n1199), .A1(n680), .B0(n1200), .B1(n667), .Y(n693) );
  OAI22X2 U797 ( .A0(n1199), .A1(n601), .B0(n1200), .B1(n542), .Y(n604) );
  INVX4 U798 ( .A(n1339), .Y(n832) );
  NAND2X2 U799 ( .A(n832), .B(n1295), .Y(n799) );
  CLKINVX3 U800 ( .A(n1340), .Y(n136) );
  AOI21X4 U801 ( .A0(n832), .A1(n1296), .B0(n136), .Y(n798) );
  INVX4 U802 ( .A(n141), .Y(n739) );
  NOR2X1 U803 ( .A(n523), .B(n527), .Y(n142) );
  NOR2X1 U804 ( .A(n1347), .B(n1348), .Y(n475) );
  OAI21XL U805 ( .A0(n1325), .A1(n518), .B0(n1326), .Y(n365) );
  OAI21XL U806 ( .A0(n1321), .A1(n1324), .B0(n1322), .Y(n143) );
  AOI21XL U807 ( .A0(n144), .A1(n365), .B0(n143), .Y(n145) );
  NOR2X1 U808 ( .A(n1346), .B(n1345), .Y(n359) );
  NOR2XL U809 ( .A(n1317), .B(n1315), .Y(n147) );
  NOR2XL U810 ( .A(n1282), .B(n1313), .Y(n187) );
  NAND2XL U811 ( .A(n187), .B(n1212), .Y(n149) );
  NAND2X1 U812 ( .A(n1346), .B(n1345), .Y(n360) );
  OAI21XL U813 ( .A0(n1319), .A1(n360), .B0(n1320), .Y(n291) );
  OAI21XL U814 ( .A0(n1315), .A1(n1318), .B0(n1316), .Y(n146) );
  AOI21X1 U815 ( .A0(n291), .A1(n147), .B0(n146), .Y(n1290) );
  OAI21XL U816 ( .A0(n1290), .A1(n1313), .B0(n1314), .Y(n188) );
  OAI21XL U817 ( .A0(n1293), .A1(n149), .B0(n148), .Y(n151) );
  XOR2X1 U818 ( .A(B[12]), .B(B[13]), .Y(n152) );
  BUFX3 U819 ( .A(n397), .Y(n1176) );
  XNOR2X1 U820 ( .A(n1138), .B(A[20]), .Y(n167) );
  BUFX3 U821 ( .A(n398), .Y(n1177) );
  XNOR2X1 U822 ( .A(n1138), .B(A[21]), .Y(n163) );
  BUFX3 U823 ( .A(n234), .Y(n1196) );
  XNOR2XL U824 ( .A(n922), .B(A[24]), .Y(n228) );
  INVX8 U825 ( .A(n920), .Y(n922) );
  XNOR2XL U826 ( .A(n922), .B(A[25]), .Y(n155) );
  XOR2X1 U827 ( .A(B[14]), .B(B[15]), .Y(n157) );
  XNOR2X2 U828 ( .A(B[14]), .B(B[13]), .Y(n713) );
  XNOR2XL U829 ( .A(n1168), .B(A[18]), .Y(n166) );
  XNOR2X1 U830 ( .A(n867), .B(A[22]), .Y(n193) );
  XNOR2XL U831 ( .A(n867), .B(A[23]), .Y(n164) );
  OAI22XL U832 ( .A0(n1137), .A1(n193), .B0(n7), .B1(n164), .Y(n169) );
  XOR2X1 U833 ( .A(B[8]), .B(B[9]), .Y(n158) );
  XNOR2X4 U834 ( .A(B[8]), .B(B[7]), .Y(n904) );
  NAND2X2 U835 ( .A(n158), .B(n904), .Y(n906) );
  XNOR2XL U836 ( .A(n331), .B(A[25]), .Y(n160) );
  XNOR2X1 U837 ( .A(n1138), .B(A[22]), .Y(n177) );
  XNOR2X1 U838 ( .A(n867), .B(A[24]), .Y(n176) );
  OAI22XL U839 ( .A0(n1199), .A1(n197), .B0(n1200), .B1(n166), .Y(n200) );
  CMPR32X1 U840 ( .A(n170), .B(n169), .C(n168), .CO(n186), .S(n209) );
  CMPR32X1 U841 ( .A(n173), .B(n172), .C(n171), .CO(n213), .S(n208) );
  INVX8 U842 ( .A(n850), .Y(n867) );
  XNOR2X1 U843 ( .A(n867), .B(A[25]), .Y(n1135) );
  OAI22X1 U844 ( .A0(n1137), .A1(n176), .B0(n7), .B1(n1135), .Y(n1155) );
  CMPR32X1 U845 ( .A(n180), .B(n179), .C(n178), .CO(n1145), .S(n185) );
  CMPR32X1 U846 ( .A(n183), .B(n182), .C(n181), .CO(n1144), .S(n184) );
  CMPR32X1 U847 ( .A(n186), .B(n185), .C(n184), .CO(n1131), .S(n212) );
  NAND2XL U848 ( .A(n1130), .B(n1129), .Y(mult_x_1_n152) );
  INVXL U849 ( .A(n187), .Y(n190) );
  INVXL U850 ( .A(n188), .Y(n189) );
  XNOR2X1 U851 ( .A(n867), .B(A[21]), .Y(n198) );
  XNOR2X1 U852 ( .A(n1138), .B(A[18]), .Y(n232) );
  XNOR2XL U853 ( .A(n331), .B(A[22]), .Y(n230) );
  INVXL U854 ( .A(n203), .Y(n225) );
  CMPR32X1 U855 ( .A(n201), .B(n200), .C(n199), .CO(n210), .S(n247) );
  CMPR32X1 U856 ( .A(n204), .B(n203), .C(n202), .CO(n171), .S(n246) );
  ADDFHX1 U857 ( .A(n207), .B(n206), .CI(n205), .CO(n250), .S(n245) );
  CMPR32X1 U858 ( .A(n210), .B(n209), .C(n208), .CO(n211), .S(n248) );
  CMPR32X1 U859 ( .A(n213), .B(n212), .C(n211), .CO(n1130), .S(n214) );
  NOR2XL U860 ( .A(n215), .B(n214), .Y(mult_x_1_n160) );
  NAND2XL U861 ( .A(n215), .B(n214), .Y(mult_x_1_n161) );
  CLKINVX3 U862 ( .A(B[5]), .Y(n929) );
  OAI22X1 U863 ( .A0(n986), .A1(n271), .B0(n9), .B1(n220), .Y(n240) );
  CMPR32X1 U864 ( .A(n224), .B(n223), .C(n222), .CO(n205), .S(n261) );
  XNOR2X1 U865 ( .A(n922), .B(A[23]), .Y(n236) );
  OAI22XL U866 ( .A0(n924), .A1(n236), .B0(n6), .B1(n228), .Y(n244) );
  XNOR2X1 U867 ( .A(n1138), .B(A[17]), .Y(n233) );
  XNOR2XL U868 ( .A(n1194), .B(A[13]), .Y(n235) );
  NOR2XL U869 ( .A(n234), .B(n235), .Y(n278) );
  INVXL U870 ( .A(n240), .Y(n277) );
  XNOR2X1 U871 ( .A(n922), .B(A[22]), .Y(n273) );
  OAI22XL U872 ( .A0(n924), .A1(n273), .B0(n6), .B1(n236), .Y(n282) );
  INVX8 U873 ( .A(n714), .Y(n1184) );
  OAI22X1 U874 ( .A0(n1199), .A1(n272), .B0(n1200), .B1(n237), .Y(n281) );
  XNOR2XL U875 ( .A(n867), .B(A[18]), .Y(n276) );
  CMPR32X1 U876 ( .A(n241), .B(n240), .C(n239), .CO(n262), .S(n301) );
  CMPR32X1 U877 ( .A(n244), .B(n243), .C(n242), .CO(n285), .S(n300) );
  CMPR32X1 U878 ( .A(n247), .B(n246), .C(n245), .CO(n249), .S(n286) );
  CMPR32X1 U879 ( .A(n250), .B(n249), .C(n248), .CO(n215), .S(n251) );
  NOR2XL U880 ( .A(n252), .B(n251), .Y(mult_x_1_n169) );
  NAND2XL U881 ( .A(n252), .B(n251), .Y(mult_x_1_n170) );
  AOI21XL U882 ( .A0(n291), .A1(n294), .B0(n254), .Y(n255) );
  XNOR2X1 U883 ( .A(n259), .B(n258), .Y(PRODUCT[32]) );
  CMPR32X1 U884 ( .A(n262), .B(n261), .C(n260), .CO(n288), .S(n299) );
  CMPR32X1 U885 ( .A(n265), .B(n264), .C(n263), .CO(n284), .S(n305) );
  XNOR2XL U886 ( .A(n1194), .B(A[12]), .Y(n267) );
  NOR2XL U887 ( .A(n234), .B(n267), .Y(n330) );
  INVXL U888 ( .A(n981), .Y(n268) );
  OAI22XL U889 ( .A0(n550), .A1(n327), .B0(n9), .B1(n271), .Y(n314) );
  OAI22X1 U890 ( .A0(n1199), .A1(n311), .B0(n1200), .B1(n272), .Y(n313) );
  XNOR2X1 U891 ( .A(n922), .B(A[21]), .Y(n309) );
  OAI22XL U892 ( .A0(n924), .A1(n309), .B0(n6), .B1(n273), .Y(n312) );
  XNOR2XL U893 ( .A(n331), .B(A[19]), .Y(n332) );
  BUFX3 U894 ( .A(n904), .Y(n995) );
  OAI22XL U895 ( .A0(n912), .A1(n332), .B0(n995), .B1(n274), .Y(n317) );
  XNOR2X1 U896 ( .A(n1138), .B(A[15]), .Y(n326) );
  XNOR2XL U897 ( .A(n867), .B(A[17]), .Y(n333) );
  OAI22XL U898 ( .A0(n1137), .A1(n333), .B0(n7), .B1(n276), .Y(n315) );
  ADDFHX1 U899 ( .A(n285), .B(n284), .CI(n283), .CO(n287), .S(n297) );
  CMPR32X1 U900 ( .A(n288), .B(n287), .C(n286), .CO(n252), .S(n289) );
  NOR2XL U901 ( .A(n290), .B(n289), .Y(mult_x_1_n176) );
  NAND2XL U902 ( .A(n290), .B(n289), .Y(mult_x_1_n177) );
  OAI21X1 U903 ( .A0(n1293), .A1(n293), .B0(n292), .Y(n296) );
  NAND2X1 U904 ( .A(n294), .B(n1318), .Y(n295) );
  ADDFHX1 U905 ( .A(n299), .B(n298), .CI(n297), .CO(n290), .S(n322) );
  CMPR32X1 U906 ( .A(n302), .B(n301), .C(n300), .CO(n283), .S(n356) );
  CMPR32X1 U907 ( .A(n305), .B(n304), .C(n303), .CO(n298), .S(n355) );
  XNOR2X1 U908 ( .A(n922), .B(A[20]), .Y(n334) );
  NOR2XL U909 ( .A(n234), .B(n310), .Y(n375) );
  NOR2XL U910 ( .A(n322), .B(n321), .Y(mult_x_1_n183) );
  NAND2XL U911 ( .A(n322), .B(n321), .Y(mult_x_1_n184) );
  OAI21X1 U912 ( .A0(n1293), .A1(n359), .B0(n360), .Y(n325) );
  NAND2X1 U913 ( .A(n323), .B(n1320), .Y(n324) );
  XNOR2X2 U914 ( .A(n325), .B(n324), .Y(PRODUCT[30]) );
  XNOR2X1 U915 ( .A(n867), .B(A[16]), .Y(n339) );
  OAI22XL U916 ( .A0(n1137), .A1(n339), .B0(n7), .B1(n333), .Y(n346) );
  XNOR2X1 U917 ( .A(n922), .B(A[19]), .Y(n395) );
  XNOR2X1 U918 ( .A(n1184), .B(A[11]), .Y(n396) );
  OR2X2 U919 ( .A(n381), .B(n380), .Y(n345) );
  XNOR2X1 U920 ( .A(n867), .B(A[15]), .Y(n382) );
  BUFX3 U921 ( .A(n953), .Y(n1128) );
  BUFX3 U922 ( .A(n764), .Y(n942) );
  CMPR32X1 U923 ( .A(n347), .B(n346), .C(n345), .CO(n351), .S(n409) );
  CMPR32X1 U924 ( .A(n353), .B(n352), .C(n351), .CO(n1076), .S(n406) );
  ADDFHX1 U925 ( .A(n356), .B(n355), .CI(n354), .CO(n321), .S(n357) );
  NOR2XL U926 ( .A(n358), .B(n357), .Y(mult_x_1_n194) );
  NAND2XL U927 ( .A(n358), .B(n357), .Y(mult_x_1_n195) );
  NAND2X1 U928 ( .A(n361), .B(n360), .Y(n362) );
  INVXL U929 ( .A(n363), .Y(n432) );
  NOR2XL U930 ( .A(n432), .B(n1323), .Y(n367) );
  INVX1 U931 ( .A(n364), .Y(n517) );
  NAND2XL U932 ( .A(n367), .B(n517), .Y(n368) );
  INVXL U933 ( .A(n365), .Y(n433) );
  INVXL U934 ( .A(n1321), .Y(n369) );
  OAI22X1 U935 ( .A0(n942), .A1(n390), .B0(n378), .B1(n1128), .Y(n389) );
  NOR2XL U936 ( .A(n234), .B(n379), .Y(n388) );
  XNOR2X1 U937 ( .A(n867), .B(A[14]), .Y(n412) );
  XNOR2XL U938 ( .A(n331), .B(A[16]), .Y(n449) );
  XNOR2XL U939 ( .A(n668), .B(A[8]), .Y(n391) );
  NOR2XL U940 ( .A(n234), .B(n391), .Y(n450) );
  XNOR2X1 U941 ( .A(n1184), .B(A[10]), .Y(n444) );
  OAI22X4 U942 ( .A0(n1199), .A1(n444), .B0(n1200), .B1(n396), .Y(n447) );
  BUFX3 U943 ( .A(n397), .Y(n812) );
  BUFX3 U944 ( .A(n398), .Y(n819) );
  OAI22X1 U945 ( .A0(n812), .A1(n445), .B0(n819), .B1(n399), .Y(n446) );
  CMPR32X1 U946 ( .A(n402), .B(n401), .C(n400), .CO(n394), .S(n425) );
  XNOR2X1 U947 ( .A(n867), .B(A[13]), .Y(n455) );
  OAI22X1 U948 ( .A0(n1137), .A1(n455), .B0(n7), .B1(n412), .Y(n460) );
  ADDFHX1 U949 ( .A(n423), .B(n422), .CI(n421), .CO(n429), .S(n471) );
  CMPR32X1 U950 ( .A(n426), .B(n425), .C(n424), .CO(n427), .S(n470) );
  NAND2XL U951 ( .A(n517), .B(n363), .Y(n436) );
  INVXL U952 ( .A(n433), .Y(n434) );
  ADDFHX1 U953 ( .A(n442), .B(n441), .CI(n440), .CO(n430), .S(n474) );
  XNOR2X1 U954 ( .A(n1184), .B(A[9]), .Y(n487) );
  XNOR2XL U955 ( .A(n331), .B(A[15]), .Y(n492) );
  OAI22XL U956 ( .A0(n912), .A1(n492), .B0(n904), .B1(n449), .Y(n463) );
  ADDHXL U957 ( .A(n451), .B(n450), .CO(n418), .S(n462) );
  OAI22X1 U958 ( .A0(n942), .A1(n495), .B0(n452), .B1(n1128), .Y(n494) );
  XNOR2X1 U959 ( .A(n668), .B(A[7]), .Y(n453) );
  NOR2XL U960 ( .A(n234), .B(n453), .Y(n493) );
  XNOR2X1 U961 ( .A(n867), .B(A[12]), .Y(n497) );
  OAI22X2 U962 ( .A0(n992), .A1(n498), .B0(n990), .B1(n456), .Y(n501) );
  OAI22X1 U963 ( .A0(n986), .A1(n499), .B0(n9), .B1(n457), .Y(n500) );
  CMPR32X1 U964 ( .A(n463), .B(n461), .C(n462), .CO(n464), .S(n509) );
  ADDFHX1 U965 ( .A(n469), .B(n468), .CI(n467), .CO(n472), .S(n512) );
  ADDFHX1 U966 ( .A(n472), .B(n471), .CI(n470), .CO(n441), .S(n483) );
  NOR2XL U967 ( .A(n474), .B(n473), .Y(mult_x_1_n215) );
  NAND2XL U968 ( .A(n517), .B(n519), .Y(n479) );
  INVXL U969 ( .A(n518), .Y(n476) );
  OAI21XL U970 ( .A0(n635), .A1(n479), .B0(n478), .Y(n482) );
  INVXL U971 ( .A(n1325), .Y(n480) );
  XNOR2X1 U972 ( .A(n482), .B(n481), .Y(PRODUCT[26]) );
  ADDFHX1 U973 ( .A(n485), .B(n484), .CI(n483), .CO(n473), .S(n516) );
  XNOR2X1 U974 ( .A(n922), .B(A[16]), .Y(n578) );
  XNOR2X1 U975 ( .A(n1184), .B(A[8]), .Y(n580) );
  OAI22X1 U976 ( .A0(n812), .A1(n582), .B0(n819), .B1(n488), .Y(n1086) );
  XNOR2XL U977 ( .A(n331), .B(A[14]), .Y(n593) );
  OAI22XL U978 ( .A0(n912), .A1(n593), .B0(n904), .B1(n492), .Y(n505) );
  XNOR2XL U979 ( .A(n668), .B(A[6]), .Y(n496) );
  NOR2XL U980 ( .A(n234), .B(n496), .Y(n595) );
  OAI22X1 U981 ( .A0(n986), .A1(n564), .B0(n9), .B1(n499), .Y(n590) );
  CMPR32X1 U982 ( .A(n505), .B(n504), .C(n503), .CO(n506), .S(n1098) );
  CMPR32X1 U983 ( .A(n514), .B(n513), .C(n512), .CO(n484), .S(n1080) );
  NOR2XL U984 ( .A(n516), .B(n515), .Y(mult_x_1_n226) );
  NAND2XL U985 ( .A(n516), .B(n515), .Y(mult_x_1_n227) );
  NAND2XL U986 ( .A(n522), .B(n535), .Y(n526) );
  OAI21XL U987 ( .A0(n635), .A1(n526), .B0(n525), .Y(n531) );
  NAND2X1 U988 ( .A(n529), .B(n528), .Y(n530) );
  XNOR2X2 U989 ( .A(n531), .B(n530), .Y(PRODUCT[24]) );
  INVXL U990 ( .A(n1327), .Y(n538) );
  XNOR2X1 U991 ( .A(n1184), .B(A[6]), .Y(n542) );
  OAI22XL U992 ( .A0(n812), .A1(n602), .B0(n819), .B1(n543), .Y(n603) );
  XNOR2X1 U993 ( .A(n922), .B(A[15]), .Y(n579) );
  OAI22X1 U994 ( .A0(n924), .A1(n541), .B0(n6), .B1(n579), .Y(n577) );
  OAI22X2 U995 ( .A0(n1199), .A1(n542), .B0(n1200), .B1(n581), .Y(n576) );
  XNOR2XL U996 ( .A(n331), .B(A[12]), .Y(n566) );
  OAI22XL U997 ( .A0(n906), .A1(n606), .B0(n995), .B1(n566), .Y(n553) );
  XNOR2XL U998 ( .A(n668), .B(A[4]), .Y(n544) );
  NOR2XL U999 ( .A(n234), .B(n544), .Y(n570) );
  OAI22X1 U1000 ( .A0(n942), .A1(n609), .B0(n545), .B1(n1128), .Y(n608) );
  XNOR2X1 U1001 ( .A(n668), .B(A[3]), .Y(n546) );
  XNOR2X1 U1002 ( .A(n867), .B(A[8]), .Y(n611) );
  XNOR2XL U1003 ( .A(n981), .B(A[16]), .Y(n613) );
  OAI22X2 U1004 ( .A0(n992), .A1(n613), .B0(n990), .B1(n548), .Y(n615) );
  XNOR2X1 U1005 ( .A(n867), .B(A[10]), .Y(n561) );
  OAI22X1 U1006 ( .A0(n869), .A1(n547), .B0(n7), .B1(n561), .Y(n559) );
  OAI22X1 U1007 ( .A0(n992), .A1(n548), .B0(n990), .B1(n563), .Y(n558) );
  OAI22XL U1008 ( .A0(n550), .A1(n549), .B0(n9), .B1(n565), .Y(n557) );
  CMPR32X1 U1009 ( .A(n553), .B(n551), .C(n552), .CO(n554), .S(n623) );
  CMPR32X1 U1010 ( .A(n556), .B(n555), .C(n554), .CO(n1121), .S(n627) );
  OAI22X1 U1011 ( .A0(n869), .A1(n561), .B0(n454), .B1(n560), .Y(n589) );
  OAI22X1 U1012 ( .A0(n992), .A1(n563), .B0(n990), .B1(n562), .Y(n588) );
  XNOR2XL U1013 ( .A(n331), .B(A[13]), .Y(n594) );
  OAI22XL U1014 ( .A0(n906), .A1(n566), .B0(n995), .B1(n594), .Y(n586) );
  OAI22X1 U1015 ( .A0(n942), .A1(n568), .B0(n567), .B1(n1128), .Y(n598) );
  XNOR2XL U1016 ( .A(n668), .B(A[5]), .Y(n569) );
  NOR2XL U1017 ( .A(n234), .B(n569), .Y(n597) );
  ADDHXL U1018 ( .A(n571), .B(n570), .CO(n584), .S(n552) );
  ADDFHX1 U1019 ( .A(n574), .B(n573), .CI(n572), .CO(n1112), .S(n626) );
  OAI22X1 U1020 ( .A0(n924), .A1(n579), .B0(n6), .B1(n578), .Y(n1085) );
  OAI22X2 U1021 ( .A0(n1199), .A1(n581), .B0(n1200), .B1(n580), .Y(n1084) );
  OAI22X1 U1022 ( .A0(n812), .A1(n583), .B0(n819), .B1(n582), .Y(n1083) );
  CMPR32X1 U1023 ( .A(n586), .B(n585), .C(n584), .CO(n1107), .S(n572) );
  OAI22XL U1024 ( .A0(n912), .A1(n594), .B0(n904), .B1(n593), .Y(n1091) );
  ADDHXL U1025 ( .A(n596), .B(n595), .CO(n503), .S(n1090) );
  XNOR2X1 U1026 ( .A(n922), .B(A[12]), .Y(n644) );
  OAI22XL U1027 ( .A0(n912), .A1(n639), .B0(n995), .B1(n606), .Y(n619) );
  OAI22X1 U1028 ( .A0(n942), .A1(n647), .B0(n609), .B1(n1128), .Y(n646) );
  XNOR2XL U1029 ( .A(n668), .B(A[2]), .Y(n610) );
  NOR2XL U1030 ( .A(n234), .B(n610), .Y(n645) );
  XNOR2X1 U1031 ( .A(n1184), .B(A[3]), .Y(n667) );
  OAI22X2 U1032 ( .A0(n1199), .A1(n667), .B0(n1200), .B1(n612), .Y(n676) );
  CMPR32X1 U1033 ( .A(n619), .B(n618), .C(n617), .CO(n620), .S(n661) );
  ADDFHX1 U1034 ( .A(n625), .B(n624), .CI(n623), .CO(n628), .S(n664) );
  NOR2XL U1035 ( .A(n630), .B(n629), .Y(mult_x_1_n262) );
  INVXL U1036 ( .A(n631), .Y(n633) );
  NAND2X1 U1037 ( .A(n633), .B(n632), .Y(n634) );
  XOR2X1 U1038 ( .A(n635), .B(n634), .Y(PRODUCT[21]) );
  INVXL U1039 ( .A(n1329), .Y(n636) );
  XNOR2XL U1040 ( .A(n331), .B(A[9]), .Y(n672) );
  OAI22XL U1041 ( .A0(n812), .A1(n670), .B0(n819), .B1(n641), .Y(n652) );
  OAI22XL U1042 ( .A0(n924), .A1(n671), .B0(n6), .B1(n644), .Y(n657) );
  XNOR2X1 U1043 ( .A(n981), .B(A[14]), .Y(n683) );
  OAI22X2 U1044 ( .A0(n992), .A1(n683), .B0(n990), .B1(n649), .Y(n686) );
  OAI22X1 U1045 ( .A0(n986), .A1(n688), .B0(n9), .B1(n651), .Y(n685) );
  CMPR32X1 U1046 ( .A(n654), .B(n653), .C(n652), .CO(n660), .S(n698) );
  CMPR32X1 U1047 ( .A(n657), .B(n656), .C(n655), .CO(n658), .S(n697) );
  CMPR32X1 U1048 ( .A(n660), .B(n659), .C(n658), .CO(n1127), .S(n701) );
  CMPR32X1 U1049 ( .A(n666), .B(n665), .C(n664), .CO(n1123), .S(n1125) );
  XNOR2X1 U1050 ( .A(n1184), .B(A[2]), .Y(n680) );
  NOR2XL U1051 ( .A(n234), .B(n669), .Y(n692) );
  OAI22XL U1052 ( .A0(n812), .A1(n684), .B0(n819), .B1(n670), .Y(n691) );
  XNOR2XL U1053 ( .A(n922), .B(A[10]), .Y(n690) );
  OAI22XL U1054 ( .A0(n924), .A1(n690), .B0(n6), .B1(n671), .Y(n696) );
  OAI22XL U1055 ( .A0(n912), .A1(n682), .B0(n995), .B1(n672), .Y(n695) );
  ADDHXL U1056 ( .A(n674), .B(n673), .CO(n655), .S(n694) );
  XNOR2X1 U1057 ( .A(n1184), .B(A[1]), .Y(n719) );
  OAI22X1 U1058 ( .A0(n912), .A1(n718), .B0(n995), .B1(n682), .Y(n729) );
  OAI22X1 U1059 ( .A0(n992), .A1(n725), .B0(n990), .B1(n683), .Y(n728) );
  OAI22X1 U1060 ( .A0(n812), .A1(n721), .B0(n819), .B1(n684), .Y(n727) );
  OAI22X1 U1061 ( .A0(n986), .A1(n749), .B0(n9), .B1(n688), .Y(n732) );
  XNOR2X1 U1062 ( .A(n922), .B(A[9]), .Y(n726) );
  OAI22XL U1063 ( .A0(n924), .A1(n726), .B0(n6), .B1(n690), .Y(n730) );
  ADDFX2 U1064 ( .A(n693), .B(n692), .CI(n691), .CO(n710), .S(n747) );
  CMPR32X1 U1065 ( .A(n696), .B(n695), .C(n694), .CO(n709), .S(n746) );
  NOR2XL U1066 ( .A(n704), .B(n703), .Y(mult_x_1_n273) );
  NAND2XL U1067 ( .A(n704), .B(n703), .Y(mult_x_1_n274) );
  CMPR32X1 U1068 ( .A(n707), .B(n706), .C(n705), .CO(n703), .S(n737) );
  CMPR32X1 U1069 ( .A(n710), .B(n709), .C(n708), .CO(n707), .S(n745) );
  XNOR2X1 U1070 ( .A(n1184), .B(A[0]), .Y(n720) );
  XNOR2X1 U1071 ( .A(n867), .B(A[4]), .Y(n757) );
  XNOR2XL U1072 ( .A(n922), .B(A[8]), .Y(n763) );
  CMPR32X1 U1073 ( .A(n729), .B(n728), .C(n727), .CO(n723), .S(n776) );
  NOR2XL U1074 ( .A(n737), .B(n736), .Y(mult_x_1_n276) );
  NAND2XL U1075 ( .A(n737), .B(n736), .Y(mult_x_1_n277) );
  INVXL U1076 ( .A(n1336), .Y(n738) );
  INVXL U1077 ( .A(n1333), .Y(n740) );
  XNOR2X1 U1078 ( .A(n867), .B(A[3]), .Y(n813) );
  OAI22X1 U1079 ( .A0(n82), .A1(n813), .B0(n7), .B1(n757), .Y(n791) );
  XNOR2XL U1080 ( .A(n981), .B(A[11]), .Y(n788) );
  XNOR2X1 U1081 ( .A(n922), .B(A[7]), .Y(n809) );
  OAI22XL U1082 ( .A0(n924), .A1(n809), .B0(n6), .B1(n763), .Y(n815) );
  NOR2XL U1083 ( .A(n771), .B(n770), .Y(mult_x_1_n281) );
  NAND2XL U1084 ( .A(n771), .B(n770), .Y(mult_x_1_n282) );
  CMPR32X1 U1085 ( .A(n777), .B(n776), .C(n775), .CO(n767), .S(n805) );
  CMPR32X1 U1086 ( .A(n780), .B(n779), .C(n778), .CO(n777), .S(n827) );
  CMPR32X1 U1087 ( .A(n783), .B(n782), .C(n781), .CO(n795), .S(n826) );
  CMPR32X1 U1088 ( .A(n786), .B(n785), .C(n784), .CO(n781), .S(n840) );
  XNOR2XL U1089 ( .A(n331), .B(A[4]), .Y(n847) );
  OAI22XL U1090 ( .A0(n906), .A1(n847), .B0(n995), .B1(n787), .Y(n846) );
  OAI22XL U1091 ( .A0(n983), .A1(n823), .B0(n990), .B1(n788), .Y(n845) );
  ADDFHX1 U1092 ( .A(n792), .B(n791), .CI(n790), .CO(n808), .S(n838) );
  CMPR32X1 U1093 ( .A(n795), .B(n794), .C(n793), .CO(n773), .S(n803) );
  NOR2XL U1094 ( .A(n797), .B(n796), .Y(mult_x_1_n286) );
  OAI21XL U1095 ( .A0(n859), .A1(n799), .B0(n798), .Y(n802) );
  INVXL U1096 ( .A(n1337), .Y(n800) );
  NAND2XL U1097 ( .A(n800), .B(n1338), .Y(n801) );
  CMPR32X1 U1098 ( .A(n808), .B(n807), .C(n806), .CO(n793), .S(n837) );
  XNOR2XL U1099 ( .A(n922), .B(A[6]), .Y(n822) );
  OAI22XL U1100 ( .A0(n924), .A1(n822), .B0(n6), .B1(n809), .Y(n843) );
  OAI22XL U1101 ( .A0(n812), .A1(n811), .B0(n819), .B1(n810), .Y(n842) );
  XNOR2X1 U1102 ( .A(n867), .B(A[2]), .Y(n821) );
  CMPR32X1 U1103 ( .A(n816), .B(n815), .C(n814), .CO(n806), .S(n855) );
  XNOR2X1 U1104 ( .A(n922), .B(A[5]), .Y(n866) );
  OAI22XL U1105 ( .A0(n924), .A1(n866), .B0(n6), .B1(n822), .Y(n877) );
  NOR2XL U1106 ( .A(n829), .B(n828), .Y(mult_x_1_n292) );
  NAND2XL U1107 ( .A(n829), .B(n828), .Y(mult_x_1_n293) );
  INVXL U1108 ( .A(n1295), .Y(n831) );
  INVXL U1109 ( .A(n1296), .Y(n830) );
  OAI21XL U1110 ( .A0(n859), .A1(n831), .B0(n830), .Y(n834) );
  NAND2XL U1111 ( .A(n1340), .B(n832), .Y(n833) );
  XNOR2X1 U1112 ( .A(n834), .B(n833), .Y(PRODUCT[15]) );
  CMPR32X1 U1113 ( .A(n840), .B(n839), .C(n838), .CO(n825), .S(n862) );
  CMPR32X1 U1114 ( .A(n843), .B(n842), .C(n841), .CO(n856), .S(n880) );
  CMPR32X1 U1115 ( .A(n846), .B(n845), .C(n844), .CO(n839), .S(n879) );
  OAI22XL U1116 ( .A0(n1137), .A1(n850), .B0(n7), .B1(n849), .Y(n873) );
  CMPR32X1 U1117 ( .A(n853), .B(n852), .C(n851), .CO(n864), .S(n885) );
  CMPR32X1 U1118 ( .A(n856), .B(n855), .C(n854), .CO(n836), .S(n860) );
  NOR2XL U1119 ( .A(n858), .B(n857), .Y(mult_x_1_n299) );
  XOR2X1 U1120 ( .A(n859), .B(n1341), .Y(PRODUCT[14]) );
  XNOR2X1 U1121 ( .A(n8), .B(A[6]), .Y(n891) );
  ADDHXL U1122 ( .A(n874), .B(n873), .CO(n886), .S(n899) );
  CMPR32X1 U1123 ( .A(n877), .B(n876), .C(n875), .CO(n863), .S(n896) );
  INVXL U1124 ( .A(n881), .Y(mult_x_1_n304) );
  INVXL U1125 ( .A(n884), .Y(mult_x_1_n305) );
  NAND2XL U1126 ( .A(mult_x_1_n304), .B(n884), .Y(mult_x_1_n84) );
  OAI22XL U1127 ( .A0(n912), .A1(n910), .B0(n995), .B1(n889), .Y(n907) );
  XNOR2X1 U1128 ( .A(n922), .B(A[3]), .Y(n909) );
  OAI22XL U1129 ( .A0(n986), .A1(n913), .B0(n9), .B1(n891), .Y(n1025) );
  CMPR32X1 U1130 ( .A(n895), .B(n894), .C(n893), .CO(n898), .S(n914) );
  CMPR32X1 U1131 ( .A(n901), .B(n900), .C(n899), .CO(n897), .S(n1023) );
  OAI22X1 U1132 ( .A0(n764), .A1(n996), .B0(n902), .B1(n1128), .Y(n994) );
  OAI22X1 U1133 ( .A0(n906), .A1(n905), .B0(n904), .B1(n903), .Y(n993) );
  OAI22XL U1134 ( .A0(n986), .A1(n984), .B0(n9), .B1(n913), .Y(n978) );
  NOR2XL U1135 ( .A(n918), .B(n917), .Y(n1147) );
  INVXL U1136 ( .A(n1147), .Y(mult_x_1_n317) );
  OAI22X1 U1137 ( .A0(n942), .A1(n921), .B0(n997), .B1(n1128), .Y(n988) );
  NOR2BX1 U1138 ( .AN(A[0]), .B(n6), .Y(n932) );
  OAI22X2 U1139 ( .A0(n942), .A1(n927), .B0(n921), .B1(n1128), .Y(n931) );
  OAI22X1 U1140 ( .A0(n986), .A1(n937), .B0(n9), .B1(n925), .Y(n930) );
  XNOR2X1 U1141 ( .A(n922), .B(A[0]), .Y(n923) );
  OAI22XL U1142 ( .A0(n986), .A1(n925), .B0(n9), .B1(n985), .Y(n1004) );
  OAI22XL U1143 ( .A0(n986), .A1(n929), .B0(n9), .B1(n928), .Y(n939) );
  XNOR2X1 U1144 ( .A(n981), .B(A[2]), .Y(n956) );
  OAI22XL U1145 ( .A0(n986), .A1(n938), .B0(n9), .B1(n937), .Y(n965) );
  ADDHXL U1146 ( .A(n940), .B(n939), .CO(n934), .S(n964) );
  NOR2XL U1147 ( .A(n1232), .B(n1241), .Y(n977) );
  OR2X2 U1148 ( .A(n945), .B(n944), .Y(n1273) );
  OAI22X1 U1149 ( .A0(n942), .A1(n947), .B0(n955), .B1(n953), .Y(n959) );
  OAI22X1 U1150 ( .A0(n992), .A1(n948), .B0(n990), .B1(n957), .Y(n958) );
  OAI21XL U1151 ( .A0(n1270), .A1(n1267), .B0(n1268), .Y(n1265) );
  OAI22XL U1152 ( .A0(n983), .A1(n957), .B0(n990), .B1(n956), .Y(n967) );
  CMPR22X1 U1153 ( .A(n959), .B(n958), .CO(n961), .S(n952) );
  CMPR32X1 U1154 ( .A(n966), .B(n965), .C(n964), .CO(n972), .S(n971) );
  CMPR32X1 U1155 ( .A(n969), .B(n968), .C(n967), .CO(n970), .S(n962) );
  OAI21XL U1156 ( .A0(n1249), .A1(n1246), .B0(n1247), .Y(n1231) );
  NAND2XL U1157 ( .A(n975), .B(n974), .Y(n1233) );
  OAI21XL U1158 ( .A0(n1232), .A1(n1242), .B0(n1233), .Y(n976) );
  AOI21XL U1159 ( .A0(n977), .A1(n1231), .B0(n976), .Y(n1069) );
  CMPR22X1 U1160 ( .A(n994), .B(n993), .CO(n1032), .S(n1028) );
  CMPR32X1 U1161 ( .A(n1015), .B(n1014), .C(n1013), .CO(n1016), .S(n975) );
  OR2X2 U1162 ( .A(n1017), .B(n1016), .Y(n1209) );
  INVXL U1163 ( .A(n1208), .Y(n1070) );
  NAND2XL U1164 ( .A(n1019), .B(n1018), .Y(n1071) );
  INVXL U1165 ( .A(n1071), .Y(n1020) );
  CMPR32X1 U1166 ( .A(n1023), .B(n1022), .C(n1021), .CO(n917), .S(n1042) );
  CMPR32X1 U1167 ( .A(n1026), .B(n1025), .C(n1024), .CO(n915), .S(n1035) );
  CMPR32X1 U1168 ( .A(n1035), .B(n1034), .C(n1033), .CO(n1041), .S(n1040) );
  NOR2XL U1169 ( .A(n1058), .B(n1064), .Y(n1044) );
  OAI21XL U1170 ( .A0(n1058), .A1(n1065), .B0(n1059), .Y(n1043) );
  NAND2XL U1171 ( .A(n1056), .B(mult_x_1_n317), .Y(n1054) );
  OAI21XL U1172 ( .A0(n1063), .A1(n1054), .B0(n1053), .Y(mult_x_1_n309) );
  NAND2XL U1173 ( .A(n1056), .B(n1055), .Y(mult_x_1_n85) );
  XNOR2X1 U1174 ( .A(n1299), .B(n1343), .Y(PRODUCT[12]) );
  INVXL U1175 ( .A(n1058), .Y(n1060) );
  NAND2XL U1176 ( .A(n1060), .B(n1059), .Y(n1061) );
  INVXL U1177 ( .A(n1063), .Y(mult_x_1_n321) );
  INVXL U1178 ( .A(n1064), .Y(n1066) );
  NAND2XL U1179 ( .A(n1066), .B(n1065), .Y(n1067) );
  INVXL U1180 ( .A(n1069), .Y(n1211) );
  AOI21XL U1181 ( .A0(n1211), .A1(n1209), .B0(n1070), .Y(n1073) );
  ADDFHX1 U1182 ( .A(n1082), .B(n1081), .CI(n1080), .CO(n515), .S(
        mult_x_1_n554) );
  ADDFHX1 U1183 ( .A(n1088), .B(n1087), .CI(n1086), .CO(n508), .S(n1096) );
  CMPR32X1 U1184 ( .A(n1091), .B(n1089), .C(n1090), .CO(n1095), .S(n1092) );
  CMPR32X1 U1185 ( .A(n1109), .B(n1108), .C(n1107), .CO(n1118), .S(n1111) );
  ADDFHX1 U1186 ( .A(n1121), .B(n1120), .CI(n1119), .CO(mult_x_1_n601), .S(
        n630) );
  ADDFHX1 U1187 ( .A(n1124), .B(n1123), .CI(n1122), .CO(n629), .S(
        mult_x_1_n618) );
  ADDFHX1 U1188 ( .A(n1127), .B(n1126), .CI(n1125), .CO(mult_x_1_n633), .S(
        n704) );
  CMPR32X1 U1189 ( .A(n1133), .B(n1132), .C(n1131), .CO(n1150), .S(n1129) );
  CMPR32X1 U1190 ( .A(n1143), .B(n1142), .C(n1141), .CO(n1160), .S(n1133) );
  CMPR32X1 U1191 ( .A(n1146), .B(n1145), .C(n1144), .CO(n1151), .S(n1132) );
  NAND2XL U1192 ( .A(mult_x_1_n317), .B(n1148), .Y(mult_x_1_n86) );
  CMPR32X1 U1193 ( .A(n1153), .B(n1152), .C(n1151), .CO(n1164), .S(n1149) );
  CMPR32X1 U1194 ( .A(n1156), .B(n1155), .C(n1154), .CO(n1167), .S(n1153) );
  OAI22X1 U1195 ( .A0(n1176), .A1(n1159), .B0(n1177), .B1(n1174), .Y(n1188) );
  CMPR32X1 U1196 ( .A(n1162), .B(n1161), .C(n1160), .CO(n1165), .S(n1152) );
  CMPR32X1 U1197 ( .A(n1167), .B(n1166), .C(n1165), .CO(n1179), .S(n1163) );
  CMPR32X1 U1198 ( .A(n1172), .B(n1171), .C(n1170), .CO(n1181), .S(n1166) );
  CMPR32X1 U1199 ( .A(n1182), .B(n1181), .C(n1180), .CO(n1190), .S(n1178) );
  CMPR32X1 U1200 ( .A(n1188), .B(n1187), .C(n1186), .CO(n1191), .S(n1180) );
  CMPR32X1 U1201 ( .A(n1193), .B(n1192), .C(n1191), .CO(n1205), .S(n1189) );
  XOR3X2 U1202 ( .A(n1203), .B(n1202), .C(n1201), .Y(n1204) );
  OAI21XL U1203 ( .A0(n1217), .A1(n1314), .B0(n1216), .Y(n1287) );
  OAI21XL U1204 ( .A0(n1293), .A1(n1221), .B0(n1220), .Y(n1223) );
  XNOR2X1 U1205 ( .A(n1223), .B(n1222), .Y(PRODUCT[36]) );
  OAI21XL U1206 ( .A0(n1293), .A1(n1227), .B0(n1226), .Y(n1230) );
  OAI21XL U1207 ( .A0(n1244), .A1(n1241), .B0(n1242), .Y(n1236) );
  INVXL U1208 ( .A(n1232), .Y(n1234) );
  OAI21XL U1209 ( .A0(n1305), .A1(n1308), .B0(n1306), .Y(n1255) );
  OAI21XL U1210 ( .A0(n1293), .A1(n1238), .B0(n1237), .Y(n1240) );
  OAI21XL U1211 ( .A0(n1293), .A1(n1260), .B0(n1259), .Y(n1263) );
  OAI21XL U1212 ( .A0(n1284), .A1(n1301), .B0(n1302), .Y(n1285) );
  OAI21XL U1213 ( .A0(n1290), .A1(n1289), .B0(n1288), .Y(n1291) );
  OAI21XL U1214 ( .A0(n1293), .A1(n1283), .B0(n1292), .Y(n1294) );
  XNOR2XL U1215 ( .A(n1294), .B(n1300), .Y(PRODUCT[40]) );
endmodule


module FFT2048_DW02_mult_2_stage_J1_3 ( A, B, TC, CLK, PRODUCT );
  input [25:0] A;
  input [16:0] B;
  output [42:0] PRODUCT;
  input TC, CLK;
  wire   n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, mult_x_1_n665, mult_x_1_n650, mult_x_1_n649,
         mult_x_1_n634, mult_x_1_n633, mult_x_1_n618, mult_x_1_n617,
         mult_x_1_n602, mult_x_1_n601, mult_x_1_n586, mult_x_1_n585,
         mult_x_1_n570, mult_x_1_n569, mult_x_1_n554, mult_x_1_n553,
         mult_x_1_n538, mult_x_1_n537, mult_x_1_n522, mult_x_1_n521,
         mult_x_1_n508, mult_x_1_n507, mult_x_1_n494, mult_x_1_n493,
         mult_x_1_n482, mult_x_1_n481, mult_x_1_n470, mult_x_1_n322,
         mult_x_1_n318, mult_x_1_n311, mult_x_1_n310, mult_x_1_n305,
         mult_x_1_n298, mult_x_1_n293, mult_x_1_n292, mult_x_1_n287,
         mult_x_1_n286, mult_x_1_n282, mult_x_1_n281, mult_x_1_n177,
         mult_x_1_n176, mult_x_1_n170, mult_x_1_n169, mult_x_1_n161,
         mult_x_1_n160, mult_x_1_n152, mult_x_1_n151, mult_x_1_n137,
         mult_x_1_n136, mult_x_1_n130, mult_x_1_n129, mult_x_1_n121,
         mult_x_1_n120, mult_x_1_n110, mult_x_1_n109, mult_x_1_n86,
         mult_x_1_n85, mult_x_1_n84, mult_x_1_n83, mult_x_1_n58, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330;

  DFFHQXL mult_x_1_clk_r_REG8_S1 ( .D(mult_x_1_n493), .CK(CLK), .Q(n1307) );
  DFFHQXL mult_x_1_clk_r_REG11_S1 ( .D(mult_x_1_n482), .CK(CLK), .Q(n1306) );
  DFFHQXL mult_x_1_clk_r_REG12_S1 ( .D(mult_x_1_n470), .CK(CLK), .Q(n1304) );
  DFFHQXL mult_x_1_clk_r_REG10_S1 ( .D(mult_x_1_n481), .CK(CLK), .Q(n1305) );
  DFFHQXL mult_x_1_clk_r_REG16_S1 ( .D(mult_x_1_n169), .CK(CLK), .Q(n1287) );
  DFFHQX4 mult_x_1_clk_r_REG46_S1 ( .D(mult_x_1_n286), .CK(CLK), .Q(n1293) );
  DFFHQXL mult_x_1_clk_r_REG18_S1 ( .D(mult_x_1_n160), .CK(CLK), .Q(n1285) );
  DFFHQX4 mult_x_1_clk_r_REG42_S1 ( .D(mult_x_1_n665), .CK(CLK), .Q(n1329) );
  DFFHQX4 mult_x_1_clk_r_REG41_S1 ( .D(mult_x_1_n650), .CK(CLK), .Q(n1328) );
  DFFHQX4 mult_x_1_clk_r_REG40_S1 ( .D(mult_x_1_n649), .CK(CLK), .Q(n1327) );
  DFFHQX4 mult_x_1_clk_r_REG39_S1 ( .D(mult_x_1_n634), .CK(CLK), .Q(n1326) );
  DFFHQX4 mult_x_1_clk_r_REG37_S1 ( .D(mult_x_1_n618), .CK(CLK), .Q(n1324) );
  DFFHQX4 mult_x_1_clk_r_REG35_S1 ( .D(mult_x_1_n602), .CK(CLK), .Q(n1322) );
  DFFHQX4 mult_x_1_clk_r_REG34_S1 ( .D(mult_x_1_n601), .CK(CLK), .Q(n1321) );
  DFFHQX4 mult_x_1_clk_r_REG33_S1 ( .D(mult_x_1_n586), .CK(CLK), .Q(n1320) );
  DFFHQX4 mult_x_1_clk_r_REG7_S1 ( .D(mult_x_1_n508), .CK(CLK), .Q(n1310) );
  DFFHQX4 mult_x_1_clk_r_REG62_S1 ( .D(mult_x_1_n322), .CK(CLK), .Q(n1303) );
  DFFHQX4 mult_x_1_clk_r_REG57_S1 ( .D(mult_x_1_n310), .CK(CLK), .Q(n1299) );
  DFFHQX4 mult_x_1_clk_r_REG53_S1 ( .D(mult_x_1_n305), .CK(CLK), .Q(n1271) );
  DFFHQX4 mult_x_1_clk_r_REG54_S1 ( .D(n574), .CK(CLK), .Q(n1270) );
  DFFHQX4 mult_x_1_clk_r_REG51_S1 ( .D(n53), .CK(CLK), .Q(n1268) );
  DFFHQXL clk_r_REG61_S1 ( .D(n1343), .CK(CLK), .Q(PRODUCT[11]) );
  DFFHQXL mult_x_1_clk_r_REG13_S1 ( .D(mult_x_1_n177), .CK(CLK), .Q(n1290) );
  DFFHQXL mult_x_1_clk_r_REG19_S1 ( .D(mult_x_1_n152), .CK(CLK), .Q(n1284) );
  DFFHQXL mult_x_1_clk_r_REG55_S1 ( .D(mult_x_1_n85), .CK(CLK), .Q(n1300) );
  DFFHQXL mult_x_1_clk_r_REG14_S1 ( .D(mult_x_1_n176), .CK(CLK), .Q(n1289) );
  DFFHQXL mult_x_1_clk_r_REG17_S1 ( .D(mult_x_1_n161), .CK(CLK), .Q(n1286) );
  DFFHQXL mult_x_1_clk_r_REG52_S1 ( .D(mult_x_1_n84), .CK(CLK), .Q(n1298) );
  DFFHQXL clk_r_REG64_S1 ( .D(n1345), .CK(CLK), .Q(PRODUCT[9]) );
  DFFHQXL clk_r_REG63_S1 ( .D(n1344), .CK(CLK), .Q(PRODUCT[10]) );
  DFFHQXL mult_x_1_clk_r_REG49_S1 ( .D(mult_x_1_n83), .CK(CLK), .Q(n1297) );
  DFFHQXL clk_r_REG70_S1 ( .D(n1351), .CK(CLK), .Q(PRODUCT[3]) );
  DFFHQXL mult_x_1_clk_r_REG26_S1 ( .D(mult_x_1_n120), .CK(CLK), .Q(n1277) );
  DFFHQXL mult_x_1_clk_r_REG20_S1 ( .D(mult_x_1_n151), .CK(CLK), .Q(n1283) );
  DFFHQXL mult_x_1_clk_r_REG15_S1 ( .D(mult_x_1_n170), .CK(CLK), .Q(n1288) );
  DFFHQXL clk_r_REG65_S1 ( .D(n1346), .CK(CLK), .Q(PRODUCT[8]) );
  DFFHQXL clk_r_REG66_S1 ( .D(n1347), .CK(CLK), .Q(PRODUCT[7]) );
  DFFHQXL clk_r_REG67_S1 ( .D(n1348), .CK(CLK), .Q(PRODUCT[6]) );
  DFFHQXL clk_r_REG68_S1 ( .D(n1349), .CK(CLK), .Q(PRODUCT[5]) );
  DFFHQXL clk_r_REG69_S1 ( .D(n1350), .CK(CLK), .Q(PRODUCT[4]) );
  DFFHQXL clk_r_REG71_S1 ( .D(n1352), .CK(CLK), .Q(PRODUCT[2]) );
  DFFHQXL clk_r_REG72_S1 ( .D(n1353), .CK(CLK), .Q(PRODUCT[1]) );
  DFFHQXL clk_r_REG73_S1 ( .D(n1354), .CK(CLK), .Q(PRODUCT[0]) );
  DFFHQX1 mult_x_1_clk_r_REG2_S1 ( .D(mult_x_1_n537), .CK(CLK), .Q(n1313) );
  DFFHQXL mult_x_1_clk_r_REG6_S1 ( .D(mult_x_1_n507), .CK(CLK), .Q(n1309) );
  DFFHQXL mult_x_1_clk_r_REG58_S1 ( .D(mult_x_1_n86), .CK(CLK), .Q(n1301) );
  DFFHQX2 mult_x_1_clk_r_REG48_S1 ( .D(mult_x_1_n292), .CK(CLK), .Q(n1295) );
  DFFHQXL mult_x_1_clk_r_REG21_S1 ( .D(mult_x_1_n137), .CK(CLK), .Q(n1282) );
  DFFHQXL mult_x_1_clk_r_REG23_S1 ( .D(mult_x_1_n130), .CK(CLK), .Q(n1280) );
  DFFHQXL mult_x_1_clk_r_REG24_S1 ( .D(mult_x_1_n129), .CK(CLK), .Q(n1279) );
  DFFHQXL mult_x_1_clk_r_REG25_S1 ( .D(mult_x_1_n121), .CK(CLK), .Q(n1278) );
  DFFHQXL mult_x_1_clk_r_REG27_S1 ( .D(mult_x_1_n110), .CK(CLK), .Q(n1276) );
  DFFHQXL mult_x_1_clk_r_REG28_S1 ( .D(mult_x_1_n109), .CK(CLK), .Q(n1275) );
  DFFHQXL mult_x_1_clk_r_REG29_S1 ( .D(mult_x_1_n58), .CK(CLK), .Q(n1274) );
  DFFHQX1 mult_x_1_clk_r_REG59_S1 ( .D(mult_x_1_n318), .CK(CLK), .Q(n1273) );
  DFFHQX1 mult_x_1_clk_r_REG60_S1 ( .D(n1330), .CK(CLK), .Q(n1272) );
  DFFHQX1 mult_x_1_clk_r_REG43_S1 ( .D(mult_x_1_n282), .CK(CLK), .Q(n1292) );
  DFFHQXL mult_x_1_clk_r_REG9_S1 ( .D(mult_x_1_n494), .CK(CLK), .Q(n1308) );
  DFFHQXL mult_x_1_clk_r_REG22_S1 ( .D(mult_x_1_n136), .CK(CLK), .Q(n1281) );
  DFFHQX4 mult_x_1_clk_r_REG5_S1 ( .D(mult_x_1_n522), .CK(CLK), .Q(n1312) );
  DFFHQX4 mult_x_1_clk_r_REG45_S1 ( .D(mult_x_1_n287), .CK(CLK), .Q(n1294) );
  DFFHQX2 mult_x_1_clk_r_REG50_S1 ( .D(mult_x_1_n298), .CK(CLK), .Q(n1269) );
  DFFHQX1 mult_x_1_clk_r_REG56_S1 ( .D(mult_x_1_n311), .CK(CLK), .Q(n1302) );
  DFFHQX1 mult_x_1_clk_r_REG47_S1 ( .D(mult_x_1_n293), .CK(CLK), .Q(n1296) );
  DFFHQX2 mult_x_1_clk_r_REG44_S1 ( .D(mult_x_1_n281), .CK(CLK), .Q(n1291) );
  DFFHQX1 mult_x_1_clk_r_REG4_S1 ( .D(mult_x_1_n521), .CK(CLK), .Q(n1311) );
  DFFHQX1 mult_x_1_clk_r_REG30_S1 ( .D(mult_x_1_n569), .CK(CLK), .Q(n1317) );
  DFFHQX1 mult_x_1_clk_r_REG1_S1 ( .D(mult_x_1_n554), .CK(CLK), .Q(n1316) );
  DFFHQX2 mult_x_1_clk_r_REG0_S1 ( .D(mult_x_1_n553), .CK(CLK), .Q(n1315) );
  DFFHQX2 mult_x_1_clk_r_REG32_S1 ( .D(mult_x_1_n585), .CK(CLK), .Q(n1319) );
  DFFHQX2 mult_x_1_clk_r_REG3_S1 ( .D(mult_x_1_n538), .CK(CLK), .Q(n1314) );
  DFFHQX2 mult_x_1_clk_r_REG38_S1 ( .D(mult_x_1_n633), .CK(CLK), .Q(n1325) );
  DFFHQX2 mult_x_1_clk_r_REG36_S1 ( .D(mult_x_1_n617), .CK(CLK), .Q(n1323) );
  DFFHQX2 mult_x_1_clk_r_REG31_S1 ( .D(mult_x_1_n570), .CK(CLK), .Q(n1318) );
  ADDFHX1 U1 ( .A(n921), .B(n920), .CI(n919), .CO(mult_x_1_n569), .S(
        mult_x_1_n570) );
  ADDFHX1 U2 ( .A(n1082), .B(n1081), .CI(n1080), .CO(n1072), .S(n1083) );
  ADDFHX1 U3 ( .A(n918), .B(n917), .CI(n916), .CO(n886), .S(n919) );
  ADDFHX1 U4 ( .A(n1005), .B(n1004), .CI(n1003), .CO(n960), .S(n1006) );
  OAI21XL U5 ( .A0(n958), .A1(n15), .B0(n957), .Y(n11) );
  XOR2X1 U6 ( .A(n951), .B(n73), .Y(n1004) );
  XOR2X1 U7 ( .A(n876), .B(n67), .Y(n917) );
  ADDFHX1 U8 ( .A(n1064), .B(n1063), .CI(n1062), .CO(n1073), .S(n1081) );
  ADDFHX1 U9 ( .A(n881), .B(n880), .CI(n879), .CO(n884), .S(n916) );
  ADDFHX1 U10 ( .A(n1093), .B(n1092), .CI(n1091), .CO(n528), .S(n1098) );
  ADDFHX2 U11 ( .A(n1040), .B(n1039), .CI(n1038), .CO(n1049), .S(n1069) );
  ADDFHX1 U12 ( .A(n1002), .B(n1001), .CI(n1000), .CO(n1005), .S(n1044) );
  ADDFHX1 U13 ( .A(n915), .B(n914), .CI(n913), .CO(n918), .S(n957) );
  ADDFHX1 U14 ( .A(n1043), .B(n1042), .CI(n1041), .CO(n1046), .S(n1068) );
  ADDFX2 U15 ( .A(n1067), .B(n1066), .CI(n1065), .CO(n1070), .S(n1080) );
  ADDFHX1 U16 ( .A(n956), .B(n955), .CI(n954), .CO(n958), .S(n1003) );
  ADDFHX1 U17 ( .A(n446), .B(n445), .CI(n444), .CO(n1078), .S(n476) );
  ADDFX2 U18 ( .A(n770), .B(n769), .CI(n768), .CO(n138), .S(n786) );
  ADDFHX1 U19 ( .A(n1061), .B(n1060), .CI(n1059), .CO(n1082), .S(n1077) );
  ADDFHX1 U20 ( .A(n893), .B(n892), .CI(n891), .CO(n878), .S(n911) );
  ADDFHX1 U21 ( .A(n929), .B(n928), .CI(n927), .CO(n912), .S(n952) );
  ADDFHX1 U22 ( .A(n862), .B(n861), .CI(n860), .CO(n847), .S(n877) );
  CMPR32X1 U23 ( .A(n435), .B(n434), .C(n433), .CO(n1061), .S(n421) );
  OAI22X1 U24 ( .A0(n1163), .A1(n1013), .B0(n1014), .B1(n967), .Y(n1020) );
  OAI22X2 U25 ( .A0(n1163), .A1(n33), .B0(n1014), .B1(n1013), .Y(n1054) );
  ADDFHX1 U26 ( .A(n727), .B(n726), .CI(n725), .CO(n734), .S(n736) );
  XNOR2X1 U27 ( .A(n1161), .B(n966), .Y(n1013) );
  BUFX8 U28 ( .A(n1170), .Y(n1163) );
  CLKBUFX3 U29 ( .A(n984), .Y(n1116) );
  NAND2X4 U30 ( .A(n90), .B(n390), .Y(n1018) );
  INVX4 U31 ( .A(n395), .Y(n1161) );
  CLKINVX3 U32 ( .A(B[11]), .Y(n546) );
  CLKINVX3 U33 ( .A(B[15]), .Y(n395) );
  BUFX4 U34 ( .A(n1012), .Y(n965) );
  BUFX4 U35 ( .A(n595), .Y(n6) );
  NAND2X1 U36 ( .A(n96), .B(n595), .Y(n597) );
  BUFX4 U37 ( .A(B[9]), .Y(n972) );
  BUFX3 U38 ( .A(n411), .Y(n10) );
  INVX4 U39 ( .A(n653), .Y(n7) );
  BUFX3 U40 ( .A(n686), .Y(n990) );
  BUFX4 U41 ( .A(B[5]), .Y(n943) );
  BUFX3 U42 ( .A(B[1]), .Y(n648) );
  NAND2X1 U43 ( .A(n91), .B(n411), .Y(n686) );
  NAND2BXL U44 ( .AN(n315), .B(n317), .Y(n48) );
  XNOR2X1 U45 ( .A(n380), .B(n379), .Y(PRODUCT[20]) );
  OAI21XL U46 ( .A0(n533), .A1(n502), .B0(n501), .Y(n504) );
  AOI2BB1X1 U47 ( .A0N(n373), .A1N(n1293), .B0(n386), .Y(n18) );
  INVX4 U48 ( .A(n317), .Y(n1104) );
  AOI2BB1X2 U49 ( .A0N(n373), .A1N(n57), .B0(n374), .Y(n385) );
  NOR2X1 U50 ( .A(n1313), .B(n1312), .Y(n332) );
  NOR2X2 U51 ( .A(n376), .B(n381), .Y(n84) );
  NOR2X2 U52 ( .A(n1327), .B(n1326), .Y(n376) );
  NAND2X2 U53 ( .A(n1268), .B(n1270), .Y(n502) );
  NAND2X1 U54 ( .A(n1329), .B(n1328), .Y(n382) );
  NOR2X1 U55 ( .A(n1323), .B(n1322), .Y(n368) );
  NOR2X2 U56 ( .A(n1329), .B(n1328), .Y(n381) );
  XOR2XL U57 ( .A(n31), .B(n52), .Y(PRODUCT[24]) );
  XOR2XL U58 ( .A(n1104), .B(n1103), .Y(PRODUCT[21]) );
  XNOR2XL U59 ( .A(n648), .B(n966), .Y(n628) );
  XNOR2XL U60 ( .A(n963), .B(n642), .Y(n695) );
  XNOR2XL U61 ( .A(n938), .B(n650), .Y(n557) );
  XNOR2XL U62 ( .A(n648), .B(n962), .Y(n466) );
  XNOR2XL U63 ( .A(n938), .B(n980), .Y(n514) );
  XOR2XL U64 ( .A(n214), .B(n29), .Y(n28) );
  XOR2XL U65 ( .A(n938), .B(n27), .Y(n26) );
  XNOR2XL U66 ( .A(n648), .B(n933), .Y(n977) );
  XNOR2XL U67 ( .A(n938), .B(A[4]), .Y(n459) );
  XOR2XL U68 ( .A(n575), .B(n1300), .Y(PRODUCT[13]) );
  BUFX3 U69 ( .A(B[16]), .Y(n107) );
  XNOR2XL U70 ( .A(n1161), .B(A[7]), .Y(n924) );
  XNOR2XL U71 ( .A(n963), .B(A[12]), .Y(n1011) );
  XNOR2XL U72 ( .A(n7), .B(n942), .Y(n409) );
  XNOR2XL U73 ( .A(n972), .B(n1151), .Y(n249) );
  BUFX3 U74 ( .A(n392), .Y(n9) );
  BUFX3 U75 ( .A(n168), .Y(n8) );
  ADDFX2 U76 ( .A(n816), .B(n815), .CI(n814), .CO(n822), .S(n852) );
  NAND2BX1 U77 ( .AN(n470), .B(n39), .Y(n38) );
  ADDFX2 U78 ( .A(n244), .B(n243), .CI(n242), .CO(n223), .S(n283) );
  OAI21X2 U79 ( .A0(n58), .A1(n36), .B0(n35), .Y(n1048) );
  XOR2XL U80 ( .A(n23), .B(n823), .Y(mult_x_1_n522) );
  XNOR2XL U81 ( .A(n1209), .B(n1208), .Y(n1347) );
  XNOR2X1 U82 ( .A(n1189), .B(n1188), .Y(n1346) );
  NAND2XL U83 ( .A(n22), .B(n21), .Y(mult_x_1_n521) );
  NAND2XL U84 ( .A(n824), .B(n825), .Y(n21) );
  OAI21XL U85 ( .A0(n824), .A1(n825), .B0(n823), .Y(n22) );
  ADDFHX1 U86 ( .A(n1008), .B(n1007), .CI(n1006), .CO(mult_x_1_n601), .S(
        mult_x_1_n602) );
  ADDFHX2 U87 ( .A(n853), .B(n852), .CI(n851), .CO(n824), .S(n854) );
  ADDFHX1 U88 ( .A(n884), .B(n883), .CI(n882), .CO(n855), .S(n885) );
  XOR2X1 U89 ( .A(n1044), .B(n1046), .Y(n85) );
  OAI2BB1XL U90 ( .A0N(n66), .A1N(n876), .B0(n65), .Y(n887) );
  INVX1 U91 ( .A(n15), .Y(n12) );
  OAI2BB1XL U92 ( .A0N(n69), .A1N(n845), .B0(n68), .Y(n856) );
  OAI2BB1XL U93 ( .A0N(n72), .A1N(n951), .B0(n71), .Y(n961) );
  OR2XL U94 ( .A(n911), .B(n912), .Y(n75) );
  OAI2BB1XL U95 ( .A0N(n173), .A1N(n965), .B0(n172), .Y(n219) );
  OAI22XL U96 ( .A0(n1024), .A1(n114), .B0(n6), .B1(n250), .Y(n291) );
  OAI22X1 U97 ( .A0(n965), .A1(n522), .B0(n1010), .B1(n511), .Y(n539) );
  NOR2X1 U98 ( .A(n8), .B(n391), .Y(n442) );
  NOR2X1 U99 ( .A(n8), .B(n1137), .Y(n1149) );
  NOR2X1 U100 ( .A(n8), .B(n898), .Y(n931) );
  OAI22XL U101 ( .A0(n990), .A1(n807), .B0(n10), .B1(n777), .Y(n808) );
  INVX1 U102 ( .A(n9), .Y(n25) );
  INVX4 U103 ( .A(n623), .Y(n963) );
  BUFX3 U104 ( .A(n984), .Y(n5) );
  NAND2XL U105 ( .A(n32), .B(n355), .Y(n31) );
  NAND2X1 U106 ( .A(n383), .B(n382), .Y(n384) );
  AND2X2 U107 ( .A(n311), .B(n310), .Y(n51) );
  NAND2X1 U108 ( .A(n1102), .B(n1101), .Y(n1103) );
  NAND2X1 U109 ( .A(n360), .B(n146), .Y(n315) );
  AND2XL U110 ( .A(n280), .B(n1290), .Y(n281) );
  INVXL U111 ( .A(n942), .Y(n29) );
  INVXL U112 ( .A(n962), .Y(n27) );
  INVX1 U113 ( .A(n500), .Y(n533) );
  INVX1 U114 ( .A(n1303), .Y(n621) );
  NAND2X1 U115 ( .A(n1316), .B(n1317), .Y(n349) );
  XOR2X1 U116 ( .A(n824), .B(n825), .Y(n23) );
  ADDFHX1 U117 ( .A(n856), .B(n855), .CI(n854), .CO(mult_x_1_n537), .S(
        mult_x_1_n538) );
  NAND2X1 U118 ( .A(n1098), .B(n1097), .Y(n1099) );
  NAND2X1 U119 ( .A(n615), .B(n614), .Y(n1126) );
  ADDFHX1 U120 ( .A(n961), .B(n960), .CI(n959), .CO(mult_x_1_n585), .S(
        mult_x_1_n586) );
  ADDFHX1 U121 ( .A(n822), .B(n821), .CI(n820), .CO(n800), .S(n823) );
  ADDFHX1 U122 ( .A(n887), .B(n886), .CI(n885), .CO(mult_x_1_n553), .S(
        mult_x_1_n554) );
  NAND2X1 U123 ( .A(n732), .B(n731), .Y(n1199) );
  ADDFHX1 U124 ( .A(n1096), .B(n1095), .CI(n1094), .CO(n1097), .S(n571) );
  NOR2X1 U125 ( .A(n675), .B(n674), .Y(n1214) );
  NAND2X1 U126 ( .A(n675), .B(n674), .Y(n1215) );
  ADDFHX1 U127 ( .A(n613), .B(n612), .CI(n611), .CO(n616), .S(n615) );
  INVX1 U128 ( .A(n958), .Y(n13) );
  OAI2BB1X1 U129 ( .A0N(n75), .A1N(n910), .B0(n74), .Y(n921) );
  XNOR2X1 U130 ( .A(n958), .B(n15), .Y(n14) );
  ADDFHX1 U131 ( .A(n294), .B(n293), .CI(n292), .CO(n756), .S(n759) );
  OR2XL U132 ( .A(n952), .B(n953), .Y(n72) );
  OR2XL U133 ( .A(n877), .B(n878), .Y(n66) );
  ADDFHX1 U134 ( .A(n536), .B(n535), .CI(n534), .CO(n525), .S(n1096) );
  ADDFHX1 U135 ( .A(n971), .B(n970), .CI(n969), .CO(n953), .S(n998) );
  ADDFHX1 U136 ( .A(n831), .B(n830), .CI(n829), .CO(n819), .S(n846) );
  OAI22X1 U137 ( .A0(n5), .A1(n900), .B0(n9), .B1(n16), .Y(n906) );
  OAI22X1 U138 ( .A0(n5), .A1(n16), .B0(n9), .B1(n26), .Y(n872) );
  NOR2X1 U139 ( .A(n8), .B(n836), .Y(n864) );
  NOR2BX1 U140 ( .AN(n1090), .B(n1016), .Y(n549) );
  XNOR2XL U141 ( .A(n1161), .B(A[25]), .Y(n1168) );
  XNOR2XL U142 ( .A(n1161), .B(A[24]), .Y(n1162) );
  NOR2X1 U143 ( .A(n8), .B(n108), .Y(n769) );
  NOR2X1 U144 ( .A(n8), .B(n936), .Y(n974) );
  NOR2X1 U145 ( .A(n8), .B(n441), .Y(n1027) );
  NOR2BX1 U146 ( .AN(n1090), .B(n9), .Y(n600) );
  XNOR2X1 U147 ( .A(n1213), .B(n1212), .Y(PRODUCT[38]) );
  XNOR2X1 U148 ( .A(n1196), .B(n1195), .Y(PRODUCT[37]) );
  XNOR2X1 U149 ( .A(n167), .B(n166), .Y(PRODUCT[36]) );
  XNOR2X1 U150 ( .A(n1231), .B(n1230), .Y(PRODUCT[39]) );
  NOR2X1 U151 ( .A(n1255), .B(n163), .Y(n1220) );
  XNOR2X1 U152 ( .A(n504), .B(n503), .Y(PRODUCT[16]) );
  AOI21X1 U153 ( .A0(n1272), .A1(n621), .B0(n1273), .Y(n575) );
  INVXL U154 ( .A(n375), .Y(n57) );
  BUFX2 U155 ( .A(A[5]), .Y(n966) );
  BUFX2 U156 ( .A(A[9]), .Y(n937) );
  BUFX2 U157 ( .A(A[8]), .Y(n925) );
  BUFX2 U158 ( .A(A[22]), .Y(n1151) );
  BUFX2 U159 ( .A(A[16]), .Y(n902) );
  BUFX2 U160 ( .A(A[17]), .Y(n940) );
  BUFX2 U161 ( .A(A[20]), .Y(n1112) );
  INVX1 U162 ( .A(n1285), .Y(n206) );
  INVX1 U163 ( .A(n1294), .Y(n386) );
  NAND2X1 U164 ( .A(n1326), .B(n1327), .Y(n377) );
  NAND2XL U165 ( .A(n232), .B(n231), .Y(mult_x_1_n161) );
  ADDFHX1 U166 ( .A(n144), .B(n143), .CI(n142), .CO(mult_x_1_n493), .S(
        mult_x_1_n494) );
  ADDFHX2 U167 ( .A(n1073), .B(n1072), .CI(n1071), .CO(mult_x_1_n633), .S(
        mult_x_1_n634) );
  ADDFHX2 U168 ( .A(n1049), .B(n1048), .CI(n1047), .CO(mult_x_1_n617), .S(
        mult_x_1_n618) );
  INVXL U169 ( .A(n1198), .Y(n77) );
  OR2XL U170 ( .A(n1175), .B(n1174), .Y(n1177) );
  OR2X2 U171 ( .A(n715), .B(n714), .Y(n747) );
  ADDFHX1 U172 ( .A(n730), .B(n729), .CI(n728), .CO(n731), .S(n715) );
  INVXL U173 ( .A(n1077), .Y(n89) );
  NAND2XL U174 ( .A(n61), .B(n60), .Y(n804) );
  ADDFHX2 U175 ( .A(n850), .B(n849), .CI(n848), .CO(n853), .S(n882) );
  NAND2XL U176 ( .A(n846), .B(n847), .Y(n68) );
  OR2XL U177 ( .A(n846), .B(n847), .Y(n69) );
  ADDFHX1 U178 ( .A(n291), .B(n290), .CI(n289), .CO(n757), .S(n761) );
  NAND2XL U179 ( .A(n877), .B(n878), .Y(n65) );
  NAND2XL U180 ( .A(n952), .B(n953), .Y(n71) );
  NAND2XL U181 ( .A(n911), .B(n912), .Y(n74) );
  ADDFHX1 U182 ( .A(n415), .B(n414), .CI(n413), .CO(n422), .S(n478) );
  ADDFHX1 U183 ( .A(n113), .B(n112), .CI(n111), .CO(n289), .S(n137) );
  ADDFHX1 U184 ( .A(n702), .B(n701), .CI(n700), .CO(n707), .S(n709) );
  OAI21XL U185 ( .A0(n1116), .A1(n26), .B0(n24), .Y(n841) );
  ADDFHX1 U186 ( .A(n463), .B(n462), .CI(n461), .CO(n455), .S(n509) );
  NAND2BX1 U187 ( .AN(n805), .B(n25), .Y(n24) );
  OR2X2 U188 ( .A(n664), .B(n663), .Y(n662) );
  OAI2BB1XL U189 ( .A0N(n6), .A1N(n597), .B0(n176), .Y(n193) );
  AND2XL U190 ( .A(n1252), .B(n1251), .Y(n1353) );
  OR2XL U191 ( .A(n646), .B(n645), .Y(n1246) );
  XNOR2XL U192 ( .A(n107), .B(A[24]), .Y(n1167) );
  XNOR2XL U193 ( .A(n107), .B(n1159), .Y(n1160) );
  OR2XL U194 ( .A(n1250), .B(n1249), .Y(n1252) );
  XNOR2XL U195 ( .A(n107), .B(n902), .Y(n170) );
  OAI2BB1XL U196 ( .A0N(n1089), .A1N(n935), .B0(n129), .Y(n778) );
  XOR2X2 U197 ( .A(B[7]), .B(n49), .Y(n595) );
  XOR2X1 U198 ( .A(n47), .B(n308), .Y(PRODUCT[31]) );
  XNOR2X1 U199 ( .A(n235), .B(n234), .Y(PRODUCT[33]) );
  XOR2X1 U200 ( .A(B[3]), .B(B[2]), .Y(n42) );
  AND2X1 U201 ( .A(n359), .B(n358), .Y(n52) );
  NAND2X1 U202 ( .A(n84), .B(n375), .Y(n83) );
  AND2X2 U203 ( .A(n307), .B(n306), .Y(n308) );
  NAND2XL U204 ( .A(n1296), .B(n30), .Y(n503) );
  INVX1 U205 ( .A(A[12]), .Y(n17) );
  BUFX2 U206 ( .A(A[10]), .Y(n899) );
  BUFX2 U207 ( .A(A[13]), .Y(n962) );
  BUFX2 U208 ( .A(A[21]), .Y(n1136) );
  BUFX2 U209 ( .A(A[14]), .Y(n922) );
  BUFX2 U210 ( .A(A[15]), .Y(n942) );
  BUFX2 U211 ( .A(A[23]), .Y(n1159) );
  BUFX2 U212 ( .A(A[19]), .Y(n933) );
  OAI21XL U213 ( .A0(n1078), .A1(n1079), .B0(n1077), .Y(n88) );
  XNOR2X1 U214 ( .A(n1161), .B(n980), .Y(n393) );
  XNOR2X1 U215 ( .A(n367), .B(n366), .Y(PRODUCT[23]) );
  XNOR2X1 U216 ( .A(n1117), .B(n933), .Y(n210) );
  AOI21X2 U217 ( .A0(n84), .A1(n374), .B0(n81), .Y(n82) );
  OAI21XL U218 ( .A0(n1266), .A1(n279), .B0(n278), .Y(n282) );
  XOR2X1 U219 ( .A(n59), .B(n1070), .Y(n1071) );
  OAI21X2 U220 ( .A0(n13), .A1(n12), .B0(n11), .Y(n920) );
  XNOR2X1 U221 ( .A(n14), .B(n957), .Y(n959) );
  XOR3X2 U222 ( .A(n912), .B(n911), .C(n910), .Y(n15) );
  XOR2X1 U223 ( .A(n938), .B(n17), .Y(n16) );
  XOR2X2 U224 ( .A(n18), .B(n388), .Y(PRODUCT[18]) );
  AOI21X4 U225 ( .A0(n20), .A1(n500), .B0(n19), .Y(n373) );
  OAI21X4 U226 ( .A0(n501), .A1(n1295), .B0(n1296), .Y(n19) );
  OAI21X2 U227 ( .A0(n1299), .A1(n1303), .B0(n1302), .Y(n500) );
  NOR2X4 U228 ( .A(n1295), .B(n502), .Y(n20) );
  OAI22X1 U229 ( .A0(n1116), .A1(n805), .B0(n9), .B1(n28), .Y(n810) );
  OAI21XL U230 ( .A0(n1116), .A1(n28), .B0(n63), .Y(n62) );
  INVX1 U231 ( .A(n1295), .Y(n30) );
  NAND2BX1 U232 ( .AN(n356), .B(n317), .Y(n32) );
  OAI21X4 U233 ( .A0(n83), .A1(n373), .B0(n82), .Y(n317) );
  OAI21X1 U234 ( .A0(n385), .A1(n381), .B0(n382), .Y(n380) );
  AOI21X4 U235 ( .A0(n1271), .A1(n1268), .B0(n1269), .Y(n501) );
  XOR2X1 U236 ( .A(B[10]), .B(B[11]), .Y(n97) );
  OAI22X1 U237 ( .A0(n393), .A1(n1163), .B0(n1014), .B1(n33), .Y(n1030) );
  XOR2X1 U238 ( .A(n1161), .B(n34), .Y(n33) );
  INVX1 U239 ( .A(A[4]), .Y(n34) );
  OAI21X1 U240 ( .A0(n1070), .A1(n1069), .B0(n1068), .Y(n35) );
  INVX1 U241 ( .A(n1070), .Y(n36) );
  NAND2X1 U242 ( .A(n472), .B(n473), .Y(mult_x_1_n282) );
  OAI2BB1X1 U243 ( .A0N(n38), .A1N(n469), .B0(n37), .Y(n1087) );
  NAND2XL U244 ( .A(n470), .B(n471), .Y(n37) );
  INVX1 U245 ( .A(n471), .Y(n39) );
  XOR3X2 U246 ( .A(n471), .B(n470), .C(n469), .Y(n474) );
  XOR2X2 U247 ( .A(n40), .B(n51), .Y(PRODUCT[30]) );
  OAI21X1 U248 ( .A0(n1266), .A1(n312), .B0(n313), .Y(n40) );
  AOI2BB1X4 U249 ( .A0N(n48), .A1N(n150), .B0(n41), .Y(n1266) );
  OAI21X1 U250 ( .A0(n150), .A1(n348), .B0(n149), .Y(n41) );
  NAND2X2 U251 ( .A(n42), .B(n93), .Y(n987) );
  XNOR2X2 U252 ( .A(B[2]), .B(B[1]), .Y(n93) );
  OAI21XL U253 ( .A0(n1163), .A1(n45), .B0(n43), .Y(n774) );
  NAND2BX1 U254 ( .AN(n110), .B(n44), .Y(n43) );
  INVX1 U255 ( .A(n1014), .Y(n44) );
  OAI22X1 U256 ( .A0(n827), .A1(n1163), .B0(n1014), .B1(n45), .Y(n830) );
  XOR2X1 U257 ( .A(n1161), .B(n46), .Y(n45) );
  INVX1 U258 ( .A(A[11]), .Y(n46) );
  NOR2X1 U259 ( .A(n332), .B(n323), .Y(n148) );
  OAI21XL U260 ( .A0(n1266), .A1(n305), .B0(n304), .Y(n47) );
  OAI21X2 U261 ( .A0(n368), .A1(n1101), .B0(n369), .Y(n361) );
  NAND2X1 U262 ( .A(n1325), .B(n1324), .Y(n1101) );
  XOR2X1 U263 ( .A(n282), .B(n281), .Y(PRODUCT[32]) );
  INVX1 U264 ( .A(B[8]), .Y(n49) );
  XNOR2X1 U265 ( .A(n972), .B(n925), .Y(n404) );
  XOR2X1 U266 ( .A(B[8]), .B(B[9]), .Y(n96) );
  NOR2X1 U267 ( .A(n473), .B(n472), .Y(mult_x_1_n281) );
  XNOR2X1 U268 ( .A(n1161), .B(n642), .Y(n398) );
  XNOR2X1 U269 ( .A(n1161), .B(n650), .Y(n399) );
  XNOR2X2 U270 ( .A(B[14]), .B(B[13]), .Y(n104) );
  XNOR2X2 U271 ( .A(B[10]), .B(B[9]), .Y(n392) );
  XNOR2X1 U272 ( .A(n963), .B(A[4]), .Y(n581) );
  XNOR2X1 U273 ( .A(n963), .B(n933), .Y(n788) );
  XNOR2X1 U274 ( .A(n963), .B(n980), .Y(n601) );
  XNOR2X1 U275 ( .A(n963), .B(n650), .Y(n696) );
  XNOR2X1 U276 ( .A(n963), .B(A[18]), .Y(n826) );
  XNOR2X1 U277 ( .A(n963), .B(n922), .Y(n964) );
  XNOR2X1 U278 ( .A(n7), .B(A[24]), .Y(n128) );
  NOR2X1 U279 ( .A(n8), .B(n773), .Y(n781) );
  XNOR2X1 U280 ( .A(n107), .B(n937), .Y(n773) );
  XNOR2X1 U281 ( .A(n648), .B(A[25]), .Y(n772) );
  XNOR2X1 U282 ( .A(n648), .B(n902), .Y(n396) );
  XNOR2X1 U283 ( .A(n648), .B(n899), .Y(n579) );
  XNOR2X1 U284 ( .A(n648), .B(n942), .Y(n397) );
  XNOR2X1 U285 ( .A(n648), .B(n937), .Y(n593) );
  XOR2X1 U286 ( .A(B[14]), .B(B[15]), .Y(n99) );
  XNOR2X1 U287 ( .A(n938), .B(n922), .Y(n805) );
  XNOR2X1 U288 ( .A(n64), .B(n62), .Y(n815) );
  INVXL U289 ( .A(n1259), .Y(n162) );
  XOR2XL U290 ( .A(B[6]), .B(B[7]), .Y(n98) );
  CLKBUFX8 U291 ( .A(n597), .Y(n1024) );
  INVXL U292 ( .A(n1254), .Y(n163) );
  XNOR2XL U293 ( .A(n943), .B(n925), .Y(n524) );
  XNOR2X1 U294 ( .A(n1117), .B(n650), .Y(n512) );
  XNOR2XL U295 ( .A(n7), .B(A[25]), .Y(n94) );
  XNOR2XL U296 ( .A(n943), .B(A[24]), .Y(n123) );
  XNOR2X1 U297 ( .A(n1117), .B(n902), .Y(n121) );
  BUFX3 U298 ( .A(A[2]), .Y(n642) );
  BUFX3 U299 ( .A(A[3]), .Y(n980) );
  OAI21XL U300 ( .A0(n1289), .A1(n306), .B0(n1290), .Y(n151) );
  INVXL U301 ( .A(n1277), .Y(n1222) );
  INVXL U302 ( .A(n1253), .Y(n1225) );
  NAND2XL U303 ( .A(n1194), .B(n1280), .Y(n1195) );
  NAND2XL U304 ( .A(n387), .B(n1292), .Y(n388) );
  XNOR2XL U305 ( .A(n943), .B(n922), .Y(n989) );
  XNOR2XL U306 ( .A(n943), .B(n962), .Y(n437) );
  XNOR2XL U307 ( .A(n943), .B(A[11]), .Y(n447) );
  NAND2X2 U308 ( .A(n97), .B(n392), .Y(n984) );
  OAI22XL U309 ( .A0(n979), .A1(n396), .B0(n440), .B1(n1089), .Y(n443) );
  NAND2BXL U310 ( .AN(n1090), .B(n107), .Y(n391) );
  XNOR2XL U311 ( .A(n943), .B(A[25]), .Y(n237) );
  OAI22X1 U312 ( .A0(n990), .A1(n123), .B0(n10), .B1(n237), .Y(n262) );
  XNOR2X1 U313 ( .A(n1117), .B(n940), .Y(n254) );
  XNOR2XL U314 ( .A(n943), .B(n1159), .Y(n103) );
  XNOR2XL U315 ( .A(n943), .B(n1151), .Y(n765) );
  OAI22XL U316 ( .A0(n965), .A1(n788), .B0(n1010), .B1(n106), .Y(n775) );
  BUFX3 U317 ( .A(A[1]), .Y(n650) );
  XNOR2XL U318 ( .A(n7), .B(n642), .Y(n658) );
  XNOR2XL U319 ( .A(n943), .B(n650), .Y(n638) );
  NOR2XL U320 ( .A(n8), .B(n1152), .Y(n1165) );
  INVXL U321 ( .A(n1153), .Y(n1154) );
  OAI22XL U322 ( .A0(n979), .A1(n897), .B0(n866), .B1(n976), .Y(n896) );
  CMPR32X1 U323 ( .A(n993), .B(n992), .C(n991), .CO(n1002), .S(n1042) );
  OAI22XL U324 ( .A0(n990), .A1(n988), .B0(n10), .B1(n944), .Y(n991) );
  OAI22XL U325 ( .A0(n56), .A1(n985), .B0(n93), .B1(n941), .Y(n992) );
  OAI22XL U326 ( .A0(n5), .A1(n982), .B0(n9), .B1(n939), .Y(n993) );
  OAI22XL U327 ( .A0(n1163), .A1(n1162), .B0(n1014), .B1(n1168), .Y(n1173) );
  OAI22X2 U328 ( .A0(n1163), .A1(n924), .B0(n1014), .B1(n889), .Y(n928) );
  OAI22XL U329 ( .A0(n1024), .A1(n973), .B0(n6), .B1(n930), .Y(n950) );
  NOR2XL U330 ( .A(n1304), .B(n1305), .Y(n275) );
  NOR2X1 U331 ( .A(n1307), .B(n1306), .Y(n309) );
  INVXL U332 ( .A(n1286), .Y(n159) );
  NAND2XL U333 ( .A(n206), .B(n158), .Y(n161) );
  NOR2XL U334 ( .A(n1281), .B(n1279), .Y(n1219) );
  INVXL U335 ( .A(n1281), .Y(n1191) );
  INVXL U336 ( .A(n1283), .Y(n158) );
  INVXL U337 ( .A(n1287), .Y(n233) );
  INVXL U338 ( .A(n332), .Y(n334) );
  INVXL U339 ( .A(n337), .Y(n350) );
  NAND2BXL U340 ( .AN(n1090), .B(n972), .Y(n594) );
  XNOR2XL U341 ( .A(n7), .B(n937), .Y(n559) );
  XNOR2X1 U342 ( .A(n963), .B(A[6]), .Y(n522) );
  XNOR2XL U343 ( .A(n943), .B(n899), .Y(n464) );
  NAND2BXL U344 ( .AN(n1090), .B(n943), .Y(n629) );
  XNOR2XL U345 ( .A(n963), .B(n1090), .Y(n625) );
  XNOR2XL U346 ( .A(n7), .B(n966), .Y(n683) );
  XNOR2XL U347 ( .A(n943), .B(n642), .Y(n626) );
  XNOR2XL U348 ( .A(n943), .B(n980), .Y(n685) );
  NOR2XL U349 ( .A(n275), .B(n1289), .Y(n152) );
  NOR2XL U350 ( .A(n161), .B(n1287), .Y(n1254) );
  NOR2XL U351 ( .A(n1253), .B(n1275), .Y(n1258) );
  NAND2XL U352 ( .A(n1220), .B(n1219), .Y(n1211) );
  OAI21XL U353 ( .A0(n533), .A1(n531), .B0(n530), .Y(n532) );
  INVXL U354 ( .A(n1271), .Y(n530) );
  XOR2X1 U355 ( .A(n533), .B(n1298), .Y(PRODUCT[14]) );
  OAI22XL U356 ( .A0(n990), .A1(n524), .B0(n10), .B1(n491), .Y(n540) );
  OAI22XL U357 ( .A0(n56), .A1(n523), .B0(n93), .B1(n490), .Y(n541) );
  XNOR2XL U358 ( .A(n943), .B(A[7]), .Y(n560) );
  CMPR32X1 U359 ( .A(n549), .B(n548), .C(n547), .CO(n554), .S(n576) );
  OAI22XL U360 ( .A0(n979), .A1(n544), .B0(n520), .B1(n1089), .Y(n548) );
  OAI22XL U361 ( .A0(n984), .A1(n557), .B0(n9), .B1(n521), .Y(n547) );
  NAND2BXL U362 ( .AN(n1090), .B(n938), .Y(n545) );
  INVXL U363 ( .A(n1114), .Y(n1115) );
  CMPR32X1 U364 ( .A(n517), .B(n516), .C(n515), .CO(n508), .S(n551) );
  OAI22XL U365 ( .A0(n990), .A1(n491), .B0(n10), .B1(n464), .Y(n517) );
  OAI22X1 U366 ( .A0(n965), .A1(n511), .B0(n1010), .B1(n465), .Y(n516) );
  OAI22XL U367 ( .A0(n56), .A1(n490), .B0(n93), .B1(n460), .Y(n492) );
  OAI22XL U368 ( .A0(n1024), .A1(n489), .B0(n6), .B1(n458), .Y(n494) );
  OAI22XL U369 ( .A0(n56), .A1(n690), .B0(n93), .B1(n689), .Y(n724) );
  XNOR2XL U370 ( .A(n943), .B(n1136), .Y(n777) );
  OAI22XL U371 ( .A0(n1024), .A1(n832), .B0(n6), .B1(n780), .Y(n813) );
  NAND2BXL U372 ( .AN(n1090), .B(n1161), .Y(n394) );
  OAI22XL U373 ( .A0(n935), .A1(n450), .B0(n397), .B1(n1089), .Y(n448) );
  OAI22X1 U374 ( .A0(n1163), .A1(n400), .B0(n1014), .B1(n399), .Y(n462) );
  NOR2XL U375 ( .A(n8), .B(n174), .Y(n195) );
  INVXL U376 ( .A(n175), .Y(n176) );
  OAI22XL U377 ( .A0(n1116), .A1(n179), .B0(n9), .B1(n191), .Y(n196) );
  OAI22XL U378 ( .A0(n1163), .A1(n177), .B0(n1014), .B1(n189), .Y(n198) );
  INVXL U379 ( .A(n485), .Y(n454) );
  OAI22XL U380 ( .A0(n965), .A1(n465), .B0(n1010), .B1(n420), .Y(n480) );
  OAI22XL U381 ( .A0(n56), .A1(n460), .B0(n93), .B1(n412), .Y(n482) );
  OAI22XL U382 ( .A0(n979), .A1(n466), .B0(n450), .B1(n1089), .Y(n487) );
  OAI22XL U383 ( .A0(n1018), .A1(n512), .B0(n1016), .B1(n451), .Y(n486) );
  NOR2BX1 U384 ( .AN(n1090), .B(n1014), .Y(n488) );
  NOR2XL U385 ( .A(n8), .B(n170), .Y(n221) );
  XNOR2XL U386 ( .A(n1161), .B(n940), .Y(n213) );
  CMPR32X1 U387 ( .A(n257), .B(n256), .C(n255), .CO(n286), .S(n293) );
  INVXL U388 ( .A(n262), .Y(n255) );
  NOR2XL U389 ( .A(n8), .B(n122), .Y(n256) );
  XNOR2XL U390 ( .A(n7), .B(n650), .Y(n659) );
  XNOR2XL U391 ( .A(n7), .B(A[4]), .Y(n627) );
  NAND2XL U392 ( .A(n1254), .B(n1258), .Y(n1261) );
  INVXL U393 ( .A(n1256), .Y(n1224) );
  NAND2XL U394 ( .A(n1220), .B(n1225), .Y(n1228) );
  INVXL U395 ( .A(n1275), .Y(n1229) );
  ADDFX2 U396 ( .A(n569), .B(n568), .CI(n567), .CO(n1095), .S(n608) );
  INVXL U397 ( .A(n1166), .Y(n1148) );
  OAI22XL U398 ( .A0(n1163), .A1(n1135), .B0(n1014), .B1(n1147), .Y(n1150) );
  NOR2XL U399 ( .A(n8), .B(n190), .Y(n1121) );
  OAI22XL U400 ( .A0(n1163), .A1(n189), .B0(n1014), .B1(n1119), .Y(n1122) );
  INVXL U401 ( .A(n1133), .Y(n1120) );
  INVXL U402 ( .A(n772), .Y(n129) );
  OR2X2 U403 ( .A(n9), .B(n127), .Y(n63) );
  CMPR32X1 U404 ( .A(n1021), .B(n1020), .C(n1019), .CO(n999), .S(n1039) );
  OAI22XL U405 ( .A0(n965), .A1(n1009), .B0(n1010), .B1(n964), .Y(n1021) );
  OAI22XL U406 ( .A0(n1024), .A1(n1023), .B0(n6), .B1(n1022), .Y(n1037) );
  OAI22XL U407 ( .A0(n990), .A1(n989), .B0(n10), .B1(n988), .Y(n1032) );
  OAI22XL U408 ( .A0(n56), .A1(n986), .B0(n93), .B1(n985), .Y(n1033) );
  OAI22XL U409 ( .A0(n1024), .A1(n1022), .B0(n6), .B1(n973), .Y(n996) );
  CMPR32X1 U410 ( .A(n1055), .B(n1054), .C(n1053), .CO(n1040), .S(n1063) );
  OAI22XL U411 ( .A0(n1012), .A1(n1011), .B0(n1010), .B1(n1009), .Y(n1055) );
  OAI22XL U412 ( .A0(n990), .A1(n416), .B0(n10), .B1(n437), .Y(n433) );
  OAI22XL U413 ( .A0(n965), .A1(n420), .B0(n1010), .B1(n419), .Y(n424) );
  OAI22XL U414 ( .A0(n990), .A1(n447), .B0(n10), .B1(n416), .Y(n426) );
  OAI22XL U415 ( .A0(n1012), .A1(n419), .B0(n1010), .B1(n439), .Y(n432) );
  OAI22XL U416 ( .A0(n1024), .A1(n404), .B0(n6), .B1(n436), .Y(n431) );
  OAI22XL U417 ( .A0(n1116), .A1(n215), .B0(n9), .B1(n209), .Y(n224) );
  INVXL U418 ( .A(n101), .Y(n130) );
  OAI22XL U419 ( .A0(n990), .A1(n765), .B0(n10), .B1(n103), .Y(n131) );
  OAI22XL U420 ( .A0(n1024), .A1(n771), .B0(n6), .B1(n115), .Y(n135) );
  OR2XL U421 ( .A(n775), .B(n774), .Y(n133) );
  OAI22XL U422 ( .A0(n686), .A1(n639), .B0(n10), .B1(n638), .Y(n667) );
  OAI22XL U423 ( .A0(n56), .A1(n658), .B0(n93), .B1(n637), .Y(n668) );
  XNOR2XL U424 ( .A(n943), .B(n1090), .Y(n639) );
  CMPR32X1 U425 ( .A(n636), .B(n55), .C(n634), .CO(n676), .S(n675) );
  OAI22XL U426 ( .A0(n56), .A1(n637), .B0(n93), .B1(n627), .Y(n636) );
  INVX1 U427 ( .A(n54), .Y(n55) );
  INVXL U428 ( .A(n635), .Y(n54) );
  INVXL U429 ( .A(n1168), .Y(n1169) );
  NOR2XL U430 ( .A(n8), .B(n1167), .Y(n1172) );
  NOR2XL U431 ( .A(n8), .B(n1160), .Y(n1183) );
  INVXL U432 ( .A(n1173), .Y(n1182) );
  NAND2X1 U433 ( .A(n717), .B(n80), .Y(n1203) );
  NOR2X1 U434 ( .A(n732), .B(n731), .Y(n1197) );
  OAI22XL U435 ( .A0(n1024), .A1(n863), .B0(n6), .B1(n832), .Y(n844) );
  OAI22X2 U436 ( .A0(n1163), .A1(n858), .B0(n1014), .B1(n827), .Y(n861) );
  OAI22XL U437 ( .A0(n1024), .A1(n894), .B0(n6), .B1(n863), .Y(n875) );
  OAI22X2 U438 ( .A0(n1163), .A1(n889), .B0(n1014), .B1(n858), .Y(n892) );
  OAI22XL U439 ( .A0(n1024), .A1(n930), .B0(n6), .B1(n894), .Y(n909) );
  ADDFX2 U440 ( .A(n1076), .B(n1075), .CI(n1074), .CO(n1085), .S(n1088) );
  OAI22XL U441 ( .A0(n979), .A1(n1090), .B0(n643), .B1(n1089), .Y(n1250) );
  NAND2XL U442 ( .A(n644), .B(n979), .Y(n1249) );
  NAND2BXL U443 ( .AN(n1090), .B(n648), .Y(n644) );
  NAND2XL U444 ( .A(n1250), .B(n1249), .Y(n1251) );
  INVXL U445 ( .A(n1204), .Y(n1217) );
  NOR2X1 U446 ( .A(n1316), .B(n1317), .Y(n337) );
  INVXL U447 ( .A(n364), .Y(n354) );
  NAND2XL U448 ( .A(n1219), .B(n1222), .Y(n1253) );
  NOR2X1 U449 ( .A(n1311), .B(n1310), .Y(n323) );
  NOR2X1 U450 ( .A(n1100), .B(n368), .Y(n360) );
  NAND2XL U451 ( .A(n1318), .B(n1319), .Y(n358) );
  INVXL U452 ( .A(n1282), .Y(n1190) );
  NAND2XL U453 ( .A(n1220), .B(n1191), .Y(n1193) );
  INVXL U454 ( .A(n1279), .Y(n1194) );
  INVXL U455 ( .A(n306), .Y(n277) );
  NAND2XL U456 ( .A(n303), .B(n307), .Y(n279) );
  INVXL U457 ( .A(n1289), .Y(n280) );
  INVXL U458 ( .A(n303), .Y(n305) );
  INVXL U459 ( .A(n275), .Y(n307) );
  AOI21XL U460 ( .A0(n339), .A1(n320), .B0(n319), .Y(n321) );
  NAND2XL U461 ( .A(n1310), .B(n1311), .Y(n324) );
  INVXL U462 ( .A(n357), .Y(n359) );
  INVXL U463 ( .A(n361), .Y(n362) );
  NAND2XL U464 ( .A(n1320), .B(n1321), .Y(n364) );
  INVXL U465 ( .A(n1270), .Y(n531) );
  XNOR2XL U466 ( .A(n648), .B(A[11]), .Y(n544) );
  XNOR2XL U467 ( .A(n938), .B(n1090), .Y(n558) );
  XNOR2XL U468 ( .A(n943), .B(n937), .Y(n491) );
  XNOR2XL U469 ( .A(n972), .B(n966), .Y(n489) );
  XNOR2XL U470 ( .A(n7), .B(A[11]), .Y(n490) );
  XNOR2XL U471 ( .A(n972), .B(n1090), .Y(n603) );
  XNOR2XL U472 ( .A(n943), .B(n966), .Y(n604) );
  XNOR2XL U473 ( .A(n7), .B(A[7]), .Y(n689) );
  XNOR2XL U474 ( .A(n7), .B(n925), .Y(n583) );
  XNOR2XL U475 ( .A(n7), .B(n1151), .Y(n806) );
  XNOR2XL U476 ( .A(n943), .B(n1112), .Y(n807) );
  XNOR2XL U477 ( .A(n7), .B(n1136), .Y(n837) );
  XNOR2XL U478 ( .A(n943), .B(n933), .Y(n838) );
  XNOR2XL U479 ( .A(n7), .B(n1112), .Y(n868) );
  XNOR2XL U480 ( .A(n943), .B(A[18]), .Y(n869) );
  XNOR2XL U481 ( .A(n1161), .B(n1090), .Y(n400) );
  XNOR2X1 U482 ( .A(n972), .B(A[6]), .Y(n458) );
  XNOR2XL U483 ( .A(n648), .B(n940), .Y(n440) );
  XNOR2XL U484 ( .A(n107), .B(A[18]), .Y(n174) );
  XNOR2XL U485 ( .A(n963), .B(n925), .Y(n465) );
  XNOR2XL U486 ( .A(n7), .B(A[12]), .Y(n460) );
  XNOR2XL U487 ( .A(n1117), .B(n642), .Y(n451) );
  XNOR2XL U488 ( .A(n648), .B(n922), .Y(n450) );
  INVXL U489 ( .A(n171), .Y(n172) );
  XNOR2XL U490 ( .A(n963), .B(A[25]), .Y(n171) );
  XNOR2XL U491 ( .A(n107), .B(n962), .Y(n122) );
  XNOR2XL U492 ( .A(n7), .B(A[6]), .Y(n690) );
  XNOR2XL U493 ( .A(n943), .B(A[4]), .Y(n684) );
  AOI21XL U494 ( .A0(n159), .A1(n158), .B0(n157), .Y(n160) );
  INVXL U495 ( .A(n1284), .Y(n157) );
  INVXL U496 ( .A(n1278), .Y(n1221) );
  NAND2X1 U497 ( .A(n316), .B(n148), .Y(n150) );
  AOI21X2 U498 ( .A0(n146), .A1(n361), .B0(n145), .Y(n348) );
  OAI21XL U499 ( .A0(n357), .A1(n364), .B0(n358), .Y(n145) );
  NAND2XL U500 ( .A(n1191), .B(n1282), .Y(n166) );
  XNOR2X1 U501 ( .A(n156), .B(n155), .Y(PRODUCT[35]) );
  NAND2XL U502 ( .A(n158), .B(n1284), .Y(n155) );
  XNOR2X1 U503 ( .A(n208), .B(n207), .Y(PRODUCT[34]) );
  NAND2XL U504 ( .A(n206), .B(n1286), .Y(n207) );
  NAND2XL U505 ( .A(n233), .B(n1288), .Y(n234) );
  XNOR2X1 U506 ( .A(n1266), .B(n50), .Y(PRODUCT[29]) );
  AND2XL U507 ( .A(n314), .B(n313), .Y(n50) );
  XNOR2X1 U508 ( .A(n327), .B(n326), .Y(PRODUCT[28]) );
  NAND2XL U509 ( .A(n325), .B(n324), .Y(n326) );
  OAI21XL U510 ( .A0(n322), .A1(n1104), .B0(n321), .Y(n327) );
  XNOR2X1 U511 ( .A(n336), .B(n335), .Y(PRODUCT[27]) );
  OAI21XL U512 ( .A0(n1104), .A1(n331), .B0(n330), .Y(n336) );
  XNOR2X1 U513 ( .A(n346), .B(n345), .Y(PRODUCT[26]) );
  NAND2XL U514 ( .A(n370), .B(n369), .Y(n371) );
  INVXL U515 ( .A(n1293), .Y(n1105) );
  OAI22XL U516 ( .A0(n979), .A1(n520), .B0(n466), .B1(n1089), .Y(n519) );
  NAND2BXL U517 ( .AN(n1090), .B(n1117), .Y(n467) );
  INVXL U518 ( .A(n972), .Y(n596) );
  CMPR32X1 U519 ( .A(n600), .B(n599), .C(n598), .CO(n607), .S(n726) );
  OAI22XL U520 ( .A0(n1024), .A1(n602), .B0(n6), .B1(n580), .Y(n598) );
  OAI22XL U521 ( .A0(n990), .A1(n560), .B0(n10), .B1(n524), .Y(n564) );
  OAI22XL U522 ( .A0(n1012), .A1(n556), .B0(n1010), .B1(n522), .Y(n566) );
  OAI22XL U523 ( .A0(n56), .A1(n559), .B0(n93), .B1(n523), .Y(n565) );
  ADDFX2 U524 ( .A(n586), .B(n585), .CI(n584), .CO(n589), .S(n605) );
  OAI22XL U525 ( .A0(n56), .A1(n583), .B0(n93), .B1(n559), .Y(n584) );
  OAI22XL U526 ( .A0(n984), .A1(n558), .B0(n9), .B1(n557), .Y(n585) );
  OAI22XL U527 ( .A0(n965), .A1(n581), .B0(n1010), .B1(n556), .Y(n586) );
  XNOR2XL U528 ( .A(n1117), .B(A[25]), .Y(n1153) );
  XNOR2XL U529 ( .A(n107), .B(n1151), .Y(n1152) );
  XNOR2XL U530 ( .A(n107), .B(n1136), .Y(n1137) );
  XNOR2XL U531 ( .A(n107), .B(n933), .Y(n190) );
  XNOR2XL U532 ( .A(n1161), .B(n1112), .Y(n189) );
  OAI22XL U533 ( .A0(n984), .A1(n521), .B0(n9), .B1(n514), .Y(n537) );
  OAI22XL U534 ( .A0(n1018), .A1(n513), .B0(n1016), .B1(n512), .Y(n538) );
  ADDFX2 U535 ( .A(n682), .B(n681), .CI(n680), .CO(n725), .S(n730) );
  OAI22XL U536 ( .A0(n686), .A1(n684), .B0(n10), .B1(n604), .Y(n680) );
  OAI22X1 U537 ( .A0(n1024), .A1(n603), .B0(n6), .B1(n602), .Y(n681) );
  OAI22XL U538 ( .A0(n965), .A1(n695), .B0(n1010), .B1(n601), .Y(n682) );
  ADDFX2 U539 ( .A(n721), .B(n720), .CI(n719), .CO(n606), .S(n738) );
  OAI22XL U540 ( .A0(n56), .A1(n689), .B0(n93), .B1(n583), .Y(n719) );
  OAI22XL U541 ( .A0(n990), .A1(n604), .B0(n10), .B1(n582), .Y(n720) );
  OAI22X1 U542 ( .A0(n965), .A1(n601), .B0(n1010), .B1(n581), .Y(n721) );
  XNOR2XL U543 ( .A(n648), .B(n1151), .Y(n866) );
  ADDFX2 U544 ( .A(n841), .B(n840), .CI(n839), .CO(n850), .S(n880) );
  OAI22XL U545 ( .A0(n990), .A1(n838), .B0(n10), .B1(n807), .Y(n839) );
  OAI22X1 U546 ( .A0(n56), .A1(n837), .B0(n93), .B1(n806), .Y(n840) );
  XNOR2XL U547 ( .A(n648), .B(n1112), .Y(n934) );
  XNOR2XL U548 ( .A(n648), .B(n1136), .Y(n897) );
  CMPR32X1 U549 ( .A(n872), .B(n871), .C(n870), .CO(n881), .S(n914) );
  OAI22XL U550 ( .A0(n990), .A1(n869), .B0(n10), .B1(n838), .Y(n870) );
  OAI22XL U551 ( .A0(n56), .A1(n868), .B0(n93), .B1(n837), .Y(n871) );
  XNOR2X1 U552 ( .A(n938), .B(A[11]), .Y(n900) );
  XNOR2XL U553 ( .A(n7), .B(n933), .Y(n901) );
  XNOR2XL U554 ( .A(n943), .B(n940), .Y(n903) );
  CMPR32X1 U555 ( .A(n906), .B(n905), .C(n904), .CO(n915), .S(n955) );
  OAI22XL U556 ( .A0(n990), .A1(n903), .B0(n10), .B1(n869), .Y(n904) );
  OAI22XL U557 ( .A0(n56), .A1(n901), .B0(n93), .B1(n868), .Y(n905) );
  XNOR2XL U558 ( .A(n938), .B(n937), .Y(n982) );
  XNOR2XL U559 ( .A(n938), .B(n899), .Y(n939) );
  XNOR2XL U560 ( .A(n7), .B(n940), .Y(n985) );
  XNOR2XL U561 ( .A(n7), .B(A[18]), .Y(n941) );
  XNOR2XL U562 ( .A(n943), .B(n942), .Y(n988) );
  XNOR2XL U563 ( .A(n943), .B(n902), .Y(n944) );
  XNOR2X1 U564 ( .A(n972), .B(A[11]), .Y(n1022) );
  OAI22XL U565 ( .A0(n979), .A1(n978), .B0(n977), .B1(n976), .Y(n1026) );
  XNOR2XL U566 ( .A(n963), .B(n962), .Y(n1009) );
  XNOR2XL U567 ( .A(n7), .B(n962), .Y(n412) );
  XNOR2XL U568 ( .A(n972), .B(A[7]), .Y(n405) );
  XNOR2XL U569 ( .A(n1117), .B(n980), .Y(n407) );
  XNOR2XL U570 ( .A(n7), .B(n922), .Y(n410) );
  XNOR2XL U571 ( .A(n938), .B(n966), .Y(n418) );
  XNOR2XL U572 ( .A(n963), .B(n937), .Y(n420) );
  XNOR2X1 U573 ( .A(n938), .B(A[6]), .Y(n417) );
  XNOR2XL U574 ( .A(n943), .B(A[12]), .Y(n416) );
  XNOR2XL U575 ( .A(n1117), .B(A[4]), .Y(n406) );
  XNOR2XL U576 ( .A(n963), .B(n899), .Y(n419) );
  INVXL U577 ( .A(n194), .Y(n183) );
  OAI22XL U578 ( .A0(n1018), .A1(n210), .B0(n1156), .B1(n182), .Y(n216) );
  OAI22XL U579 ( .A0(n1024), .A1(n211), .B0(n6), .B1(n180), .Y(n218) );
  XNOR2XL U580 ( .A(n972), .B(n1159), .Y(n211) );
  XNOR2XL U581 ( .A(n214), .B(n902), .Y(n127) );
  OAI22X1 U582 ( .A0(n1163), .A1(n109), .B0(n1014), .B1(n125), .Y(n112) );
  ADDFX2 U583 ( .A(n120), .B(n119), .CI(n118), .CO(n294), .S(n136) );
  OAI22XL U584 ( .A0(n1024), .A1(n115), .B0(n6), .B1(n114), .Y(n120) );
  OAI22XL U585 ( .A0(n979), .A1(n656), .B0(n628), .B1(n1089), .Y(n641) );
  OAI22XL U586 ( .A0(n990), .A1(n630), .B0(n10), .B1(n629), .Y(n640) );
  INVXL U587 ( .A(n943), .Y(n630) );
  XNOR2XL U588 ( .A(n7), .B(n980), .Y(n637) );
  NAND2BXL U589 ( .AN(n1090), .B(n963), .Y(n622) );
  ADDFX2 U590 ( .A(n633), .B(n632), .CI(n631), .CO(n710), .S(n634) );
  OAI22XL U591 ( .A0(n990), .A1(n638), .B0(n10), .B1(n626), .Y(n631) );
  OAI22X1 U592 ( .A0(n979), .A1(n628), .B0(n624), .B1(n1089), .Y(n632) );
  ADDFX2 U593 ( .A(n705), .B(n704), .CI(n703), .CO(n729), .S(n706) );
  OAI22X1 U594 ( .A0(n686), .A1(n685), .B0(n10), .B1(n684), .Y(n704) );
  OAI22XL U595 ( .A0(n56), .A1(n683), .B0(n93), .B1(n690), .Y(n705) );
  OAI22XL U596 ( .A0(n965), .A1(n696), .B0(n1010), .B1(n695), .Y(n697) );
  NOR2BXL U597 ( .AN(n1090), .B(n6), .Y(n699) );
  OAI22XL U598 ( .A0(n990), .A1(n626), .B0(n10), .B1(n685), .Y(n700) );
  OAI22X1 U599 ( .A0(n965), .A1(n625), .B0(n1010), .B1(n696), .Y(n701) );
  NAND2XL U600 ( .A(n1222), .B(n1278), .Y(n1212) );
  NAND2BXL U601 ( .AN(n1090), .B(n7), .Y(n652) );
  OAI22XL U602 ( .A0(n990), .A1(n582), .B0(n10), .B1(n560), .Y(n592) );
  OAI22XL U603 ( .A0(n1024), .A1(n580), .B0(n6), .B1(n561), .Y(n591) );
  OAI22XL U604 ( .A0(n1024), .A1(n561), .B0(n6), .B1(n543), .Y(n578) );
  OAI22XL U605 ( .A0(n1018), .A1(n1118), .B0(n1156), .B1(n1138), .Y(n1141) );
  OAI22XL U606 ( .A0(n1163), .A1(n1119), .B0(n1014), .B1(n1135), .Y(n1140) );
  OAI22XL U607 ( .A0(n1018), .A1(n192), .B0(n1156), .B1(n1118), .Y(n1125) );
  NOR2XL U608 ( .A(n8), .B(n1113), .Y(n1134) );
  OAI2BB1XL U609 ( .A0N(n9), .A1N(n1116), .B0(n1115), .Y(n1132) );
  XNOR2XL U610 ( .A(n107), .B(n1112), .Y(n1113) );
  NAND2X1 U611 ( .A(n747), .B(n1187), .Y(n718) );
  OAI22XL U612 ( .A0(n1024), .A1(n780), .B0(n6), .B1(n771), .Y(n795) );
  OAI22XL U613 ( .A0(n990), .A1(n777), .B0(n10), .B1(n765), .Y(n792) );
  XNOR2XL U614 ( .A(n1117), .B(n962), .Y(n789) );
  XNOR2XL U615 ( .A(n972), .B(n902), .Y(n832) );
  OAI22XL U616 ( .A0(n935), .A1(n835), .B0(n783), .B1(n1089), .Y(n834) );
  XNOR2X1 U617 ( .A(n779), .B(n778), .Y(n64) );
  XNOR2XL U618 ( .A(n1117), .B(A[12]), .Y(n828) );
  XNOR2X1 U619 ( .A(n1161), .B(n899), .Y(n827) );
  XNOR2XL U620 ( .A(n972), .B(n942), .Y(n863) );
  XNOR2XL U621 ( .A(n963), .B(n940), .Y(n857) );
  XNOR2XL U622 ( .A(n1117), .B(A[11]), .Y(n859) );
  XNOR2XL U623 ( .A(n1161), .B(n937), .Y(n858) );
  XNOR2XL U624 ( .A(n972), .B(n922), .Y(n894) );
  XNOR2X1 U625 ( .A(n1161), .B(A[6]), .Y(n967) );
  XNOR2XL U626 ( .A(n1117), .B(n925), .Y(n968) );
  XNOR2XL U627 ( .A(n963), .B(n942), .Y(n923) );
  XNOR2XL U628 ( .A(n963), .B(n902), .Y(n888) );
  XNOR2XL U629 ( .A(n1117), .B(n937), .Y(n926) );
  XNOR2XL U630 ( .A(n1117), .B(n899), .Y(n890) );
  XNOR2XL U631 ( .A(n1161), .B(n925), .Y(n889) );
  XNOR2XL U632 ( .A(n972), .B(A[12]), .Y(n973) );
  XNOR2XL U633 ( .A(n972), .B(n962), .Y(n930) );
  CMPR32X1 U634 ( .A(n947), .B(n946), .C(n945), .CO(n956), .S(n1001) );
  OAI22XL U635 ( .A0(n990), .A1(n944), .B0(n10), .B1(n903), .Y(n945) );
  OAI22XL U636 ( .A0(n56), .A1(n941), .B0(n93), .B1(n901), .Y(n946) );
  OAI22XL U637 ( .A0(n5), .A1(n939), .B0(n9), .B1(n900), .Y(n947) );
  OAI22XL U638 ( .A0(n1012), .A1(n439), .B0(n1010), .B1(n1011), .Y(n1058) );
  OAI22XL U639 ( .A0(n1024), .A1(n436), .B0(n6), .B1(n1023), .Y(n1052) );
  OAI22XL U640 ( .A0(n56), .A1(n409), .B0(n93), .B1(n986), .Y(n1029) );
  OAI22XL U641 ( .A0(n984), .A1(n408), .B0(n9), .B1(n983), .Y(n1031) );
  NOR2XL U642 ( .A(n8), .B(n169), .Y(n187) );
  XNOR2XL U643 ( .A(n107), .B(n940), .Y(n169) );
  NAND2XL U644 ( .A(n484), .B(n454), .Y(n452) );
  ADDFX2 U645 ( .A(n527), .B(n526), .CI(n525), .CO(n506), .S(n1091) );
  ADDFX2 U646 ( .A(n269), .B(n268), .CI(n267), .CO(n271), .S(n298) );
  NOR2XL U647 ( .A(n8), .B(n212), .Y(n241) );
  OAI22X1 U648 ( .A0(n1163), .A1(n247), .B0(n1014), .B1(n213), .Y(n240) );
  INVXL U649 ( .A(n220), .Y(n242) );
  OAI22X1 U650 ( .A0(n1024), .A1(n249), .B0(n6), .B1(n211), .Y(n243) );
  OAI22X1 U651 ( .A0(n1018), .A1(n253), .B0(n1156), .B1(n210), .Y(n244) );
  OAI22XL U652 ( .A0(n1116), .A1(n126), .B0(n9), .B1(n252), .Y(n258) );
  OAI22X1 U653 ( .A0(n1163), .A1(n125), .B0(n1014), .B1(n248), .Y(n259) );
  OAI22XL U654 ( .A0(n965), .A1(n124), .B0(n1010), .B1(n246), .Y(n260) );
  OAI22XL U655 ( .A0(n1024), .A1(n250), .B0(n6), .B1(n249), .Y(n264) );
  OAI22XL U656 ( .A0(n965), .A1(n246), .B0(n1010), .B1(n245), .Y(n266) );
  CMPR32X1 U657 ( .A(n263), .B(n262), .C(n261), .CO(n285), .S(n754) );
  OAI2BB1XL U658 ( .A0N(n10), .A1N(n990), .B0(n238), .Y(n261) );
  INVXL U659 ( .A(n237), .Y(n238) );
  OAI22XL U660 ( .A0(n1116), .A1(n252), .B0(n9), .B1(n251), .Y(n288) );
  CMPR32X1 U661 ( .A(n102), .B(n101), .C(n100), .CO(n290), .S(n140) );
  OAI2BB1XL U662 ( .A0N(n93), .A1N(n56), .B0(n95), .Y(n100) );
  XNOR2XL U663 ( .A(n107), .B(A[12]), .Y(n92) );
  OAI22XL U664 ( .A0(n979), .A1(n643), .B0(n649), .B1(n1089), .Y(n646) );
  NOR2BXL U665 ( .AN(n1090), .B(n93), .Y(n645) );
  XNOR2XL U666 ( .A(n7), .B(n1090), .Y(n651) );
  NOR2BXL U667 ( .AN(n1090), .B(n10), .Y(n671) );
  OAI22XL U668 ( .A0(n979), .A1(n657), .B0(n656), .B1(n1089), .Y(n670) );
  OAI22XL U669 ( .A0(n56), .A1(n659), .B0(n93), .B1(n658), .Y(n669) );
  INVXL U670 ( .A(n1263), .Y(n1264) );
  OR2XL U671 ( .A(n1255), .B(n1261), .Y(n1265) );
  NAND2XL U672 ( .A(n1229), .B(n1276), .Y(n1230) );
  NOR2XL U673 ( .A(n655), .B(n654), .Y(n1240) );
  NAND2XL U674 ( .A(n655), .B(n654), .Y(n1241) );
  AOI21XL U675 ( .A0(n1246), .A1(n1247), .B0(n647), .Y(n1243) );
  INVXL U676 ( .A(n1245), .Y(n647) );
  NAND2BX1 U677 ( .AN(n1197), .B(n1203), .Y(n79) );
  ADDFX2 U678 ( .A(n735), .B(n734), .CI(n733), .CO(n614), .S(n740) );
  OAI22XL U679 ( .A0(n1163), .A1(n1147), .B0(n1014), .B1(n1162), .Y(n1180) );
  NAND2X1 U680 ( .A(n740), .B(n739), .Y(n1198) );
  NOR2X1 U681 ( .A(n740), .B(n739), .Y(n1200) );
  NAND2XL U682 ( .A(n779), .B(n62), .Y(n60) );
  OAI21XL U683 ( .A0(n779), .A1(n62), .B0(n778), .Y(n61) );
  NAND2XL U684 ( .A(n646), .B(n645), .Y(n1245) );
  INVXL U685 ( .A(n1251), .Y(n1247) );
  NAND2XL U686 ( .A(n664), .B(n663), .Y(n1237) );
  AOI21XL U687 ( .A0(n1238), .A1(n662), .B0(n665), .Y(n1235) );
  INVXL U688 ( .A(n1237), .Y(n665) );
  NOR2XL U689 ( .A(n673), .B(n672), .Y(n1232) );
  NAND2XL U690 ( .A(n673), .B(n672), .Y(n1233) );
  NOR2XL U691 ( .A(n1108), .B(n1107), .Y(mult_x_1_n151) );
  NOR2XL U692 ( .A(n1158), .B(n1157), .Y(mult_x_1_n120) );
  XOR2XL U693 ( .A(n1244), .B(n1243), .Y(n1351) );
  NAND2XL U694 ( .A(n1242), .B(n1241), .Y(n1244) );
  INVXL U695 ( .A(n1240), .Y(n1242) );
  XOR2X1 U696 ( .A(n743), .B(n742), .Y(n1344) );
  INVXL U697 ( .A(n1203), .Y(n743) );
  NAND2XL U698 ( .A(n747), .B(n746), .Y(n748) );
  NOR2XL U699 ( .A(n1128), .B(n1127), .Y(mult_x_1_n136) );
  XOR2X1 U700 ( .A(n78), .B(n76), .Y(n1343) );
  NOR2X1 U701 ( .A(n77), .B(n1200), .Y(n76) );
  NAND2X1 U702 ( .A(n79), .B(n1199), .Y(n78) );
  NAND2XL U703 ( .A(n1177), .B(n1176), .Y(mult_x_1_n58) );
  NAND2XL U704 ( .A(n1175), .B(n1174), .Y(n1176) );
  NOR2XL U705 ( .A(n1185), .B(n1184), .Y(mult_x_1_n109) );
  NAND2XL U706 ( .A(n1185), .B(n1184), .Y(mult_x_1_n110) );
  NAND2XL U707 ( .A(n1158), .B(n1157), .Y(mult_x_1_n121) );
  NOR2XL U708 ( .A(n1143), .B(n1142), .Y(mult_x_1_n129) );
  NAND2XL U709 ( .A(n1143), .B(n1142), .Y(mult_x_1_n130) );
  NAND2XL U710 ( .A(n1128), .B(n1127), .Y(mult_x_1_n137) );
  NAND2XL U711 ( .A(n1330), .B(n1126), .Y(mult_x_1_n86) );
  NAND2X1 U712 ( .A(n87), .B(n86), .Y(n1007) );
  NAND2X1 U713 ( .A(n1044), .B(n1046), .Y(n86) );
  OAI21XL U714 ( .A0(n1044), .A1(n1046), .B0(n1045), .Y(n87) );
  XOR2X1 U715 ( .A(n85), .B(n1045), .Y(n1047) );
  INVX1 U716 ( .A(n1069), .Y(n58) );
  OAI2BB1X1 U717 ( .A0N(n1079), .A1N(n1078), .B0(n88), .Y(n1084) );
  ADDFX2 U718 ( .A(n1088), .B(n1087), .CI(n1086), .CO(mult_x_1_n665), .S(n473)
         );
  XNOR3X2 U719 ( .A(n1079), .B(n1078), .C(n89), .Y(n1086) );
  NOR2BXL U720 ( .AN(n1090), .B(n1089), .Y(n1354) );
  XNOR2XL U721 ( .A(n1248), .B(n1247), .Y(n1352) );
  NAND2XL U722 ( .A(n1246), .B(n1245), .Y(n1248) );
  XNOR2XL U723 ( .A(n1239), .B(n1238), .Y(n1350) );
  NAND2XL U724 ( .A(n662), .B(n1237), .Y(n1239) );
  XOR2XL U725 ( .A(n1236), .B(n1235), .Y(n1349) );
  NAND2XL U726 ( .A(n1234), .B(n1233), .Y(n1236) );
  INVXL U727 ( .A(n1232), .Y(n1234) );
  XOR2XL U728 ( .A(n1218), .B(n1217), .Y(n1348) );
  NAND2XL U729 ( .A(n1216), .B(n1215), .Y(n1218) );
  INVXL U730 ( .A(n1214), .Y(n1216) );
  NAND2XL U731 ( .A(n1207), .B(n1206), .Y(n1208) );
  NAND2XL U732 ( .A(n1187), .B(n1186), .Y(n1188) );
  INVX1 U733 ( .A(B[7]), .Y(n623) );
  OR2X2 U734 ( .A(n1098), .B(n1097), .Y(n53) );
  ADDFHX1 U735 ( .A(n497), .B(n496), .CI(n495), .CO(n475), .S(n505) );
  CMPR22X1 U736 ( .A(n865), .B(n864), .CO(n842), .S(n874) );
  CMPR22X1 U737 ( .A(n932), .B(n931), .CO(n907), .S(n949) );
  CMPR22X1 U738 ( .A(n975), .B(n974), .CO(n948), .S(n995) );
  CMPR22X1 U739 ( .A(n1028), .B(n1027), .CO(n1035), .S(n1057) );
  OAI22X1 U740 ( .A0(n979), .A1(n693), .B0(n593), .B1(n1089), .Y(n692) );
  XNOR2X1 U741 ( .A(n449), .B(n448), .Y(n484) );
  AND2X1 U742 ( .A(n449), .B(n448), .Y(n457) );
  OAI22XL U743 ( .A0(n1170), .A1(n395), .B0(n104), .B1(n394), .Y(n449) );
  CMPR22X1 U744 ( .A(n782), .B(n781), .CO(n794), .S(n812) );
  CMPR22X1 U745 ( .A(n563), .B(n562), .CO(n577), .S(n590) );
  CMPR22X1 U746 ( .A(n688), .B(n687), .CO(n703), .S(n711) );
  OAI22X1 U747 ( .A0(n965), .A1(n623), .B0(n1010), .B1(n622), .Y(n687) );
  XNOR3X2 U748 ( .A(n485), .B(n484), .C(n483), .Y(n526) );
  CMPR22X1 U749 ( .A(n692), .B(n691), .CO(n727), .S(n723) );
  OAI22X1 U750 ( .A0(n597), .A1(n596), .B0(n595), .B1(n594), .Y(n691) );
  NAND2X1 U751 ( .A(n378), .B(n377), .Y(n379) );
  XNOR2X1 U752 ( .A(n372), .B(n371), .Y(PRODUCT[22]) );
  NOR2X1 U753 ( .A(n1309), .B(n1308), .Y(n312) );
  AOI21XL U754 ( .A0(n1226), .A1(n1219), .B0(n1223), .Y(n1210) );
  AOI21XL U755 ( .A0(n1226), .A1(n1225), .B0(n1224), .Y(n1227) );
  AOI21XL U756 ( .A0(n1226), .A1(n1191), .B0(n1190), .Y(n1192) );
  BUFX3 U757 ( .A(n987), .Y(n56) );
  XOR2X1 U758 ( .A(n373), .B(n1106), .Y(PRODUCT[17]) );
  XOR2X1 U759 ( .A(n1068), .B(n1069), .Y(n59) );
  XOR2X1 U760 ( .A(n877), .B(n878), .Y(n67) );
  XOR2X1 U761 ( .A(n845), .B(n70), .Y(n883) );
  XOR2X1 U762 ( .A(n846), .B(n847), .Y(n70) );
  XOR2X1 U763 ( .A(n952), .B(n953), .Y(n73) );
  OR2X2 U764 ( .A(n744), .B(n718), .Y(n80) );
  OAI21X1 U765 ( .A0(n382), .A1(n376), .B0(n377), .Y(n81) );
  NOR2X1 U766 ( .A(n677), .B(n676), .Y(n1205) );
  OAI22X1 U767 ( .A0(n1116), .A1(n546), .B0(n9), .B1(n545), .Y(n562) );
  AOI21X1 U768 ( .A0(n276), .A1(n152), .B0(n151), .Y(n1262) );
  NOR2X1 U769 ( .A(n1324), .B(n1325), .Y(n1100) );
  OAI21XL U770 ( .A0(n1266), .A1(n1255), .B0(n1262), .Y(n235) );
  OAI21XL U771 ( .A0(n1266), .A1(n205), .B0(n204), .Y(n208) );
  XNOR2X1 U772 ( .A(n352), .B(n351), .Y(PRODUCT[25]) );
  AOI21XL U773 ( .A0(n1223), .A1(n1222), .B0(n1221), .Y(n1256) );
  NAND2X1 U774 ( .A(n1309), .B(n1308), .Y(n313) );
  AOI21XL U775 ( .A0(n339), .A1(n316), .B0(n318), .Y(n330) );
  XNOR2X1 U776 ( .A(n532), .B(n1297), .Y(PRODUCT[15]) );
  XNOR2XL U777 ( .A(n7), .B(n899), .Y(n523) );
  XNOR2XL U778 ( .A(n972), .B(A[24]), .Y(n180) );
  OAI22X1 U779 ( .A0(n1163), .A1(n399), .B0(n1014), .B1(n398), .Y(n401) );
  OAI22X1 U780 ( .A0(n1018), .A1(n116), .B0(n1156), .B1(n121), .Y(n119) );
  OAI22X1 U781 ( .A0(n1163), .A1(n967), .B0(n1014), .B1(n924), .Y(n970) );
  OAI22X1 U782 ( .A0(n1163), .A1(n398), .B0(n1014), .B1(n393), .Y(n429) );
  XOR2X1 U783 ( .A(B[12]), .B(B[13]), .Y(n90) );
  XNOR2X1 U784 ( .A(B[12]), .B(B[11]), .Y(n390) );
  CLKINVX3 U785 ( .A(B[13]), .Y(n468) );
  XNOR2X1 U786 ( .A(n1117), .B(n922), .Y(n767) );
  BUFX3 U787 ( .A(n390), .Y(n1156) );
  INVX8 U788 ( .A(n468), .Y(n1117) );
  XNOR2X1 U789 ( .A(n1117), .B(n942), .Y(n116) );
  OAI22XL U790 ( .A0(n1018), .A1(n767), .B0(n1156), .B1(n116), .Y(n132) );
  XOR2X1 U791 ( .A(B[4]), .B(B[5]), .Y(n91) );
  XNOR2X1 U792 ( .A(B[4]), .B(B[3]), .Y(n411) );
  CLKINVX3 U793 ( .A(B[3]), .Y(n653) );
  OAI22X1 U794 ( .A0(n987), .A1(n128), .B0(n93), .B1(n94), .Y(n101) );
  XNOR2X1 U795 ( .A(B[16]), .B(B[15]), .Y(n168) );
  NOR2XL U796 ( .A(n168), .B(n92), .Y(n102) );
  INVXL U797 ( .A(n94), .Y(n95) );
  XNOR2X1 U798 ( .A(n972), .B(A[18]), .Y(n771) );
  XNOR2X1 U799 ( .A(n972), .B(n933), .Y(n115) );
  CLKINVX3 U800 ( .A(n546), .Y(n214) );
  XNOR2XL U801 ( .A(n214), .B(n940), .Y(n117) );
  OAI22XL U802 ( .A0(n1116), .A1(n127), .B0(n9), .B1(n117), .Y(n134) );
  XNOR2X1 U803 ( .A(B[6]), .B(B[5]), .Y(n173) );
  NAND2X2 U804 ( .A(n98), .B(n173), .Y(n1012) );
  BUFX8 U805 ( .A(n173), .Y(n1010) );
  XNOR2X1 U806 ( .A(n963), .B(n1112), .Y(n106) );
  NAND2X2 U807 ( .A(n99), .B(n104), .Y(n1170) );
  CLKBUFX8 U808 ( .A(n104), .Y(n1014) );
  XNOR2X1 U809 ( .A(n1161), .B(A[12]), .Y(n110) );
  XNOR2X1 U810 ( .A(n972), .B(n1112), .Y(n114) );
  XNOR2X1 U811 ( .A(n972), .B(n1136), .Y(n250) );
  OAI22X1 U812 ( .A0(n990), .A1(n103), .B0(n10), .B1(n123), .Y(n113) );
  XNOR2X1 U813 ( .A(n1161), .B(n962), .Y(n109) );
  XNOR2X1 U814 ( .A(n1161), .B(n922), .Y(n125) );
  XNOR2X1 U815 ( .A(n963), .B(n1136), .Y(n105) );
  XNOR2X1 U816 ( .A(n963), .B(n1151), .Y(n124) );
  OAI22XL U817 ( .A0(n965), .A1(n105), .B0(n1010), .B1(n124), .Y(n111) );
  OAI22X1 U818 ( .A0(n965), .A1(n106), .B0(n1010), .B1(n105), .Y(n770) );
  XNOR2XL U819 ( .A(n107), .B(A[11]), .Y(n108) );
  OAI22XL U820 ( .A0(n1163), .A1(n110), .B0(n1014), .B1(n109), .Y(n768) );
  XNOR2X1 U821 ( .A(n214), .B(A[18]), .Y(n126) );
  OAI22XL U822 ( .A0(n1116), .A1(n117), .B0(n9), .B1(n126), .Y(n118) );
  OAI22X1 U823 ( .A0(n1018), .A1(n121), .B0(n1156), .B1(n254), .Y(n257) );
  XNOR2X1 U824 ( .A(n963), .B(n1159), .Y(n246) );
  XNOR2X1 U825 ( .A(n1161), .B(n942), .Y(n248) );
  XNOR2X1 U826 ( .A(n214), .B(n933), .Y(n252) );
  XNOR2X1 U827 ( .A(n7), .B(n1159), .Y(n776) );
  OAI22X1 U828 ( .A0(n987), .A1(n776), .B0(n93), .B1(n128), .Y(n779) );
  INVX1 U829 ( .A(B[0]), .Y(n976) );
  BUFX3 U830 ( .A(n976), .Y(n1089) );
  NAND2X1 U831 ( .A(B[1]), .B(n976), .Y(n935) );
  CMPR32X1 U832 ( .A(n132), .B(n131), .C(n130), .CO(n141), .S(n803) );
  CMPR32X1 U833 ( .A(n135), .B(n134), .C(n133), .CO(n139), .S(n802) );
  CMPR32X1 U834 ( .A(n138), .B(n137), .C(n136), .CO(n760), .S(n797) );
  CMPR32X1 U835 ( .A(n141), .B(n140), .C(n139), .CO(n144), .S(n796) );
  NOR2X1 U836 ( .A(n1320), .B(n1321), .Y(n353) );
  NOR2X1 U837 ( .A(n1318), .B(n1319), .Y(n357) );
  NOR2X1 U838 ( .A(n353), .B(n357), .Y(n146) );
  NOR2X1 U839 ( .A(n1314), .B(n1315), .Y(n342) );
  NOR2X1 U840 ( .A(n337), .B(n342), .Y(n316) );
  NOR2X1 U841 ( .A(n1291), .B(n1293), .Y(n375) );
  OAI21X2 U842 ( .A0(n1291), .A1(n1294), .B0(n1292), .Y(n374) );
  NAND2X1 U843 ( .A(n1322), .B(n1323), .Y(n369) );
  NAND2X1 U844 ( .A(n1314), .B(n1315), .Y(n343) );
  OAI21XL U845 ( .A0(n342), .A1(n349), .B0(n343), .Y(n318) );
  NAND2XL U846 ( .A(n1312), .B(n1313), .Y(n333) );
  OAI21XL U847 ( .A0(n323), .A1(n333), .B0(n324), .Y(n147) );
  AOI21X1 U848 ( .A0(n148), .A1(n318), .B0(n147), .Y(n149) );
  NOR2X1 U849 ( .A(n312), .B(n309), .Y(n303) );
  NAND2X1 U850 ( .A(n303), .B(n152), .Y(n1255) );
  NOR2X1 U851 ( .A(n1255), .B(n1287), .Y(n202) );
  NAND2XL U852 ( .A(n202), .B(n206), .Y(n154) );
  NAND2XL U853 ( .A(n1307), .B(n1306), .Y(n310) );
  OAI21XL U854 ( .A0(n309), .A1(n313), .B0(n310), .Y(n276) );
  NAND2XL U855 ( .A(n1304), .B(n1305), .Y(n306) );
  OAI21XL U856 ( .A0(n1262), .A1(n1287), .B0(n1288), .Y(n203) );
  AOI21XL U857 ( .A0(n203), .A1(n206), .B0(n159), .Y(n153) );
  OAI21XL U858 ( .A0(n1266), .A1(n154), .B0(n153), .Y(n156) );
  INVXL U859 ( .A(n1220), .Y(n165) );
  OAI21XL U860 ( .A0(n161), .A1(n1288), .B0(n160), .Y(n1259) );
  OAI21XL U861 ( .A0(n1262), .A1(n163), .B0(n162), .Y(n1226) );
  INVXL U862 ( .A(n1226), .Y(n164) );
  OAI21XL U863 ( .A0(n1266), .A1(n165), .B0(n164), .Y(n167) );
  XNOR2X1 U864 ( .A(n1117), .B(n1112), .Y(n182) );
  XNOR2XL U865 ( .A(n1117), .B(n1136), .Y(n178) );
  OAI22XL U866 ( .A0(n1018), .A1(n182), .B0(n1156), .B1(n178), .Y(n188) );
  XNOR2X1 U867 ( .A(n963), .B(A[24]), .Y(n245) );
  OAI22X1 U868 ( .A0(n965), .A1(n245), .B0(n1010), .B1(n171), .Y(n220) );
  XNOR2X1 U869 ( .A(n1161), .B(A[18]), .Y(n181) );
  XNOR2X1 U870 ( .A(n1161), .B(n933), .Y(n177) );
  OAI22XL U871 ( .A0(n1163), .A1(n181), .B0(n1014), .B1(n177), .Y(n185) );
  XNOR2XL U872 ( .A(n214), .B(n1151), .Y(n209) );
  XNOR2XL U873 ( .A(n214), .B(n1159), .Y(n179) );
  OAI22XL U874 ( .A0(n1116), .A1(n209), .B0(n9), .B1(n179), .Y(n184) );
  XNOR2X1 U875 ( .A(n972), .B(A[25]), .Y(n175) );
  OAI22X1 U876 ( .A0(n597), .A1(n180), .B0(n6), .B1(n175), .Y(n194) );
  XNOR2XL U877 ( .A(n1117), .B(n1151), .Y(n192) );
  OAI22XL U878 ( .A0(n1018), .A1(n178), .B0(n1156), .B1(n192), .Y(n197) );
  XNOR2X1 U879 ( .A(n214), .B(A[24]), .Y(n191) );
  OAI22XL U880 ( .A0(n1170), .A1(n213), .B0(n1014), .B1(n181), .Y(n217) );
  CMPR32X1 U881 ( .A(n185), .B(n184), .C(n183), .CO(n201), .S(n226) );
  CMPR32X1 U882 ( .A(n188), .B(n187), .C(n186), .CO(n230), .S(n225) );
  XNOR2X1 U883 ( .A(n1161), .B(n1136), .Y(n1119) );
  INVX4 U884 ( .A(n546), .Y(n938) );
  XNOR2X1 U885 ( .A(n938), .B(A[25]), .Y(n1114) );
  OAI22X1 U886 ( .A0(n1116), .A1(n191), .B0(n9), .B1(n1114), .Y(n1133) );
  XNOR2X1 U887 ( .A(n1117), .B(n1159), .Y(n1118) );
  CMPR32X1 U888 ( .A(n195), .B(n194), .C(n193), .CO(n1124), .S(n200) );
  CMPR32X1 U889 ( .A(n198), .B(n197), .C(n196), .CO(n1123), .S(n199) );
  CMPR32X1 U890 ( .A(n201), .B(n200), .C(n199), .CO(n1109), .S(n229) );
  NAND2XL U891 ( .A(n1108), .B(n1107), .Y(mult_x_1_n152) );
  INVXL U892 ( .A(n202), .Y(n205) );
  INVXL U893 ( .A(n203), .Y(n204) );
  XNOR2X1 U894 ( .A(n214), .B(n1136), .Y(n215) );
  XNOR2X1 U895 ( .A(n1117), .B(A[18]), .Y(n253) );
  XNOR2X1 U896 ( .A(n107), .B(n942), .Y(n212) );
  XNOR2X1 U897 ( .A(n1161), .B(n902), .Y(n247) );
  XNOR2X1 U898 ( .A(n214), .B(n1112), .Y(n251) );
  OAI22XL U899 ( .A0(n1116), .A1(n251), .B0(n9), .B1(n215), .Y(n239) );
  CMPR32X1 U900 ( .A(n218), .B(n217), .C(n216), .CO(n227), .S(n269) );
  CMPR32X1 U901 ( .A(n221), .B(n220), .C(n219), .CO(n186), .S(n268) );
  ADDFHX1 U902 ( .A(n224), .B(n223), .CI(n222), .CO(n272), .S(n267) );
  CMPR32X1 U903 ( .A(n227), .B(n226), .C(n225), .CO(n228), .S(n270) );
  CMPR32X1 U904 ( .A(n230), .B(n229), .C(n228), .CO(n1108), .S(n231) );
  NOR2XL U905 ( .A(n232), .B(n231), .Y(mult_x_1_n160) );
  XNOR2XL U906 ( .A(n107), .B(n922), .Y(n236) );
  NOR2XL U907 ( .A(n8), .B(n236), .Y(n263) );
  CMPR32X1 U908 ( .A(n241), .B(n240), .C(n239), .CO(n222), .S(n284) );
  OAI22XL U909 ( .A0(n1170), .A1(n248), .B0(n1014), .B1(n247), .Y(n265) );
  OAI22XL U910 ( .A0(n1018), .A1(n254), .B0(n1156), .B1(n253), .Y(n287) );
  ADDFHX1 U911 ( .A(n260), .B(n259), .CI(n258), .CO(n755), .S(n292) );
  CMPR32X1 U912 ( .A(n266), .B(n265), .C(n264), .CO(n297), .S(n753) );
  CMPR32X1 U913 ( .A(n272), .B(n271), .C(n270), .CO(n232), .S(n273) );
  NOR2XL U914 ( .A(n274), .B(n273), .Y(mult_x_1_n169) );
  NAND2XL U915 ( .A(n274), .B(n273), .Y(mult_x_1_n170) );
  INVXL U916 ( .A(n276), .Y(n304) );
  AOI21XL U917 ( .A0(n276), .A1(n307), .B0(n277), .Y(n278) );
  CMPR32X1 U918 ( .A(n285), .B(n284), .C(n283), .CO(n300), .S(n752) );
  CMPR32X1 U919 ( .A(n288), .B(n287), .C(n286), .CO(n296), .S(n758) );
  ADDFHX1 U920 ( .A(n297), .B(n296), .CI(n295), .CO(n299), .S(n750) );
  CMPR32X1 U921 ( .A(n300), .B(n299), .C(n298), .CO(n274), .S(n301) );
  NOR2XL U922 ( .A(n302), .B(n301), .Y(mult_x_1_n176) );
  NAND2XL U923 ( .A(n302), .B(n301), .Y(mult_x_1_n177) );
  INVXL U924 ( .A(n309), .Y(n311) );
  INVXL U925 ( .A(n312), .Y(n314) );
  INVXL U926 ( .A(n315), .Y(n347) );
  INVXL U927 ( .A(n316), .Y(n328) );
  NOR2XL U928 ( .A(n328), .B(n332), .Y(n320) );
  NAND2XL U929 ( .A(n347), .B(n320), .Y(n322) );
  INVX1 U930 ( .A(n348), .Y(n339) );
  INVXL U931 ( .A(n318), .Y(n329) );
  OAI21XL U932 ( .A0(n329), .A1(n332), .B0(n333), .Y(n319) );
  INVXL U933 ( .A(n323), .Y(n325) );
  NAND2XL U934 ( .A(n347), .B(n316), .Y(n331) );
  NAND2XL U935 ( .A(n334), .B(n333), .Y(n335) );
  NAND2XL U936 ( .A(n347), .B(n350), .Y(n341) );
  INVXL U937 ( .A(n349), .Y(n338) );
  AOI21X1 U938 ( .A0(n339), .A1(n350), .B0(n338), .Y(n340) );
  OAI21XL U939 ( .A0(n1104), .A1(n341), .B0(n340), .Y(n346) );
  INVXL U940 ( .A(n342), .Y(n344) );
  NAND2XL U941 ( .A(n344), .B(n343), .Y(n345) );
  OAI21XL U942 ( .A0(n1104), .A1(n315), .B0(n348), .Y(n352) );
  NAND2XL U943 ( .A(n350), .B(n349), .Y(n351) );
  INVXL U944 ( .A(n353), .Y(n365) );
  NAND2XL U945 ( .A(n360), .B(n365), .Y(n356) );
  AOI21XL U946 ( .A0(n361), .A1(n365), .B0(n354), .Y(n355) );
  INVXL U947 ( .A(n360), .Y(n363) );
  OAI21XL U948 ( .A0(n1104), .A1(n363), .B0(n362), .Y(n367) );
  NAND2X1 U949 ( .A(n365), .B(n364), .Y(n366) );
  OAI21XL U950 ( .A0(n1104), .A1(n1100), .B0(n1101), .Y(n372) );
  INVXL U951 ( .A(n368), .Y(n370) );
  INVXL U952 ( .A(n376), .Y(n378) );
  INVXL U953 ( .A(n381), .Y(n383) );
  XOR2X1 U954 ( .A(n385), .B(n384), .Y(PRODUCT[19]) );
  INVXL U955 ( .A(n1291), .Y(n387) );
  XNOR2XL U956 ( .A(n107), .B(n650), .Y(n389) );
  NOR2XL U957 ( .A(n8), .B(n389), .Y(n428) );
  BUFX3 U958 ( .A(n390), .Y(n1016) );
  XNOR2XL U959 ( .A(n1117), .B(n966), .Y(n438) );
  OAI22XL U960 ( .A0(n1018), .A1(n406), .B0(n1016), .B1(n438), .Y(n427) );
  XNOR2X1 U961 ( .A(n963), .B(A[11]), .Y(n439) );
  XNOR2X1 U962 ( .A(n972), .B(n937), .Y(n436) );
  BUFX3 U963 ( .A(n935), .Y(n979) );
  BUFX3 U964 ( .A(A[0]), .Y(n1090) );
  XNOR2X1 U965 ( .A(n938), .B(A[7]), .Y(n408) );
  XNOR2X1 U966 ( .A(n938), .B(n925), .Y(n983) );
  XNOR2X1 U967 ( .A(n7), .B(n902), .Y(n986) );
  NOR2BX1 U968 ( .AN(n1090), .B(n8), .Y(n403) );
  OAI22X1 U969 ( .A0(n979), .A1(n397), .B0(n396), .B1(n1089), .Y(n402) );
  OAI22X1 U970 ( .A0(n1024), .A1(n458), .B0(n6), .B1(n405), .Y(n463) );
  OAI22XL U971 ( .A0(n1018), .A1(n451), .B0(n1016), .B1(n407), .Y(n461) );
  CMPR32X1 U972 ( .A(n403), .B(n402), .C(n401), .CO(n423), .S(n456) );
  OAI22X1 U973 ( .A0(n1024), .A1(n405), .B0(n6), .B1(n404), .Y(n415) );
  OAI22X1 U974 ( .A0(n56), .A1(n412), .B0(n93), .B1(n410), .Y(n414) );
  OAI22XL U975 ( .A0(n1018), .A1(n407), .B0(n1016), .B1(n406), .Y(n413) );
  OAI22X1 U976 ( .A0(n984), .A1(n417), .B0(n9), .B1(n408), .Y(n435) );
  OAI22X1 U977 ( .A0(n56), .A1(n410), .B0(n93), .B1(n409), .Y(n434) );
  OAI22X1 U978 ( .A0(n5), .A1(n459), .B0(n9), .B1(n418), .Y(n481) );
  OAI22X1 U979 ( .A0(n5), .A1(n418), .B0(n9), .B1(n417), .Y(n425) );
  ADDFHX1 U980 ( .A(n423), .B(n422), .CI(n421), .CO(n1079), .S(n470) );
  CMPR32X1 U981 ( .A(n426), .B(n425), .C(n424), .CO(n446), .S(n477) );
  CMPR32X1 U982 ( .A(n429), .B(n428), .C(n427), .CO(n1076), .S(n445) );
  CMPR32X1 U983 ( .A(n432), .B(n431), .C(n430), .CO(n1075), .S(n444) );
  XNOR2X1 U984 ( .A(n972), .B(n899), .Y(n1023) );
  OAI22XL U985 ( .A0(n990), .A1(n437), .B0(n10), .B1(n989), .Y(n1051) );
  XNOR2X1 U986 ( .A(n1117), .B(A[6]), .Y(n1017) );
  OAI22XL U987 ( .A0(n1018), .A1(n438), .B0(n1016), .B1(n1017), .Y(n1050) );
  XNOR2X1 U988 ( .A(n648), .B(A[18]), .Y(n978) );
  OAI22X1 U989 ( .A0(n979), .A1(n440), .B0(n978), .B1(n1089), .Y(n1028) );
  XNOR2XL U990 ( .A(n107), .B(n642), .Y(n441) );
  ADDHXL U991 ( .A(n443), .B(n442), .CO(n1056), .S(n430) );
  OAI22X1 U992 ( .A0(n990), .A1(n464), .B0(n10), .B1(n447), .Y(n485) );
  NAND2XL U993 ( .A(n452), .B(n483), .Y(n453) );
  OAI21XL U994 ( .A0(n454), .A1(n484), .B0(n453), .Y(n497) );
  ADDFHX1 U995 ( .A(n457), .B(n456), .CI(n455), .CO(n471), .S(n496) );
  OAI22X1 U996 ( .A0(n5), .A1(n514), .B0(n9), .B1(n459), .Y(n493) );
  XNOR2X1 U997 ( .A(n963), .B(A[7]), .Y(n511) );
  XNOR2X1 U998 ( .A(n648), .B(A[12]), .Y(n520) );
  OAI22XL U999 ( .A0(n1018), .A1(n468), .B0(n1156), .B1(n467), .Y(n518) );
  CMPR32X1 U1000 ( .A(n476), .B(n475), .C(n474), .CO(n472), .S(n499) );
  CMPR32X1 U1001 ( .A(n479), .B(n478), .C(n477), .CO(n469), .S(n507) );
  CMPR32X1 U1002 ( .A(n482), .B(n481), .C(n480), .CO(n479), .S(n527) );
  CMPR32X1 U1003 ( .A(n488), .B(n487), .C(n486), .CO(n483), .S(n536) );
  XNOR2X1 U1004 ( .A(n972), .B(A[4]), .Y(n543) );
  OAI22X1 U1005 ( .A0(n1024), .A1(n543), .B0(n6), .B1(n489), .Y(n542) );
  CMPR32X1 U1006 ( .A(n494), .B(n493), .C(n492), .CO(n510), .S(n534) );
  NOR2XL U1007 ( .A(n499), .B(n498), .Y(mult_x_1_n286) );
  NAND2XL U1008 ( .A(n499), .B(n498), .Y(mult_x_1_n287) );
  CMPR32X1 U1009 ( .A(n507), .B(n506), .C(n505), .CO(n498), .S(n529) );
  ADDFHX1 U1010 ( .A(n510), .B(n509), .CI(n508), .CO(n495), .S(n1093) );
  XNOR2X1 U1011 ( .A(n1117), .B(n1090), .Y(n513) );
  XNOR2X1 U1012 ( .A(n938), .B(n642), .Y(n521) );
  ADDHXL U1013 ( .A(n519), .B(n518), .CO(n515), .S(n555) );
  XNOR2X1 U1014 ( .A(n963), .B(n966), .Y(n556) );
  NOR2XL U1015 ( .A(n529), .B(n528), .Y(mult_x_1_n292) );
  NAND2XL U1016 ( .A(n529), .B(n528), .Y(mult_x_1_n293) );
  CMPR32X1 U1017 ( .A(n539), .B(n538), .C(n537), .CO(n552), .S(n569) );
  ADDFX2 U1018 ( .A(n542), .B(n541), .CI(n540), .CO(n535), .S(n568) );
  XNOR2X1 U1019 ( .A(n972), .B(n980), .Y(n561) );
  OAI22X1 U1020 ( .A0(n979), .A1(n579), .B0(n544), .B1(n1089), .Y(n563) );
  CMPR32X1 U1021 ( .A(n552), .B(n551), .C(n550), .CO(n1092), .S(n1094) );
  ADDFHX1 U1022 ( .A(n555), .B(n554), .CI(n553), .CO(n550), .S(n610) );
  XNOR2X1 U1023 ( .A(n943), .B(A[6]), .Y(n582) );
  XNOR2X1 U1024 ( .A(n972), .B(n642), .Y(n580) );
  CMPR32X1 U1025 ( .A(n566), .B(n565), .C(n564), .CO(n553), .S(n587) );
  NOR2XL U1026 ( .A(n571), .B(n570), .Y(n572) );
  NAND2XL U1027 ( .A(n571), .B(n570), .Y(n573) );
  INVXL U1028 ( .A(n573), .Y(mult_x_1_n305) );
  INVXL U1029 ( .A(n572), .Y(n574) );
  NAND2XL U1030 ( .A(n574), .B(n573), .Y(mult_x_1_n84) );
  CMPR32X1 U1031 ( .A(n578), .B(n577), .C(n576), .CO(n567), .S(n613) );
  OAI22XL U1032 ( .A0(n979), .A1(n593), .B0(n579), .B1(n1089), .Y(n599) );
  XNOR2X1 U1033 ( .A(n972), .B(n650), .Y(n602) );
  ADDFHX1 U1034 ( .A(n589), .B(n588), .CI(n587), .CO(n609), .S(n611) );
  CMPR32X1 U1035 ( .A(n592), .B(n591), .C(n590), .CO(n588), .S(n735) );
  XNOR2X1 U1036 ( .A(n648), .B(n925), .Y(n693) );
  CMPR32X1 U1037 ( .A(n607), .B(n606), .C(n605), .CO(n612), .S(n733) );
  OR2X2 U1038 ( .A(n615), .B(n614), .Y(n1330) );
  CMPR32X1 U1039 ( .A(n610), .B(n609), .C(n608), .CO(n570), .S(n617) );
  OR2X2 U1040 ( .A(n617), .B(n616), .Y(n620) );
  NAND2XL U1041 ( .A(n620), .B(n1330), .Y(mult_x_1_n310) );
  INVXL U1042 ( .A(n1126), .Y(mult_x_1_n318) );
  NAND2XL U1043 ( .A(n617), .B(n616), .Y(n619) );
  INVXL U1044 ( .A(n619), .Y(n618) );
  AOI21XL U1045 ( .A0(n620), .A1(mult_x_1_n318), .B0(n618), .Y(mult_x_1_n311)
         );
  NAND2XL U1046 ( .A(n620), .B(n619), .Y(mult_x_1_n85) );
  XNOR2XL U1047 ( .A(n621), .B(n1301), .Y(PRODUCT[12]) );
  XNOR2X1 U1048 ( .A(n648), .B(A[6]), .Y(n624) );
  XNOR2X1 U1049 ( .A(n648), .B(A[7]), .Y(n694) );
  OAI22X1 U1050 ( .A0(n979), .A1(n624), .B0(n694), .B1(n1089), .Y(n688) );
  NOR2BX1 U1051 ( .AN(n1090), .B(n1010), .Y(n633) );
  OAI22X1 U1052 ( .A0(n987), .A1(n627), .B0(n93), .B1(n683), .Y(n702) );
  XNOR2X1 U1053 ( .A(n648), .B(A[4]), .Y(n656) );
  ADDHXL U1054 ( .A(n641), .B(n640), .CO(n635), .S(n666) );
  NOR2XL U1055 ( .A(n1205), .B(n1214), .Y(n679) );
  XNOR2X1 U1056 ( .A(n648), .B(n650), .Y(n643) );
  XNOR2X1 U1057 ( .A(n648), .B(n642), .Y(n649) );
  XNOR2X1 U1058 ( .A(n648), .B(n980), .Y(n657) );
  OAI22X1 U1059 ( .A0(n979), .A1(n649), .B0(n657), .B1(n1089), .Y(n661) );
  OAI22X1 U1060 ( .A0(n56), .A1(n651), .B0(n93), .B1(n659), .Y(n660) );
  OAI22XL U1061 ( .A0(n56), .A1(n653), .B0(n93), .B1(n652), .Y(n654) );
  OAI21XL U1062 ( .A0(n1243), .A1(n1240), .B0(n1241), .Y(n1238) );
  CMPR22X1 U1063 ( .A(n661), .B(n660), .CO(n663), .S(n655) );
  CMPR32X1 U1064 ( .A(n668), .B(n667), .C(n666), .CO(n674), .S(n673) );
  CMPR32X1 U1065 ( .A(n671), .B(n670), .C(n669), .CO(n672), .S(n664) );
  OAI21XL U1066 ( .A0(n1235), .A1(n1232), .B0(n1233), .Y(n1204) );
  NAND2XL U1067 ( .A(n677), .B(n676), .Y(n1206) );
  OAI21XL U1068 ( .A0(n1205), .A1(n1215), .B0(n1206), .Y(n678) );
  AOI21X1 U1069 ( .A0(n679), .A1(n1204), .B0(n678), .Y(n744) );
  OAI22XL U1070 ( .A0(n979), .A1(n694), .B0(n693), .B1(n1089), .Y(n698) );
  CMPR32X1 U1071 ( .A(n699), .B(n698), .C(n697), .CO(n722), .S(n708) );
  CMPR32X1 U1072 ( .A(n708), .B(n707), .C(n706), .CO(n714), .S(n713) );
  CMPR32X1 U1073 ( .A(n711), .B(n710), .C(n709), .CO(n712), .S(n677) );
  OR2X2 U1074 ( .A(n713), .B(n712), .Y(n1187) );
  NAND2XL U1075 ( .A(n713), .B(n712), .Y(n1186) );
  INVXL U1076 ( .A(n1186), .Y(n745) );
  NAND2XL U1077 ( .A(n715), .B(n714), .Y(n746) );
  INVXL U1078 ( .A(n746), .Y(n716) );
  AOI21X1 U1079 ( .A0(n747), .A1(n745), .B0(n716), .Y(n717) );
  CMPR32X1 U1080 ( .A(n724), .B(n723), .C(n722), .CO(n737), .S(n728) );
  CMPR32X1 U1081 ( .A(n738), .B(n737), .C(n736), .CO(n739), .S(n732) );
  INVXL U1082 ( .A(n1197), .Y(n741) );
  NAND2XL U1083 ( .A(n741), .B(n1199), .Y(n742) );
  INVXL U1084 ( .A(n744), .Y(n1189) );
  AOI21XL U1085 ( .A0(n1189), .A1(n1187), .B0(n745), .Y(n749) );
  XOR2X1 U1086 ( .A(n749), .B(n748), .Y(n1345) );
  ADDFHX1 U1087 ( .A(n752), .B(n751), .CI(n750), .CO(n302), .S(mult_x_1_n470)
         );
  CMPR32X1 U1088 ( .A(n755), .B(n754), .C(n753), .CO(n295), .S(n764) );
  CMPR32X1 U1089 ( .A(n758), .B(n757), .C(n756), .CO(n751), .S(n763) );
  ADDFHX1 U1090 ( .A(n761), .B(n760), .CI(n759), .CO(n762), .S(n143) );
  CMPR32X1 U1091 ( .A(n764), .B(n763), .C(n762), .CO(mult_x_1_n481), .S(
        mult_x_1_n482) );
  XNOR2XL U1092 ( .A(n107), .B(n899), .Y(n766) );
  NOR2XL U1093 ( .A(n8), .B(n766), .Y(n791) );
  OAI22XL U1094 ( .A0(n1018), .A1(n789), .B0(n1156), .B1(n767), .Y(n790) );
  XNOR2X1 U1095 ( .A(n972), .B(n940), .Y(n780) );
  XNOR2X1 U1096 ( .A(n648), .B(A[24]), .Y(n783) );
  OAI22X1 U1097 ( .A0(n979), .A1(n783), .B0(n772), .B1(n1089), .Y(n782) );
  XNOR2X1 U1098 ( .A(n775), .B(n774), .Y(n793) );
  OAI22X1 U1099 ( .A0(n56), .A1(n806), .B0(n93), .B1(n776), .Y(n809) );
  XNOR2X1 U1100 ( .A(n648), .B(n1159), .Y(n835) );
  XNOR2XL U1101 ( .A(n107), .B(n925), .Y(n784) );
  NOR2XL U1102 ( .A(n8), .B(n784), .Y(n833) );
  CMPR32X1 U1103 ( .A(n787), .B(n786), .C(n785), .CO(n801), .S(n821) );
  OAI22X1 U1104 ( .A0(n965), .A1(n826), .B0(n1010), .B1(n788), .Y(n831) );
  OAI22XL U1105 ( .A0(n1018), .A1(n828), .B0(n1016), .B1(n789), .Y(n829) );
  CMPR32X1 U1106 ( .A(n792), .B(n791), .C(n790), .CO(n787), .S(n818) );
  CMPR32X1 U1107 ( .A(n795), .B(n794), .C(n793), .CO(n785), .S(n817) );
  CMPR32X1 U1108 ( .A(n798), .B(n797), .C(n796), .CO(n142), .S(n799) );
  ADDFHX1 U1109 ( .A(n801), .B(n800), .CI(n799), .CO(mult_x_1_n507), .S(
        mult_x_1_n508) );
  CMPR32X1 U1110 ( .A(n804), .B(n803), .C(n802), .CO(n798), .S(n825) );
  ADDFHX1 U1111 ( .A(n810), .B(n809), .CI(n808), .CO(n816), .S(n849) );
  CMPR32X1 U1112 ( .A(n813), .B(n812), .C(n811), .CO(n814), .S(n848) );
  CMPR32X1 U1113 ( .A(n819), .B(n818), .C(n817), .CO(n820), .S(n851) );
  OAI22X1 U1114 ( .A0(n965), .A1(n857), .B0(n1010), .B1(n826), .Y(n862) );
  OAI22XL U1115 ( .A0(n1018), .A1(n859), .B0(n1016), .B1(n828), .Y(n860) );
  ADDHXL U1116 ( .A(n834), .B(n833), .CO(n811), .S(n843) );
  OAI22X1 U1117 ( .A0(n979), .A1(n866), .B0(n835), .B1(n976), .Y(n865) );
  XNOR2XL U1118 ( .A(n107), .B(A[7]), .Y(n836) );
  CMPR32X1 U1119 ( .A(n844), .B(n842), .C(n843), .CO(n845), .S(n879) );
  OAI22X1 U1120 ( .A0(n965), .A1(n888), .B0(n1010), .B1(n857), .Y(n893) );
  OAI22XL U1121 ( .A0(n1018), .A1(n890), .B0(n1016), .B1(n859), .Y(n891) );
  XNOR2XL U1122 ( .A(n107), .B(A[6]), .Y(n867) );
  NOR2XL U1123 ( .A(n8), .B(n867), .Y(n895) );
  CMPR32X1 U1124 ( .A(n875), .B(n874), .C(n873), .CO(n876), .S(n913) );
  OAI22X1 U1125 ( .A0(n965), .A1(n923), .B0(n1010), .B1(n888), .Y(n929) );
  OAI22XL U1126 ( .A0(n1018), .A1(n926), .B0(n1016), .B1(n890), .Y(n927) );
  ADDHXL U1127 ( .A(n896), .B(n895), .CO(n873), .S(n908) );
  OAI22X1 U1128 ( .A0(n935), .A1(n934), .B0(n897), .B1(n1089), .Y(n932) );
  XNOR2XL U1129 ( .A(n107), .B(n966), .Y(n898) );
  CMPR32X1 U1130 ( .A(n909), .B(n907), .C(n908), .CO(n910), .S(n954) );
  OAI22X1 U1131 ( .A0(n965), .A1(n964), .B0(n1010), .B1(n923), .Y(n971) );
  OAI22XL U1132 ( .A0(n1018), .A1(n968), .B0(n1016), .B1(n926), .Y(n969) );
  OAI22X1 U1133 ( .A0(n935), .A1(n977), .B0(n934), .B1(n1089), .Y(n975) );
  XNOR2XL U1134 ( .A(n107), .B(A[4]), .Y(n936) );
  CMPR32X1 U1135 ( .A(n950), .B(n949), .C(n948), .CO(n951), .S(n1000) );
  XNOR2XL U1136 ( .A(n1117), .B(A[7]), .Y(n1015) );
  OAI22XL U1137 ( .A0(n1018), .A1(n1015), .B0(n1016), .B1(n968), .Y(n1019) );
  XNOR2XL U1138 ( .A(n107), .B(n980), .Y(n981) );
  NOR2XL U1139 ( .A(n8), .B(n981), .Y(n1025) );
  OAI22X1 U1140 ( .A0(n5), .A1(n983), .B0(n9), .B1(n982), .Y(n1034) );
  CMPR32X1 U1141 ( .A(n996), .B(n995), .C(n994), .CO(n997), .S(n1041) );
  CMPR32X1 U1142 ( .A(n999), .B(n998), .C(n997), .CO(n1008), .S(n1045) );
  OAI22XL U1143 ( .A0(n1018), .A1(n1017), .B0(n1016), .B1(n1015), .Y(n1053) );
  ADDHXL U1144 ( .A(n1026), .B(n1025), .CO(n994), .S(n1036) );
  CMPR32X1 U1145 ( .A(n1031), .B(n1030), .C(n1029), .CO(n1067), .S(n1074) );
  ADDFX2 U1146 ( .A(n1034), .B(n1033), .CI(n1032), .CO(n1043), .S(n1066) );
  CMPR32X1 U1147 ( .A(n1037), .B(n1035), .C(n1036), .CO(n1038), .S(n1065) );
  CMPR32X1 U1148 ( .A(n1052), .B(n1051), .C(n1050), .CO(n1064), .S(n1060) );
  CMPR32X1 U1149 ( .A(n1058), .B(n1057), .C(n1056), .CO(n1062), .S(n1059) );
  CMPR32X1 U1150 ( .A(n1085), .B(n1084), .C(n1083), .CO(mult_x_1_n649), .S(
        mult_x_1_n650) );
  NAND2XL U1151 ( .A(n53), .B(n1099), .Y(mult_x_1_n83) );
  INVXL U1152 ( .A(n1099), .Y(mult_x_1_n298) );
  INVXL U1153 ( .A(n1100), .Y(n1102) );
  NAND2XL U1154 ( .A(n1105), .B(n1294), .Y(n1106) );
  CMPR32X1 U1155 ( .A(n1111), .B(n1110), .C(n1109), .CO(n1128), .S(n1107) );
  XNOR2X1 U1156 ( .A(n1117), .B(A[24]), .Y(n1138) );
  XNOR2X1 U1157 ( .A(n1161), .B(n1151), .Y(n1135) );
  CMPR32X1 U1158 ( .A(n1122), .B(n1121), .C(n1120), .CO(n1139), .S(n1111) );
  CMPR32X1 U1159 ( .A(n1125), .B(n1124), .C(n1123), .CO(n1129), .S(n1110) );
  CMPR32X1 U1160 ( .A(n1131), .B(n1130), .C(n1129), .CO(n1143), .S(n1127) );
  CMPR32X1 U1161 ( .A(n1134), .B(n1133), .C(n1132), .CO(n1146), .S(n1131) );
  XNOR2X1 U1162 ( .A(n1161), .B(n1159), .Y(n1147) );
  OAI22X1 U1163 ( .A0(n1018), .A1(n1138), .B0(n1156), .B1(n1153), .Y(n1166) );
  CMPR32X1 U1164 ( .A(n1141), .B(n1140), .C(n1139), .CO(n1144), .S(n1130) );
  CMPR32X1 U1165 ( .A(n1146), .B(n1145), .C(n1144), .CO(n1158), .S(n1142) );
  CMPR32X1 U1166 ( .A(n1150), .B(n1149), .C(n1148), .CO(n1179), .S(n1145) );
  OAI2BB1X1 U1167 ( .A0N(n1156), .A1N(n1018), .B0(n1154), .Y(n1164) );
  CMPR32X1 U1168 ( .A(n1166), .B(n1165), .C(n1164), .CO(n1181), .S(n1178) );
  OAI2BB1X1 U1169 ( .A0N(n1014), .A1N(n1170), .B0(n1169), .Y(n1171) );
  XOR3X2 U1170 ( .A(n1173), .B(n1172), .C(n1171), .Y(n1174) );
  CMPR32X1 U1171 ( .A(n1180), .B(n1179), .C(n1178), .CO(n1185), .S(n1157) );
  CMPR32X1 U1172 ( .A(n1183), .B(n1182), .C(n1181), .CO(n1175), .S(n1184) );
  OAI21XL U1173 ( .A0(n1266), .A1(n1193), .B0(n1192), .Y(n1196) );
  NOR2XL U1174 ( .A(n1200), .B(n1197), .Y(n1202) );
  OAI21XL U1175 ( .A0(n1200), .A1(n1199), .B0(n1198), .Y(n1201) );
  AOI21XL U1176 ( .A0(n1203), .A1(n1202), .B0(n1201), .Y(mult_x_1_n322) );
  OAI21XL U1177 ( .A0(n1217), .A1(n1214), .B0(n1215), .Y(n1209) );
  INVXL U1178 ( .A(n1205), .Y(n1207) );
  OAI21XL U1179 ( .A0(n1279), .A1(n1282), .B0(n1280), .Y(n1223) );
  OAI21XL U1180 ( .A0(n1266), .A1(n1211), .B0(n1210), .Y(n1213) );
  OAI21XL U1181 ( .A0(n1266), .A1(n1228), .B0(n1227), .Y(n1231) );
  OAI21XL U1182 ( .A0(n1256), .A1(n1275), .B0(n1276), .Y(n1257) );
  AOI21XL U1183 ( .A0(n1259), .A1(n1258), .B0(n1257), .Y(n1260) );
  OAI21XL U1184 ( .A0(n1262), .A1(n1261), .B0(n1260), .Y(n1263) );
  OAI21XL U1185 ( .A0(n1266), .A1(n1265), .B0(n1264), .Y(n1267) );
  XNOR2XL U1186 ( .A(n1267), .B(n1274), .Y(PRODUCT[40]) );
endmodule


module FFT2048_DW02_mult_2_stage_J1_2 ( A, B, TC, CLK, PRODUCT );
  input [25:0] A;
  input [16:0] B;
  output [42:0] PRODUCT;
  input TC, CLK;
  wire   n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, mult_x_1_n649, mult_x_1_n634, mult_x_1_n633,
         mult_x_1_n618, mult_x_1_n601, mult_x_1_n586, mult_x_1_n585,
         mult_x_1_n570, mult_x_1_n569, mult_x_1_n554, mult_x_1_n553,
         mult_x_1_n538, mult_x_1_n537, mult_x_1_n522, mult_x_1_n521,
         mult_x_1_n508, mult_x_1_n316, mult_x_1_n309, mult_x_1_n307,
         mult_x_1_n306, mult_x_1_n296, mult_x_1_n295, mult_x_1_n293,
         mult_x_1_n292, mult_x_1_n287, mult_x_1_n286, mult_x_1_n282,
         mult_x_1_n281, mult_x_1_n277, mult_x_1_n276, mult_x_1_n263,
         mult_x_1_n262, mult_x_1_n198, mult_x_1_n197, mult_x_1_n195,
         mult_x_1_n194, mult_x_1_n184, mult_x_1_n183, mult_x_1_n177,
         mult_x_1_n176, mult_x_1_n170, mult_x_1_n169, mult_x_1_n161,
         mult_x_1_n160, mult_x_1_n152, mult_x_1_n151, mult_x_1_n137,
         mult_x_1_n136, mult_x_1_n130, mult_x_1_n129, mult_x_1_n121,
         mult_x_1_n120, mult_x_1_n110, mult_x_1_n109, mult_x_1_n85,
         mult_x_1_n84, mult_x_1_n83, mult_x_1_n58, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305;

  DFFHQXL mult_x_1_clk_r_REG10_S1 ( .D(mult_x_1_n194), .CK(CLK), .Q(n1269) );
  DFFHQXL mult_x_1_clk_r_REG7_S1 ( .D(mult_x_1_n198), .CK(CLK), .Q(n1272) );
  DFFHQXL mult_x_1_clk_r_REG8_S1 ( .D(mult_x_1_n197), .CK(CLK), .Q(n1271) );
  DFFHQXL mult_x_1_clk_r_REG16_S1 ( .D(mult_x_1_n169), .CK(CLK), .Q(n1263) );
  DFFHQXL mult_x_1_clk_r_REG18_S1 ( .D(mult_x_1_n160), .CK(CLK), .Q(n1261) );
  DFFHQXL mult_x_1_clk_r_REG20_S1 ( .D(mult_x_1_n151), .CK(CLK), .Q(n1259) );
  DFFHQXL mult_x_1_clk_r_REG12_S1 ( .D(mult_x_1_n183), .CK(CLK), .Q(n1267) );
  DFFHQX4 mult_x_1_clk_r_REG40_S1 ( .D(mult_x_1_n649), .CK(CLK), .Q(n1305) );
  DFFHQX4 mult_x_1_clk_r_REG39_S1 ( .D(mult_x_1_n634), .CK(CLK), .Q(n1304) );
  DFFHQX4 mult_x_1_clk_r_REG38_S1 ( .D(mult_x_1_n633), .CK(CLK), .Q(n1303) );
  DFFHQX4 mult_x_1_clk_r_REG37_S1 ( .D(mult_x_1_n618), .CK(CLK), .Q(n1302) );
  DFFHQX4 mult_x_1_clk_r_REG34_S1 ( .D(mult_x_1_n601), .CK(CLK), .Q(n1301) );
  DFFHQX4 mult_x_1_clk_r_REG33_S1 ( .D(mult_x_1_n586), .CK(CLK), .Q(n1300) );
  DFFHQX4 mult_x_1_clk_r_REG30_S1 ( .D(mult_x_1_n569), .CK(CLK), .Q(n1297) );
  DFFHQX4 mult_x_1_clk_r_REG1_S1 ( .D(mult_x_1_n554), .CK(CLK), .Q(n1296) );
  DFFHQX4 mult_x_1_clk_r_REG0_S1 ( .D(mult_x_1_n553), .CK(CLK), .Q(n1295) );
  DFFHQX4 mult_x_1_clk_r_REG3_S1 ( .D(mult_x_1_n538), .CK(CLK), .Q(n1294) );
  DFFHQX4 mult_x_1_clk_r_REG56_S1 ( .D(mult_x_1_n309), .CK(CLK), .Q(n1288) );
  DFFHQX4 mult_x_1_clk_r_REG50_S1 ( .D(mult_x_1_n296), .CK(CLK), .Q(n1287) );
  DFFHQXL mult_x_1_clk_r_REG49_S1 ( .D(mult_x_1_n83), .CK(CLK), .Q(n1284) );
  DFFHQX4 mult_x_1_clk_r_REG51_S1 ( .D(mult_x_1_n295), .CK(CLK), .Q(n1283) );
  DFFHQX4 mult_x_1_clk_r_REG48_S1 ( .D(mult_x_1_n292), .CK(CLK), .Q(n1281) );
  DFFHQX4 mult_x_1_clk_r_REG45_S1 ( .D(mult_x_1_n287), .CK(CLK), .Q(n1280) );
  DFFHQX1 mult_x_1_clk_r_REG53_S1 ( .D(mult_x_1_n307), .CK(CLK), .Q(n1249) );
  DFFHQX1 mult_x_1_clk_r_REG54_S1 ( .D(mult_x_1_n306), .CK(CLK), .Q(n1248) );
  DFFHQXL clk_r_REG57_S1 ( .D(n1319), .CK(CLK), .Q(PRODUCT[12]) );
  DFFHQXL mult_x_1_clk_r_REG9_S1 ( .D(mult_x_1_n195), .CK(CLK), .Q(n1270) );
  DFFHQXL mult_x_1_clk_r_REG21_S1 ( .D(mult_x_1_n137), .CK(CLK), .Q(n1258) );
  DFFHQXL mult_x_1_clk_r_REG11_S1 ( .D(mult_x_1_n184), .CK(CLK), .Q(n1268) );
  DFFHQXL mult_x_1_clk_r_REG13_S1 ( .D(mult_x_1_n177), .CK(CLK), .Q(n1266) );
  DFFHQXL mult_x_1_clk_r_REG14_S1 ( .D(mult_x_1_n176), .CK(CLK), .Q(n1265) );
  DFFHQXL clk_r_REG60_S1 ( .D(n1321), .CK(CLK), .Q(PRODUCT[10]) );
  DFFHQXL clk_r_REG61_S1 ( .D(n1322), .CK(CLK), .Q(PRODUCT[9]) );
  DFFHQXL mult_x_1_clk_r_REG15_S1 ( .D(mult_x_1_n170), .CK(CLK), .Q(n1264) );
  DFFHQXL mult_x_1_clk_r_REG19_S1 ( .D(mult_x_1_n152), .CK(CLK), .Q(n1260) );
  DFFHQXL mult_x_1_clk_r_REG17_S1 ( .D(mult_x_1_n161), .CK(CLK), .Q(n1262) );
  DFFHQXL clk_r_REG59_S1 ( .D(n1320), .CK(CLK), .Q(PRODUCT[11]) );
  DFFHQXL clk_r_REG63_S1 ( .D(n1324), .CK(CLK), .Q(PRODUCT[7]) );
  DFFHQXL mult_x_1_clk_r_REG25_S1 ( .D(mult_x_1_n121), .CK(CLK), .Q(n1254) );
  DFFHQX1 mult_x_1_clk_r_REG35_S1 ( .D(mult_x_1_n263), .CK(CLK), .Q(n1274) );
  DFFHQXL clk_r_REG62_S1 ( .D(n1323), .CK(CLK), .Q(PRODUCT[8]) );
  DFFHQXL clk_r_REG64_S1 ( .D(n1325), .CK(CLK), .Q(PRODUCT[6]) );
  DFFHQXL clk_r_REG65_S1 ( .D(n1326), .CK(CLK), .Q(PRODUCT[5]) );
  DFFHQXL clk_r_REG66_S1 ( .D(n1327), .CK(CLK), .Q(PRODUCT[4]) );
  DFFHQXL clk_r_REG67_S1 ( .D(n1328), .CK(CLK), .Q(PRODUCT[3]) );
  DFFHQXL clk_r_REG68_S1 ( .D(n1329), .CK(CLK), .Q(PRODUCT[2]) );
  DFFHQXL clk_r_REG70_S1 ( .D(n1331), .CK(CLK), .Q(PRODUCT[0]) );
  DFFHQXL clk_r_REG69_S1 ( .D(n1330), .CK(CLK), .Q(PRODUCT[1]) );
  DFFHQXL mult_x_1_clk_r_REG52_S1 ( .D(mult_x_1_n84), .CK(CLK), .Q(n1285) );
  DFFHQXL mult_x_1_clk_r_REG23_S1 ( .D(mult_x_1_n130), .CK(CLK), .Q(n1256) );
  DFFHQXL mult_x_1_clk_r_REG24_S1 ( .D(mult_x_1_n129), .CK(CLK), .Q(n1255) );
  DFFHQXL mult_x_1_clk_r_REG26_S1 ( .D(mult_x_1_n120), .CK(CLK), .Q(n1253) );
  DFFHQXL mult_x_1_clk_r_REG27_S1 ( .D(mult_x_1_n110), .CK(CLK), .Q(n1252) );
  DFFHQXL mult_x_1_clk_r_REG28_S1 ( .D(mult_x_1_n109), .CK(CLK), .Q(n1251) );
  DFFHQXL mult_x_1_clk_r_REG29_S1 ( .D(mult_x_1_n58), .CK(CLK), .Q(n1250) );
  DFFHQXL mult_x_1_clk_r_REG58_S1 ( .D(mult_x_1_n316), .CK(CLK), .Q(n1289) );
  DFFHQXL mult_x_1_clk_r_REG22_S1 ( .D(mult_x_1_n136), .CK(CLK), .Q(n1257) );
  DFFHQX1 mult_x_1_clk_r_REG47_S1 ( .D(mult_x_1_n293), .CK(CLK), .Q(n1282) );
  DFFHQX2 mult_x_1_clk_r_REG36_S1 ( .D(mult_x_1_n262), .CK(CLK), .Q(n1273) );
  DFFHQXL mult_x_1_clk_r_REG55_S1 ( .D(mult_x_1_n85), .CK(CLK), .Q(n1286) );
  DFFHQX1 mult_x_1_clk_r_REG46_S1 ( .D(mult_x_1_n286), .CK(CLK), .Q(n1279) );
  DFFHQX1 mult_x_1_clk_r_REG42_S1 ( .D(mult_x_1_n276), .CK(CLK), .Q(n1275) );
  DFFHQX1 mult_x_1_clk_r_REG43_S1 ( .D(mult_x_1_n282), .CK(CLK), .Q(n1278) );
  DFFHQX2 mult_x_1_clk_r_REG44_S1 ( .D(mult_x_1_n281), .CK(CLK), .Q(n1277) );
  DFFHQX2 mult_x_1_clk_r_REG2_S1 ( .D(mult_x_1_n537), .CK(CLK), .Q(n1293) );
  DFFHQX2 mult_x_1_clk_r_REG4_S1 ( .D(mult_x_1_n521), .CK(CLK), .Q(n1291) );
  DFFHQX2 mult_x_1_clk_r_REG5_S1 ( .D(mult_x_1_n522), .CK(CLK), .Q(n1292) );
  DFFHQX2 mult_x_1_clk_r_REG32_S1 ( .D(mult_x_1_n585), .CK(CLK), .Q(n1299) );
  DFFHQX2 mult_x_1_clk_r_REG31_S1 ( .D(mult_x_1_n570), .CK(CLK), .Q(n1298) );
  DFFHQX2 mult_x_1_clk_r_REG6_S1 ( .D(mult_x_1_n508), .CK(CLK), .Q(n1290) );
  DFFHQX1 mult_x_1_clk_r_REG41_S1 ( .D(mult_x_1_n277), .CK(CLK), .Q(n1276) );
  ADDFHX1 U1 ( .A(n872), .B(n871), .CI(n870), .CO(n565), .S(mult_x_1_n508) );
  ADDFHX1 U2 ( .A(n563), .B(n562), .CI(n561), .CO(n520), .S(n564) );
  ADDFHX2 U3 ( .A(n499), .B(n498), .CI(n497), .CO(n516), .S(n562) );
  ADDFHX2 U4 ( .A(n742), .B(n741), .CI(n740), .CO(n715), .S(n747) );
  ADDFHX2 U5 ( .A(n894), .B(n893), .CI(n892), .CO(n871), .S(n895) );
  CMPR32X1 U6 ( .A(n992), .B(n991), .C(n990), .CO(n995), .S(n1037) );
  CMPR32X1 U7 ( .A(n957), .B(n956), .C(n955), .CO(n960), .S(n993) );
  CMPR32X1 U8 ( .A(n924), .B(n923), .C(n922), .CO(n927), .S(n958) );
  OAI21X2 U9 ( .A0(n81), .A1(n80), .B0(n79), .Y(n22) );
  ADDFHX1 U10 ( .A(n464), .B(n463), .CI(n462), .CO(n457), .S(n517) );
  ADDFHX1 U11 ( .A(n954), .B(n953), .CI(n952), .CO(n963), .S(n994) );
  ADDFHX2 U12 ( .A(n834), .B(n833), .CI(n832), .CO(n805), .S(n841) );
  CMPR32X1 U13 ( .A(n1036), .B(n1035), .C(n1034), .CO(n1039), .S(n1112) );
  ADDFX2 U14 ( .A(n1051), .B(n1050), .CI(n1049), .CO(n1120), .S(n1046) );
  CMPR32X1 U15 ( .A(n366), .B(n365), .C(n364), .CO(n409), .S(n404) );
  ADDFX2 U16 ( .A(n727), .B(n726), .CI(n725), .CO(n742), .S(n772) );
  ADDFHX1 U17 ( .A(n837), .B(n836), .CI(n835), .CO(n840), .S(n839) );
  NAND3BX1 U18 ( .AN(n857), .B(n856), .C(n7), .Y(n13) );
  CMPR32X1 U19 ( .A(n506), .B(n505), .C(n504), .CO(n515), .S(n874) );
  CMPR32X1 U20 ( .A(n477), .B(n476), .C(n475), .CO(n480), .S(n510) );
  ADDFHX1 U21 ( .A(n804), .B(n803), .CI(n802), .CO(n780), .S(n832) );
  ADDFHX1 U22 ( .A(n719), .B(n718), .CI(n717), .CO(n706), .S(n749) );
  ADDFHX1 U23 ( .A(n1005), .B(n1004), .CI(n1003), .CO(n989), .S(n1032) );
  CMPR32X1 U24 ( .A(n810), .B(n809), .C(n808), .CO(n802), .S(n837) );
  ADDHXL U25 ( .A(n795), .B(n794), .CO(n791), .S(n825) );
  CMPR32X1 U26 ( .A(n761), .B(n760), .C(n759), .CO(n756), .S(n810) );
  ADDFHX1 U27 ( .A(n233), .B(n232), .CI(n231), .CO(n850), .S(n244) );
  CMPR32X1 U28 ( .A(n798), .B(n797), .C(n796), .CO(n824), .S(n817) );
  ADDFX2 U29 ( .A(n688), .B(n687), .CI(n686), .CO(n695), .S(n726) );
  CMPR32X1 U30 ( .A(n650), .B(n649), .C(n648), .CO(n661), .S(n693) );
  CLKINVX3 U31 ( .A(n252), .Y(n500) );
  ADDFX2 U32 ( .A(n212), .B(n211), .CI(n210), .CO(n232), .S(n219) );
  CMPR32X1 U33 ( .A(n179), .B(n178), .C(n177), .CO(n185), .S(n184) );
  ADDFHX1 U34 ( .A(n222), .B(n221), .CI(n220), .CO(n223), .S(n186) );
  BUFX8 U35 ( .A(n470), .Y(n10) );
  CLKBUFX8 U36 ( .A(n1165), .Y(n1143) );
  BUFX4 U37 ( .A(n256), .Y(n6) );
  CLKBUFX8 U38 ( .A(n1061), .Y(n1140) );
  XNOR2X2 U39 ( .A(B[16]), .B(B[15]), .Y(n1013) );
  CMPR32X1 U40 ( .A(n176), .B(n175), .C(n174), .CO(n221), .S(n177) );
  CLKINVX4 U41 ( .A(n252), .Y(n976) );
  XOR2X1 U42 ( .A(B[11]), .B(B[10]), .Y(n58) );
  OAI22X1 U43 ( .A0(n1074), .A1(n156), .B0(n1072), .B1(n197), .Y(n199) );
  NAND2X1 U44 ( .A(n257), .B(n1165), .Y(n470) );
  CLKINVX3 U45 ( .A(B[13]), .Y(n739) );
  OAI22X1 U46 ( .A0(n11), .A1(n101), .B0(n168), .B1(n96), .Y(n18) );
  INVX4 U47 ( .A(B[11]), .Y(n252) );
  BUFX4 U48 ( .A(n100), .Y(n11) );
  INVX4 U49 ( .A(n106), .Y(n979) );
  NAND2X1 U50 ( .A(n98), .B(n381), .Y(n734) );
  INVX4 U51 ( .A(n530), .Y(n5) );
  OAI21XL U52 ( .A0(n1246), .A1(n452), .B0(n451), .Y(n455) );
  XOR2X1 U53 ( .A(n486), .B(n485), .Y(PRODUCT[30]) );
  XOR2X1 U54 ( .A(n586), .B(n585), .Y(PRODUCT[27]) );
  XOR2X1 U55 ( .A(n66), .B(n59), .Y(PRODUCT[24]) );
  XOR2X1 U56 ( .A(n1246), .B(n522), .Y(PRODUCT[29]) );
  XNOR2X1 U57 ( .A(n596), .B(n595), .Y(PRODUCT[26]) );
  OAI21XL U58 ( .A0(n1089), .A1(n591), .B0(n590), .Y(n596) );
  OAI21XL U59 ( .A0(n608), .A1(n1089), .B0(n607), .Y(n66) );
  INVXL U60 ( .A(n598), .Y(n589) );
  AOI21X1 U61 ( .A0(n569), .A1(n93), .B0(n92), .Y(n43) );
  NAND2X1 U62 ( .A(n1301), .B(n1300), .Y(n614) );
  AOI21X2 U63 ( .A0(n279), .A1(n612), .B0(n65), .Y(n598) );
  OAI21XL U64 ( .A0(n1089), .A1(n568), .B0(n598), .Y(n602) );
  NAND3BX2 U65 ( .AN(n42), .B(n40), .C(n1282), .Y(n39) );
  XOR2XL U66 ( .A(n579), .B(n578), .Y(PRODUCT[28]) );
  XNOR2XL U67 ( .A(n5), .B(A[6]), .Y(n97) );
  XNOR2XL U68 ( .A(B[3]), .B(A[6]), .Y(n162) );
  XNOR2XL U69 ( .A(B[3]), .B(A[9]), .Y(n241) );
  XNOR2XL U70 ( .A(n979), .B(A[9]), .Y(n766) );
  XNOR2XL U71 ( .A(B[16]), .B(A[7]), .Y(n909) );
  XNOR2XL U72 ( .A(B[3]), .B(A[17]), .Y(n1019) );
  XNOR2XL U73 ( .A(B[3]), .B(A[16]), .Y(n674) );
  XNOR2XL U74 ( .A(B[3]), .B(A[13]), .Y(n696) );
  XNOR2XL U75 ( .A(B[16]), .B(A[16]), .Y(n324) );
  XNOR2XL U76 ( .A(n979), .B(A[24]), .Y(n429) );
  XNOR2XL U77 ( .A(n976), .B(A[25]), .Y(n253) );
  XNOR2XL U78 ( .A(n979), .B(A[21]), .Y(n537) );
  BUFX4 U79 ( .A(n155), .Y(n1072) );
  XNOR2XL U80 ( .A(n1001), .B(A[21]), .Y(n322) );
  XNOR2XL U81 ( .A(n5), .B(A[1]), .Y(n118) );
  ADDFX2 U82 ( .A(n813), .B(n812), .CI(n811), .CO(n822), .S(n831) );
  XOR2X1 U83 ( .A(n31), .B(n693), .Y(n741) );
  AOI21XL U84 ( .A0(n856), .A1(n7), .B0(n8), .Y(n91) );
  XOR2XL U85 ( .A(n1194), .B(n1193), .Y(n1325) );
  AOI21XL U86 ( .A0(n1086), .A1(n843), .B0(n842), .Y(mult_x_1_n296) );
  XOR2X1 U87 ( .A(n869), .B(n868), .Y(n1322) );
  NAND2XL U88 ( .A(n1086), .B(n1085), .Y(mult_x_1_n83) );
  NOR2X1 U89 ( .A(n806), .B(n805), .Y(mult_x_1_n292) );
  XNOR2X1 U90 ( .A(n1183), .B(n1182), .Y(n1323) );
  ADDFHX2 U91 ( .A(n773), .B(n772), .CI(n771), .CO(n748), .S(n779) );
  ADDFHX2 U92 ( .A(n1120), .B(n1119), .CI(n1118), .CO(n1128), .S(n1079) );
  INVXL U93 ( .A(n73), .Y(n14) );
  ADDFHX1 U94 ( .A(n825), .B(n824), .CI(n823), .CO(n820), .S(n848) );
  NAND2BXL U95 ( .AN(n651), .B(n9), .Y(n48) );
  NOR2X1 U96 ( .A(n1162), .B(n324), .Y(n363) );
  NOR2X1 U97 ( .A(n1162), .B(n632), .Y(n657) );
  OAI2BB1XL U98 ( .A0N(n6), .A1N(n1140), .B0(n1139), .Y(n1145) );
  NOR2X1 U99 ( .A(n1162), .B(n1137), .Y(n1146) );
  NOR2X1 U100 ( .A(n1162), .B(n1141), .Y(n1160) );
  NOR2X1 U101 ( .A(n1162), .B(n378), .Y(n400) );
  OAI2BB1X1 U102 ( .A0N(n173), .A1N(n18), .B0(n16), .Y(n178) );
  NOR2X1 U103 ( .A(n149), .B(n148), .Y(n1190) );
  NOR2X1 U104 ( .A(n1013), .B(n909), .Y(n938) );
  NOR2X1 U105 ( .A(n1013), .B(n532), .Y(n542) );
  NAND2X1 U106 ( .A(n415), .B(n1266), .Y(n416) );
  AND2X1 U107 ( .A(n349), .B(n1262), .Y(n350) );
  NOR2X1 U108 ( .A(n592), .B(n587), .Y(n566) );
  NAND2X1 U109 ( .A(n711), .B(n1278), .Y(n712) );
  NAND2X1 U110 ( .A(n628), .B(n1276), .Y(n629) );
  INVX1 U111 ( .A(n605), .Y(n615) );
  NAND2X1 U112 ( .A(n1292), .B(n1293), .Y(n583) );
  XOR2X1 U113 ( .A(n864), .B(n863), .Y(n1321) );
  NAND2XL U114 ( .A(n806), .B(n805), .Y(mult_x_1_n293) );
  ADDFHX1 U115 ( .A(n749), .B(n748), .CI(n747), .CO(n743), .S(n775) );
  INVX1 U116 ( .A(n854), .Y(n1092) );
  CLKINVX3 U117 ( .A(n32), .Y(n1086) );
  NOR2X2 U118 ( .A(n841), .B(n840), .Y(n32) );
  ADDFHX1 U119 ( .A(n1129), .B(n1128), .CI(n1127), .CO(n1130), .S(
        mult_x_1_n618) );
  ADDFHX1 U120 ( .A(n1114), .B(n1113), .CI(n1112), .CO(n1041), .S(n1124) );
  ADDFHX1 U121 ( .A(n1105), .B(n1104), .CI(n1103), .CO(n1123), .S(n1118) );
  NAND2BXL U122 ( .AN(n689), .B(n9), .Y(n23) );
  NOR2X1 U123 ( .A(n1162), .B(n323), .Y(n338) );
  NOR2X1 U124 ( .A(n1162), .B(n259), .Y(n298) );
  INVXL U125 ( .A(n38), .Y(n36) );
  AND2XL U126 ( .A(n228), .B(n90), .Y(n818) );
  NOR2X1 U127 ( .A(n1162), .B(n261), .Y(n307) );
  INVXL U128 ( .A(n201), .Y(n15) );
  NOR2X1 U129 ( .A(n1162), .B(n355), .Y(n384) );
  ADDFHX1 U130 ( .A(n1054), .B(n1053), .CI(n1052), .CO(n1117), .S(n1044) );
  NOR2X1 U131 ( .A(n1162), .B(n251), .Y(n269) );
  NOR2X1 U132 ( .A(n1162), .B(n271), .Y(n1135) );
  NAND2XL U133 ( .A(n71), .B(n70), .Y(n69) );
  NAND2X1 U134 ( .A(n149), .B(n148), .Y(n1191) );
  OR2X2 U135 ( .A(n138), .B(n137), .Y(n136) );
  XNOR2XL U136 ( .A(B[16]), .B(A[21]), .Y(n271) );
  XNOR2XL U137 ( .A(B[16]), .B(A[24]), .Y(n1161) );
  XNOR2X1 U138 ( .A(n321), .B(n320), .Y(PRODUCT[35]) );
  XNOR2X1 U139 ( .A(n1198), .B(n1197), .Y(PRODUCT[38]) );
  XNOR2X1 U140 ( .A(n1179), .B(n1178), .Y(PRODUCT[37]) );
  XNOR2X1 U141 ( .A(n296), .B(n295), .Y(PRODUCT[36]) );
  XNOR2X1 U142 ( .A(n1211), .B(n1210), .Y(PRODUCT[39]) );
  XNOR2X2 U143 ( .A(n455), .B(n454), .Y(PRODUCT[31]) );
  NAND2X1 U144 ( .A(n94), .B(n96), .Y(n100) );
  OAI22X1 U145 ( .A0(n1011), .A1(n736), .B0(n723), .B1(n1084), .Y(n760) );
  NOR2X1 U146 ( .A(n1235), .B(n292), .Y(n1200) );
  CLKINVX3 U147 ( .A(B[1]), .Y(n530) );
  XNOR2X1 U148 ( .A(n778), .B(n777), .Y(PRODUCT[16]) );
  INVX1 U149 ( .A(n1087), .Y(n93) );
  NAND2X1 U150 ( .A(n521), .B(n1272), .Y(n522) );
  INVX1 U151 ( .A(n1261), .Y(n349) );
  NAND3X1 U152 ( .A(n13), .B(n12), .C(n858), .Y(n855) );
  NAND2X1 U153 ( .A(n1090), .B(n854), .Y(n250) );
  NAND2XL U154 ( .A(n744), .B(n743), .Y(mult_x_1_n282) );
  ADDFHX2 U155 ( .A(n716), .B(n715), .CI(n714), .CO(n708), .S(n744) );
  ADDFHX2 U156 ( .A(n1048), .B(n1047), .CI(n1046), .CO(n1080), .S(n1082) );
  NAND2X1 U157 ( .A(n249), .B(n248), .Y(n854) );
  INVXL U158 ( .A(mult_x_1_n307), .Y(n843) );
  ADDFHX2 U159 ( .A(n781), .B(n780), .CI(n779), .CO(n774), .S(n806) );
  XNOR2X1 U160 ( .A(n1189), .B(n1188), .Y(n1324) );
  INVX1 U161 ( .A(n861), .Y(n7) );
  INVX1 U162 ( .A(n862), .Y(n8) );
  INVXL U163 ( .A(n852), .Y(n89) );
  INVXL U164 ( .A(n1083), .Y(n21) );
  NAND2X1 U165 ( .A(n839), .B(n838), .Y(mult_x_1_n307) );
  ADDFHX2 U166 ( .A(n1123), .B(n1122), .CI(n1121), .CO(n1125), .S(n1127) );
  INVXL U167 ( .A(n694), .Y(n29) );
  ADDFHX2 U168 ( .A(n406), .B(n405), .CI(n404), .CO(n408), .S(n444) );
  OR2XL U169 ( .A(n1170), .B(n1169), .Y(n1172) );
  ADDFHX1 U170 ( .A(n828), .B(n827), .CI(n826), .CO(n847), .S(n849) );
  ADDFHX1 U171 ( .A(n989), .B(n988), .CI(n987), .CO(n998), .S(n1038) );
  NAND2BXL U172 ( .AN(n663), .B(n53), .Y(n52) );
  NAND2XL U173 ( .A(n663), .B(n55), .Y(n51) );
  ADDFHX1 U174 ( .A(n701), .B(n700), .CI(n699), .CO(n694), .S(n751) );
  OAI2BB1XL U175 ( .A0N(n35), .A1N(n731), .B0(n33), .Y(n725) );
  NAND2BXL U176 ( .AN(n732), .B(n36), .Y(n35) );
  INVXL U177 ( .A(n34), .Y(n33) );
  INVXL U178 ( .A(n695), .Y(n30) );
  OR2X2 U179 ( .A(n184), .B(n183), .Y(n1180) );
  ADDFHX1 U180 ( .A(n512), .B(n511), .CI(n510), .CO(n498), .S(n559) );
  INVXL U181 ( .A(n217), .Y(n74) );
  ADDFHX1 U182 ( .A(n437), .B(n436), .CI(n435), .CO(n421), .S(n479) );
  ADDFHX1 U183 ( .A(n672), .B(n671), .CI(n670), .CO(n1051), .S(n680) );
  ADDFHX1 U184 ( .A(n200), .B(n199), .CI(n198), .CO(n216), .S(n222) );
  ADDFHX1 U185 ( .A(n1099), .B(n1098), .CI(n1097), .CO(n1033), .S(n1107) );
  ADDFHX1 U186 ( .A(n1096), .B(n1095), .CI(n1094), .CO(n1108), .S(n1116) );
  INVXL U187 ( .A(n85), .Y(n84) );
  XNOR2X1 U188 ( .A(n17), .B(n173), .Y(n180) );
  XNOR2X1 U189 ( .A(n172), .B(n18), .Y(n17) );
  INVXL U190 ( .A(n193), .Y(n71) );
  INVX1 U191 ( .A(n1074), .Y(n9) );
  NAND2BXL U192 ( .AN(n651), .B(n25), .Y(n24) );
  INVXL U193 ( .A(n55), .Y(n53) );
  OAI2BB1XL U194 ( .A0N(n381), .A1N(n1024), .B0(n380), .Y(n398) );
  INVXL U195 ( .A(n1072), .Y(n25) );
  AND2XL U196 ( .A(n1224), .B(n1223), .Y(n1330) );
  OR2XL U197 ( .A(n1222), .B(n1221), .Y(n1224) );
  NAND2BXL U198 ( .AN(A[0]), .B(n979), .Y(n105) );
  INVX1 U199 ( .A(B[3]), .Y(n426) );
  XOR2X1 U200 ( .A(B[2]), .B(B[3]), .Y(n99) );
  INVX2 U201 ( .A(B[5]), .Y(n106) );
  OR2XL U202 ( .A(n1235), .B(n1241), .Y(n1245) );
  NAND2X1 U203 ( .A(B[1]), .B(n940), .Y(n119) );
  AND2X2 U204 ( .A(n577), .B(n576), .Y(n578) );
  AND2X2 U205 ( .A(n584), .B(n583), .Y(n585) );
  NAND2XL U206 ( .A(n375), .B(n1264), .Y(n376) );
  INVXL U207 ( .A(n618), .Y(n92) );
  AND2X2 U208 ( .A(n484), .B(n1270), .Y(n485) );
  INVXL U209 ( .A(A[10]), .Y(n50) );
  INVXL U210 ( .A(A[14]), .Y(n56) );
  INVXL U211 ( .A(A[13]), .Y(n57) );
  INVXL U212 ( .A(A[8]), .Y(n27) );
  INVXL U213 ( .A(A[6]), .Y(n77) );
  INVXL U214 ( .A(A[0]), .Y(n86) );
  NOR2X1 U215 ( .A(n1295), .B(n1294), .Y(n592) );
  BUFX8 U216 ( .A(n493), .Y(n1074) );
  XOR2X1 U217 ( .A(B[8]), .B(B[9]), .Y(n154) );
  OAI21XL U218 ( .A0(n1072), .A1(n49), .B0(n48), .Y(n663) );
  XOR2X1 U219 ( .A(n732), .B(n38), .Y(n37) );
  AOI21X2 U220 ( .A0(n285), .A1(n569), .B0(n284), .Y(n483) );
  NOR2X1 U221 ( .A(n1300), .B(n1301), .Y(n605) );
  NAND2X1 U222 ( .A(n603), .B(n279), .Y(n568) );
  OAI22X1 U223 ( .A0(n1016), .A1(n252), .B0(n877), .B1(n190), .Y(n90) );
  NAND3X1 U224 ( .A(n855), .B(n1090), .C(n1093), .Y(n88) );
  XNOR2X1 U225 ( .A(n904), .B(A[2]), .Y(n196) );
  OAI2BB1X1 U226 ( .A0N(n83), .A1N(n201), .B0(n82), .Y(n233) );
  XNOR2X1 U227 ( .A(B[2]), .B(B[1]), .Y(n126) );
  NAND2X1 U228 ( .A(n225), .B(n226), .Y(n858) );
  NAND2BX1 U229 ( .AN(n857), .B(n8), .Y(n12) );
  OAI21X1 U230 ( .A0(n865), .A1(n189), .B0(n188), .Y(n856) );
  NOR2X1 U231 ( .A(n226), .B(n225), .Y(n857) );
  XOR3X2 U232 ( .A(n217), .B(n216), .C(n73), .Y(n61) );
  OAI21X1 U233 ( .A0(n14), .A1(n74), .B0(n72), .Y(n245) );
  XOR2X1 U234 ( .A(n15), .B(n75), .Y(n73) );
  OAI21XL U235 ( .A0(n173), .A1(n18), .B0(n172), .Y(n16) );
  OAI21XL U236 ( .A0(n1185), .A1(n1191), .B0(n1186), .Y(n152) );
  NOR2X1 U237 ( .A(n151), .B(n150), .Y(n1185) );
  XNOR2X4 U238 ( .A(B[6]), .B(B[5]), .Y(n96) );
  XNOR3X2 U239 ( .A(n21), .B(n22), .C(n1082), .Y(n709) );
  NAND2XL U240 ( .A(n20), .B(n19), .Y(mult_x_1_n649) );
  NAND2XL U241 ( .A(n22), .B(n1083), .Y(n19) );
  OAI21XL U242 ( .A0(n1083), .A1(n22), .B0(n1082), .Y(n20) );
  OAI21XL U243 ( .A0(n1072), .A1(n26), .B0(n23), .Y(n701) );
  OAI21XL U244 ( .A0(n1074), .A1(n26), .B0(n24), .Y(n646) );
  XOR2X1 U245 ( .A(n904), .B(n27), .Y(n26) );
  OAI21XL U246 ( .A0(n30), .A1(n29), .B0(n28), .Y(n707) );
  OAI21XL U247 ( .A0(n694), .A1(n695), .B0(n693), .Y(n28) );
  XOR2X1 U248 ( .A(n695), .B(n694), .Y(n31) );
  AND2XL U249 ( .A(n732), .B(n38), .Y(n34) );
  XOR2X1 U250 ( .A(n731), .B(n37), .Y(n783) );
  OAI22X1 U251 ( .A0(n10), .A1(n691), .B0(n1143), .B1(n690), .Y(n38) );
  NAND3X2 U252 ( .A(n39), .B(n622), .C(n278), .Y(n45) );
  AOI21X1 U253 ( .A0(n39), .A1(n622), .B0(n621), .Y(n630) );
  AOI21X1 U254 ( .A0(n39), .A1(n745), .B0(n710), .Y(n713) );
  XNOR2X1 U255 ( .A(n746), .B(n39), .Y(PRODUCT[17]) );
  NAND3BX4 U256 ( .AN(n1281), .B(n41), .C(n1288), .Y(n40) );
  CLKINVX3 U257 ( .A(n1283), .Y(n41) );
  NOR2X1 U258 ( .A(n1281), .B(n1287), .Y(n42) );
  NOR2X2 U259 ( .A(n623), .B(n1275), .Y(n278) );
  NOR2X2 U260 ( .A(n1305), .B(n1304), .Y(n623) );
  XOR2X1 U261 ( .A(n43), .B(n620), .Y(PRODUCT[22]) );
  NAND3BX4 U262 ( .AN(n46), .B(n45), .C(n44), .Y(n569) );
  NAND2X1 U263 ( .A(n278), .B(n621), .Y(n44) );
  XOR2X1 U264 ( .A(n351), .B(n350), .Y(PRODUCT[34]) );
  OAI21XL U265 ( .A0(n623), .A1(n1276), .B0(n624), .Y(n46) );
  OAI21X1 U266 ( .A0(n1280), .A1(n1277), .B0(n1278), .Y(n621) );
  XOR3X2 U267 ( .A(n707), .B(n706), .C(n705), .Y(n714) );
  OAI21XL U268 ( .A0(n1074), .A1(n49), .B0(n47), .Y(n1064) );
  OR2X2 U269 ( .A(n1073), .B(n1072), .Y(n47) );
  XOR2X1 U270 ( .A(n904), .B(n50), .Y(n49) );
  OAI2BB1X1 U271 ( .A0N(n52), .A1N(n662), .B0(n51), .Y(n1045) );
  XOR2X1 U272 ( .A(n662), .B(n54), .Y(n660) );
  XOR2X1 U273 ( .A(n663), .B(n55), .Y(n54) );
  OAI22X1 U274 ( .A0(n1024), .A1(n652), .B0(n1022), .B1(n675), .Y(n55) );
  XNOR2X1 U275 ( .A(n106), .B(n56), .Y(n675) );
  XNOR2X1 U276 ( .A(n106), .B(n57), .Y(n652) );
  NAND2X4 U277 ( .A(n58), .B(n193), .Y(n1016) );
  XNOR2X4 U278 ( .A(B[10]), .B(B[9]), .Y(n193) );
  NAND2X1 U279 ( .A(n1305), .B(n1304), .Y(n624) );
  XOR2X1 U280 ( .A(n1285), .B(n844), .Y(PRODUCT[14]) );
  INVX1 U281 ( .A(n1288), .Y(n844) );
  NOR2X1 U282 ( .A(n1291), .B(n1290), .Y(n575) );
  XNOR2X1 U283 ( .A(B[8]), .B(B[7]), .Y(n155) );
  INVX4 U284 ( .A(n569), .Y(n1089) );
  OAI21X1 U285 ( .A0(n582), .A1(n62), .B0(n63), .Y(n586) );
  BUFX3 U286 ( .A(n1089), .Y(n62) );
  INVXL U287 ( .A(n1239), .Y(n291) );
  NAND2X1 U288 ( .A(n99), .B(n126), .Y(n242) );
  BUFX3 U289 ( .A(n242), .Y(n1020) );
  BUFX3 U290 ( .A(n381), .Y(n1022) );
  INVXL U291 ( .A(n1234), .Y(n292) );
  OAI21X2 U292 ( .A0(n618), .A1(n1273), .B0(n1274), .Y(n612) );
  INVXL U293 ( .A(n1233), .Y(n1205) );
  CLKBUFX8 U294 ( .A(B[9]), .Y(n904) );
  XOR2X1 U295 ( .A(B[6]), .B(B[7]), .Y(n94) );
  XNOR2XL U296 ( .A(n5), .B(A[16]), .Y(n634) );
  XNOR2XL U297 ( .A(n500), .B(A[24]), .Y(n266) );
  XNOR2XL U298 ( .A(n904), .B(A[7]), .Y(n689) );
  XNOR2XL U299 ( .A(n904), .B(A[24]), .Y(n331) );
  XNOR2XL U300 ( .A(n904), .B(A[23]), .Y(n354) );
  XNOR2XL U301 ( .A(n1132), .B(A[17]), .Y(n356) );
  XNOR2XL U302 ( .A(n1132), .B(A[16]), .Y(n389) );
  XNOR2XL U303 ( .A(n904), .B(A[22]), .Y(n390) );
  XNOR2XL U304 ( .A(n1142), .B(A[14]), .Y(n430) );
  NAND2XL U305 ( .A(n1177), .B(n1256), .Y(n1178) );
  NAND2XL U306 ( .A(n319), .B(n1260), .Y(n320) );
  CLKINVX3 U307 ( .A(n685), .Y(n1132) );
  XNOR2X1 U308 ( .A(n1142), .B(A[3]), .Y(n633) );
  XNOR2XL U309 ( .A(n976), .B(A[7]), .Y(n637) );
  BUFX3 U310 ( .A(n734), .Y(n1024) );
  XNOR2XL U311 ( .A(n1132), .B(A[21]), .Y(n258) );
  XNOR2XL U312 ( .A(n1132), .B(A[20]), .Y(n264) );
  XNOR2XL U313 ( .A(n500), .B(A[21]), .Y(n357) );
  XNOR2XL U314 ( .A(n1132), .B(A[24]), .Y(n1144) );
  INVXL U315 ( .A(n1138), .Y(n1139) );
  XNOR2XL U316 ( .A(n1132), .B(A[23]), .Y(n1133) );
  NOR2X1 U317 ( .A(n224), .B(n223), .Y(n861) );
  OAI22XL U318 ( .A0(n1020), .A1(n113), .B0(n1018), .B1(n103), .Y(n112) );
  OAI22XL U319 ( .A0(n1020), .A1(n132), .B0(n1018), .B1(n113), .Y(n142) );
  NAND2X1 U320 ( .A(n224), .B(n223), .Y(n862) );
  OAI22XL U321 ( .A0(n10), .A1(n1144), .B0(n1143), .B1(n1163), .Y(n1168) );
  INVXL U322 ( .A(n1262), .Y(n316) );
  NAND2XL U323 ( .A(n349), .B(n319), .Y(n290) );
  INVXL U324 ( .A(n1257), .Y(n1174) );
  INVXL U325 ( .A(n1259), .Y(n319) );
  NOR2XL U326 ( .A(n290), .B(n1263), .Y(n1234) );
  NOR2XL U327 ( .A(n1233), .B(n1251), .Y(n1238) );
  NOR2X1 U328 ( .A(n570), .B(n64), .Y(n63) );
  INVX1 U329 ( .A(n1279), .Y(n745) );
  NAND2BXL U330 ( .AN(A[0]), .B(n904), .Y(n163) );
  XNOR2XL U331 ( .A(B[3]), .B(A[10]), .Y(n765) );
  XNOR2XL U332 ( .A(n964), .B(A[6]), .Y(n786) );
  XNOR2XL U333 ( .A(n964), .B(A[7]), .Y(n785) );
  XNOR2XL U334 ( .A(n904), .B(A[5]), .Y(n762) );
  XNOR2XL U335 ( .A(n904), .B(A[6]), .Y(n728) );
  XNOR2XL U336 ( .A(B[3]), .B(A[11]), .Y(n764) );
  XNOR2XL U337 ( .A(n904), .B(A[0]), .Y(n156) );
  XNOR2XL U338 ( .A(n904), .B(A[1]), .Y(n197) );
  NOR2X1 U339 ( .A(n193), .B(n86), .Y(n85) );
  OAI22XL U340 ( .A0(n1074), .A1(n197), .B0(n1072), .B1(n196), .Y(n201) );
  NAND2BXL U341 ( .AN(A[0]), .B(n976), .Y(n190) );
  OAI22XL U342 ( .A0(n1011), .A1(n194), .B0(n229), .B1(n1084), .Y(n228) );
  XNOR2XL U343 ( .A(n904), .B(A[3]), .Y(n227) );
  XNOR2XL U344 ( .A(n904), .B(A[4]), .Y(n763) );
  XNOR2XL U345 ( .A(n5), .B(A[22]), .Y(n941) );
  XNOR2XL U346 ( .A(n5), .B(A[19]), .Y(n1010) );
  XNOR2XL U347 ( .A(n976), .B(A[10]), .Y(n1014) );
  XNOR2XL U348 ( .A(n5), .B(A[17]), .Y(n655) );
  XNOR2XL U349 ( .A(n5), .B(A[18]), .Y(n676) );
  XNOR2XL U350 ( .A(n976), .B(A[9]), .Y(n1015) );
  XNOR2XL U351 ( .A(B[3]), .B(A[12]), .Y(n730) );
  OAI22X1 U352 ( .A0(n10), .A1(n685), .B0(n1143), .B1(n684), .Y(n721) );
  NAND2BXL U353 ( .AN(A[0]), .B(n1142), .Y(n684) );
  XNOR2XL U354 ( .A(n1132), .B(A[18]), .Y(n332) );
  XNOR2XL U355 ( .A(n979), .B(A[25]), .Y(n379) );
  XNOR2XL U356 ( .A(n964), .B(A[23]), .Y(n395) );
  XNOR2XL U357 ( .A(n500), .B(A[19]), .Y(n397) );
  XNOR2XL U358 ( .A(B[3]), .B(A[25]), .Y(n427) );
  XNOR2XL U359 ( .A(n904), .B(A[21]), .Y(n424) );
  XNOR2XL U360 ( .A(n904), .B(A[20]), .Y(n432) );
  XNOR2XL U361 ( .A(n964), .B(A[2]), .Y(n167) );
  CLKINVX2 U362 ( .A(B[7]), .Y(n325) );
  XNOR2XL U363 ( .A(B[3]), .B(A[5]), .Y(n157) );
  XNOR2XL U364 ( .A(n964), .B(A[1]), .Y(n168) );
  INVXL U365 ( .A(n1236), .Y(n1204) );
  NAND2XL U366 ( .A(n1200), .B(n1205), .Y(n1208) );
  INVXL U367 ( .A(n1251), .Y(n1209) );
  NAND2XL U368 ( .A(n1234), .B(n1238), .Y(n1241) );
  NAND2XL U369 ( .A(n1202), .B(n1254), .Y(n1197) );
  OAI22XL U370 ( .A0(n242), .A1(n206), .B0(n1018), .B1(n209), .Y(n210) );
  NOR2BXL U371 ( .AN(A[0]), .B(n1143), .Y(n761) );
  OAI22XL U372 ( .A0(n1020), .A1(n209), .B0(n1018), .B1(n241), .Y(n234) );
  OAI22XL U373 ( .A0(n11), .A1(n207), .B0(n96), .B1(n240), .Y(n236) );
  OAI22X1 U374 ( .A0(n1016), .A1(n208), .B0(n877), .B1(n230), .Y(n235) );
  XNOR2XL U375 ( .A(n964), .B(A[20]), .Y(n495) );
  XNOR2XL U376 ( .A(n904), .B(A[17]), .Y(n541) );
  OAI22XL U377 ( .A0(n1024), .A1(n488), .B0(n1022), .B1(n429), .Y(n474) );
  OAI22X1 U378 ( .A0(n10), .A1(n471), .B0(n1143), .B1(n430), .Y(n473) );
  OAI22X1 U379 ( .A0(n1020), .A1(n502), .B0(n1018), .B1(n427), .Y(n490) );
  XNOR2XL U380 ( .A(n904), .B(A[19]), .Y(n492) );
  XNOR2XL U381 ( .A(n904), .B(A[18]), .Y(n529) );
  XNOR2XL U382 ( .A(n904), .B(A[16]), .Y(n905) );
  OAI22XL U383 ( .A0(n1011), .A1(n908), .B0(n544), .B1(n940), .Y(n907) );
  XNOR2XL U384 ( .A(n964), .B(A[18]), .Y(n898) );
  XNOR2XL U385 ( .A(n904), .B(A[15]), .Y(n937) );
  XNOR2XL U386 ( .A(n964), .B(A[17]), .Y(n931) );
  XNOR2X1 U387 ( .A(n1142), .B(A[8]), .Y(n966) );
  XNOR2XL U388 ( .A(n964), .B(A[16]), .Y(n965) );
  XNOR2XL U389 ( .A(n964), .B(A[15]), .Y(n999) );
  XNOR2X1 U390 ( .A(n1142), .B(A[6]), .Y(n1057) );
  XNOR2XL U391 ( .A(n964), .B(A[14]), .Y(n1055) );
  XNOR2X1 U392 ( .A(n1142), .B(A[5]), .Y(n1058) );
  OAI22XL U393 ( .A0(n10), .A1(n690), .B0(n1143), .B1(n635), .Y(n686) );
  NOR2BXL U394 ( .AN(A[0]), .B(n1013), .Y(n688) );
  XNOR2X1 U395 ( .A(n1142), .B(A[4]), .Y(n665) );
  OAI22XL U396 ( .A0(n1016), .A1(n304), .B0(n877), .B1(n266), .Y(n308) );
  OAI2BB1XL U397 ( .A0N(n1072), .A1N(n1074), .B0(n263), .Y(n305) );
  INVXL U398 ( .A(n262), .Y(n263) );
  XNOR2XL U399 ( .A(n500), .B(A[22]), .Y(n352) );
  CMPR32X1 U400 ( .A(n363), .B(n362), .C(n361), .CO(n337), .S(n405) );
  OAI2BB1XL U401 ( .A0N(n96), .A1N(n11), .B0(n327), .Y(n361) );
  INVXL U402 ( .A(n326), .Y(n327) );
  INVXL U403 ( .A(n362), .Y(n385) );
  OAI22XL U404 ( .A0(n1074), .A1(n390), .B0(n1072), .B1(n354), .Y(n386) );
  OAI22XL U405 ( .A0(n1016), .A1(n391), .B0(n877), .B1(n357), .Y(n382) );
  OAI22XL U406 ( .A0(n10), .A1(n389), .B0(n1143), .B1(n356), .Y(n383) );
  CMPR32X1 U407 ( .A(n491), .B(n490), .C(n489), .CO(n466), .S(n514) );
  OAI2BB1XL U408 ( .A0N(n1018), .A1N(n1020), .B0(n428), .Y(n489) );
  NOR2X1 U409 ( .A(n1013), .B(n425), .Y(n491) );
  INVXL U410 ( .A(n427), .Y(n428) );
  XNOR2XL U411 ( .A(B[3]), .B(A[4]), .Y(n103) );
  OAI22XL U412 ( .A0(n10), .A1(n258), .B0(n1143), .B1(n270), .Y(n274) );
  OAI22XL U413 ( .A0(n10), .A1(n270), .B0(n1143), .B1(n1133), .Y(n1136) );
  INVXL U414 ( .A(n1147), .Y(n1134) );
  OAI22XL U415 ( .A0(n11), .A1(n698), .B0(n96), .B1(n641), .Y(n702) );
  OAI22XL U416 ( .A0(n1024), .A1(n720), .B0(n1022), .B1(n640), .Y(n704) );
  OAI22X1 U417 ( .A0(n697), .A1(n1016), .B0(n193), .B1(n76), .Y(n703) );
  CMPR32X1 U418 ( .A(n644), .B(n643), .C(n642), .CO(n682), .S(n718) );
  OAI22X1 U419 ( .A0(n10), .A1(n635), .B0(n1143), .B1(n633), .Y(n644) );
  OAI22XL U420 ( .A0(n11), .A1(n641), .B0(n96), .B1(n654), .Y(n647) );
  OAI22XL U421 ( .A0(n734), .A1(n640), .B0(n1022), .B1(n652), .Y(n648) );
  OAI22X1 U422 ( .A0(n637), .A1(n193), .B0(n1016), .B1(n76), .Y(n650) );
  OAI22XL U423 ( .A0(n119), .A1(n131), .B0(n130), .B1(n1084), .Y(n144) );
  OAI22XL U424 ( .A0(n242), .A1(n133), .B0(n1018), .B1(n132), .Y(n143) );
  NOR2BXL U425 ( .AN(A[0]), .B(n1022), .Y(n145) );
  INVXL U426 ( .A(n1163), .Y(n1164) );
  NOR2XL U427 ( .A(n1162), .B(n1161), .Y(n1167) );
  INVXL U428 ( .A(n1168), .Y(n1159) );
  NAND2XL U429 ( .A(n853), .B(n852), .Y(n1091) );
  OAI22XL U430 ( .A0(n1011), .A1(A[0]), .B0(n118), .B1(n1084), .Y(n1222) );
  NAND2XL U431 ( .A(n120), .B(n1011), .Y(n1221) );
  NAND2BXL U432 ( .AN(A[0]), .B(n5), .Y(n120) );
  NAND2XL U433 ( .A(n1222), .B(n1221), .Y(n1223) );
  NOR2XL U434 ( .A(n129), .B(n128), .Y(n1212) );
  AOI21XL U435 ( .A0(n1218), .A1(n1219), .B0(n123), .Y(n1215) );
  INVXL U436 ( .A(n1217), .Y(n123) );
  NAND2XL U437 ( .A(n129), .B(n128), .Y(n1213) );
  NAND2XL U438 ( .A(n138), .B(n137), .Y(n1225) );
  AOI21XL U439 ( .A0(n1226), .A1(n136), .B0(n139), .Y(n1231) );
  INVXL U440 ( .A(n1225), .Y(n139) );
  INVXL U441 ( .A(n1184), .Y(n1193) );
  NAND2XL U442 ( .A(n1199), .B(n1202), .Y(n1233) );
  NOR2XL U443 ( .A(n1257), .B(n1255), .Y(n1199) );
  NAND2XL U444 ( .A(n566), .B(n281), .Y(n283) );
  NOR2XL U445 ( .A(n581), .B(n567), .Y(n572) );
  INVXL U446 ( .A(n566), .Y(n581) );
  INVXL U447 ( .A(n568), .Y(n597) );
  NOR2X1 U448 ( .A(n1296), .B(n1297), .Y(n587) );
  NOR2X1 U449 ( .A(n1302), .B(n1303), .Y(n1087) );
  INVXL U450 ( .A(n1258), .Y(n1173) );
  NAND2XL U451 ( .A(n1200), .B(n1174), .Y(n1176) );
  INVXL U452 ( .A(n1255), .Y(n1177) );
  AOI21XL U453 ( .A0(n316), .A1(n319), .B0(n288), .Y(n289) );
  INVXL U454 ( .A(n1260), .Y(n288) );
  AOI21XL U455 ( .A0(n1203), .A1(n1202), .B0(n1201), .Y(n1236) );
  INVXL U456 ( .A(n1254), .Y(n1201) );
  NAND2XL U457 ( .A(n1200), .B(n1199), .Y(n1196) );
  INVXL U458 ( .A(n1253), .Y(n1202) );
  INVXL U459 ( .A(n1263), .Y(n375) );
  INVXL U460 ( .A(n1268), .Y(n412) );
  NAND2XL U461 ( .A(n449), .B(n453), .Y(n414) );
  INVXL U462 ( .A(n1265), .Y(n415) );
  INVXL U463 ( .A(n1267), .Y(n453) );
  AOI21XL U464 ( .A0(n589), .A1(n572), .B0(n571), .Y(n573) );
  OAI21XL U465 ( .A0(n580), .A1(n567), .B0(n583), .Y(n571) );
  NAND2XL U466 ( .A(n572), .B(n597), .Y(n574) );
  NAND2XL U467 ( .A(n1290), .B(n1291), .Y(n576) );
  NAND2XL U468 ( .A(n597), .B(n566), .Y(n582) );
  INVXL U469 ( .A(n567), .Y(n584) );
  AOI21XL U470 ( .A0(n589), .A1(n600), .B0(n588), .Y(n590) );
  INVXL U471 ( .A(n599), .Y(n588) );
  NAND2XL U472 ( .A(n597), .B(n600), .Y(n591) );
  INVXL U473 ( .A(n592), .Y(n594) );
  OAI21X1 U474 ( .A0(n609), .A1(n614), .B0(n610), .Y(n65) );
  INVXL U475 ( .A(n587), .Y(n600) );
  INVXL U476 ( .A(n609), .Y(n611) );
  NAND2X1 U477 ( .A(n1302), .B(n1303), .Y(n618) );
  INVXL U478 ( .A(n1280), .Y(n710) );
  XNOR2XL U479 ( .A(n5), .B(A[14]), .Y(n723) );
  XNOR2XL U480 ( .A(n976), .B(A[0]), .Y(n208) );
  XNOR2XL U481 ( .A(n964), .B(A[4]), .Y(n207) );
  XNOR2XL U482 ( .A(n976), .B(A[1]), .Y(n230) );
  CLKINVX3 U483 ( .A(B[15]), .Y(n685) );
  NOR2BXL U484 ( .AN(n202), .B(n86), .Y(n70) );
  XNOR2XL U485 ( .A(n5), .B(A[25]), .Y(n531) );
  XNOR2XL U486 ( .A(n5), .B(A[24]), .Y(n544) );
  XNOR2XL U487 ( .A(n5), .B(A[23]), .Y(n908) );
  XNOR2XL U488 ( .A(n976), .B(A[14]), .Y(n876) );
  XNOR2XL U489 ( .A(n979), .B(A[20]), .Y(n879) );
  XNOR2XL U490 ( .A(n5), .B(A[20]), .Y(n1009) );
  XNOR2XL U491 ( .A(n5), .B(A[15]), .Y(n683) );
  XNOR2XL U492 ( .A(n1132), .B(A[19]), .Y(n303) );
  XNOR2XL U493 ( .A(n500), .B(A[23]), .Y(n304) );
  XNOR2XL U494 ( .A(n964), .B(A[25]), .Y(n326) );
  XNOR2XL U495 ( .A(n500), .B(A[20]), .Y(n391) );
  NOR2XL U496 ( .A(n1013), .B(n393), .Y(n437) );
  OAI22X1 U497 ( .A0(n1140), .A1(n433), .B0(n6), .B1(n394), .Y(n436) );
  NAND2XL U498 ( .A(n1174), .B(n1258), .Y(n295) );
  OAI21XL U499 ( .A0(n1246), .A1(n348), .B0(n347), .Y(n351) );
  OAI21XL U500 ( .A0(n483), .A1(n1271), .B0(n1272), .Y(n486) );
  OAI21XL U501 ( .A0(n574), .A1(n1089), .B0(n573), .Y(n579) );
  NAND2X1 U502 ( .A(n619), .B(n1274), .Y(n620) );
  XNOR2X1 U503 ( .A(n617), .B(n616), .Y(PRODUCT[23]) );
  OAI21XL U504 ( .A0(n844), .A1(n1283), .B0(n1287), .Y(n778) );
  XOR2X1 U505 ( .A(n1289), .B(n1286), .Y(PRODUCT[13]) );
  INVXL U506 ( .A(n904), .Y(n164) );
  CMPR32X1 U507 ( .A(n215), .B(n214), .C(n213), .CO(n218), .S(n220) );
  OAI22XL U508 ( .A0(n242), .A1(n162), .B0(n1018), .B1(n206), .Y(n215) );
  OAI22XL U509 ( .A0(n1024), .A1(n243), .B0(n1022), .B1(n767), .Y(n799) );
  OAI22XL U510 ( .A0(n242), .A1(n241), .B0(n1018), .B1(n765), .Y(n800) );
  NAND2BXL U511 ( .AN(A[0]), .B(n1001), .Y(n738) );
  OAI22XL U512 ( .A0(n1024), .A1(n767), .B0(n1022), .B1(n766), .Y(n814) );
  OAI22XL U513 ( .A0(n1074), .A1(n763), .B0(n1072), .B1(n762), .Y(n816) );
  OAI22XL U514 ( .A0(n1020), .A1(n765), .B0(n1018), .B1(n764), .Y(n815) );
  XNOR2XL U515 ( .A(n1132), .B(A[22]), .Y(n270) );
  OAI22XL U516 ( .A0(n1016), .A1(n790), .B0(n193), .B1(n789), .Y(n811) );
  OAI22XL U517 ( .A0(n11), .A1(n786), .B0(n96), .B1(n785), .Y(n813) );
  CMPR32X1 U518 ( .A(n793), .B(n792), .C(n791), .CO(n782), .S(n821) );
  OAI22XL U519 ( .A0(n734), .A1(n766), .B0(n1022), .B1(n733), .Y(n793) );
  OAI22XL U520 ( .A0(n11), .A1(n785), .B0(n96), .B1(n735), .Y(n792) );
  OAI22XL U521 ( .A0(n1140), .A1(n724), .B0(n6), .B1(n692), .Y(n731) );
  ADDFX2 U522 ( .A(n770), .B(n769), .CI(n768), .CO(n784), .S(n808) );
  OAI22XL U523 ( .A0(n1020), .A1(n764), .B0(n1018), .B1(n730), .Y(n768) );
  OAI22XL U524 ( .A0(n1016), .A1(n789), .B0(n193), .B1(n729), .Y(n769) );
  OAI22XL U525 ( .A0(n1024), .A1(n158), .B0(n1022), .B1(n205), .Y(n198) );
  ADDFX2 U526 ( .A(n239), .B(n238), .CI(n237), .CO(n827), .S(n246) );
  OAI22X1 U527 ( .A0(n1074), .A1(n196), .B0(n1072), .B1(n227), .Y(n238) );
  OAI22XL U528 ( .A0(n1024), .A1(n204), .B0(n1022), .B1(n243), .Y(n239) );
  NAND3X1 U529 ( .A(n69), .B(n68), .C(n67), .Y(n75) );
  NAND2BXL U530 ( .AN(n202), .B(n86), .Y(n67) );
  NAND2BXL U531 ( .AN(n202), .B(n193), .Y(n68) );
  NAND2XL U532 ( .A(n202), .B(n85), .Y(n82) );
  NAND2BXL U533 ( .AN(n202), .B(n84), .Y(n83) );
  OAI22X1 U534 ( .A0(n1140), .A1(n487), .B0(n6), .B1(n433), .Y(n476) );
  INVXL U535 ( .A(n531), .Y(n503) );
  XNOR2XL U536 ( .A(n500), .B(A[15]), .Y(n535) );
  OAI22XL U537 ( .A0(n1074), .A1(n905), .B0(n1072), .B1(n541), .Y(n885) );
  ADDFX2 U538 ( .A(n882), .B(n881), .CI(n880), .CO(n888), .S(n923) );
  OAI22XL U539 ( .A0(n1024), .A1(n879), .B0(n1022), .B1(n537), .Y(n880) );
  OAI22XL U540 ( .A0(n1020), .A1(n878), .B0(n1018), .B1(n536), .Y(n881) );
  OAI22XL U541 ( .A0(n1016), .A1(n876), .B0(n877), .B1(n535), .Y(n882) );
  XNOR2XL U542 ( .A(n904), .B(A[14]), .Y(n971) );
  OAI22XL U543 ( .A0(n1011), .A1(n974), .B0(n941), .B1(n940), .Y(n973) );
  CMPR32X1 U544 ( .A(n915), .B(n914), .C(n913), .CO(n924), .S(n956) );
  OAI22XL U545 ( .A0(n1024), .A1(n912), .B0(n1022), .B1(n879), .Y(n913) );
  OAI22XL U546 ( .A0(n1020), .A1(n911), .B0(n1018), .B1(n878), .Y(n914) );
  OAI22XL U547 ( .A0(n1016), .A1(n910), .B0(n877), .B1(n876), .Y(n915) );
  OAI22XL U548 ( .A0(n1024), .A1(n945), .B0(n1022), .B1(n912), .Y(n946) );
  OAI22XL U549 ( .A0(n1020), .A1(n944), .B0(n1018), .B1(n911), .Y(n947) );
  OAI22XL U550 ( .A0(n1016), .A1(n943), .B0(n193), .B1(n910), .Y(n948) );
  OAI22XL U551 ( .A0(n1024), .A1(n980), .B0(n1022), .B1(n945), .Y(n981) );
  OAI22XL U552 ( .A0(n1020), .A1(n978), .B0(n1018), .B1(n944), .Y(n982) );
  OAI22XL U553 ( .A0(n1016), .A1(n977), .B0(n193), .B1(n943), .Y(n983) );
  OAI22XL U554 ( .A0(n1011), .A1(n676), .B0(n1010), .B1(n1084), .Y(n1078) );
  ADDFX2 U555 ( .A(n1027), .B(n1026), .CI(n1025), .CO(n1036), .S(n1110) );
  OAI22X1 U556 ( .A0(n1020), .A1(n1017), .B0(n1018), .B1(n978), .Y(n1026) );
  OAI22XL U557 ( .A0(n1020), .A1(n1019), .B0(n1018), .B1(n1017), .Y(n1069) );
  OAI22XL U558 ( .A0(n1015), .A1(n1016), .B0(n1014), .B1(n193), .Y(n1070) );
  XNOR2XL U559 ( .A(n1142), .B(A[2]), .Y(n635) );
  XNOR2XL U560 ( .A(n964), .B(A[10]), .Y(n641) );
  XOR2XL U561 ( .A(n976), .B(n77), .Y(n76) );
  XNOR2XL U562 ( .A(n979), .B(A[12]), .Y(n640) );
  XNOR2XL U563 ( .A(n904), .B(A[9]), .Y(n651) );
  XNOR2XL U564 ( .A(n964), .B(A[11]), .Y(n654) );
  OAI22XL U565 ( .A0(n1011), .A1(n634), .B0(n655), .B1(n1084), .Y(n658) );
  NAND2BXL U566 ( .AN(A[0]), .B(B[16]), .Y(n632) );
  CMPR32X1 U567 ( .A(n1067), .B(n1066), .C(n1065), .CO(n1105), .S(n1050) );
  OAI22XL U568 ( .A0(n1024), .A1(n675), .B0(n1022), .B1(n1023), .Y(n1065) );
  OAI22XL U569 ( .A0(n1020), .A1(n674), .B0(n1018), .B1(n1019), .Y(n1066) );
  OAI22XL U570 ( .A0(n1016), .A1(n673), .B0(n877), .B1(n1015), .Y(n1067) );
  OAI22XL U571 ( .A0(n11), .A1(n735), .B0(n96), .B1(n698), .Y(n753) );
  OAI22XL U572 ( .A0(n1020), .A1(n730), .B0(n1018), .B1(n696), .Y(n755) );
  OAI22XL U573 ( .A0(n1016), .A1(n729), .B0(n193), .B1(n697), .Y(n754) );
  OAI22XL U574 ( .A0(n734), .A1(n733), .B0(n1022), .B1(n720), .Y(n758) );
  OAI22XL U575 ( .A0(n1074), .A1(n354), .B0(n1072), .B1(n331), .Y(n360) );
  OAI22XL U576 ( .A0(n1140), .A1(n353), .B0(n6), .B1(n333), .Y(n358) );
  OAI22XL U577 ( .A0(n10), .A1(n356), .B0(n1143), .B1(n332), .Y(n359) );
  OAI22XL U578 ( .A0(n1074), .A1(n424), .B0(n1072), .B1(n390), .Y(n401) );
  OAI22XL U579 ( .A0(n11), .A1(n395), .B0(n96), .B1(n388), .Y(n403) );
  OAI22XL U580 ( .A0(n10), .A1(n396), .B0(n1143), .B1(n389), .Y(n402) );
  INVXL U581 ( .A(n379), .Y(n380) );
  ADDFX2 U582 ( .A(n440), .B(n439), .CI(n438), .CO(n461), .S(n478) );
  OAI22XL U583 ( .A0(n1016), .A1(n434), .B0(n877), .B1(n397), .Y(n438) );
  OAI22X1 U584 ( .A0(n10), .A1(n430), .B0(n1143), .B1(n396), .Y(n439) );
  ADDFX2 U585 ( .A(n423), .B(n422), .CI(n421), .CO(n442), .S(n464) );
  OAI22XL U586 ( .A0(n1016), .A1(n397), .B0(n877), .B1(n391), .Y(n423) );
  OAI22X1 U587 ( .A0(n1140), .A1(n394), .B0(n6), .B1(n392), .Y(n422) );
  OAI22XL U588 ( .A0(n1074), .A1(n432), .B0(n1072), .B1(n424), .Y(n467) );
  XNOR2X1 U589 ( .A(n5), .B(A[2]), .Y(n124) );
  XNOR2XL U590 ( .A(n5), .B(A[4]), .Y(n130) );
  XNOR2XL U591 ( .A(n5), .B(A[3]), .Y(n131) );
  ADDFX2 U592 ( .A(n171), .B(n170), .CI(n169), .CO(n213), .S(n179) );
  OAI22X1 U593 ( .A0(n1011), .A1(n166), .B0(n165), .B1(n1084), .Y(n170) );
  NOR2BXL U594 ( .AN(A[0]), .B(n1072), .Y(n171) );
  OAI22XL U595 ( .A0(n11), .A1(n168), .B0(n96), .B1(n167), .Y(n169) );
  NAND2BXL U596 ( .AN(A[0]), .B(n964), .Y(n95) );
  OAI22XL U597 ( .A0(n1024), .A1(n102), .B0(n1022), .B1(n159), .Y(n172) );
  OAI22XL U598 ( .A0(n1011), .A1(n104), .B0(n97), .B1(n1084), .Y(n108) );
  OAI22XL U599 ( .A0(n1024), .A1(n114), .B0(n1022), .B1(n102), .Y(n107) );
  NOR2BXL U600 ( .AN(A[0]), .B(n96), .Y(n109) );
  NAND2XL U601 ( .A(n1209), .B(n1252), .Y(n1210) );
  INVXL U602 ( .A(n1243), .Y(n1244) );
  ADDFX2 U603 ( .A(n831), .B(n830), .CI(n829), .CO(n836), .S(n846) );
  OAI2BB1XL U604 ( .A0N(n877), .A1N(n1016), .B0(n254), .Y(n267) );
  INVXL U605 ( .A(n253), .Y(n254) );
  ADDFX2 U606 ( .A(n784), .B(n783), .CI(n782), .CO(n771), .S(n834) );
  CMPR32X1 U607 ( .A(n528), .B(n527), .C(n526), .CO(n512), .S(n547) );
  OAI22XL U608 ( .A0(n11), .A1(n495), .B0(n96), .B1(n468), .Y(n528) );
  OAI22XL U609 ( .A0(n10), .A1(n496), .B0(n1143), .B1(n471), .Y(n526) );
  CMPR32X1 U610 ( .A(n554), .B(n553), .C(n552), .CO(n548), .S(n890) );
  OAI22XL U611 ( .A0(n1024), .A1(n537), .B0(n1022), .B1(n523), .Y(n554) );
  NOR2XL U612 ( .A(n1013), .B(n524), .Y(n553) );
  OAI22XL U613 ( .A0(n1074), .A1(n541), .B0(n1072), .B1(n529), .Y(n557) );
  INVXL U614 ( .A(n490), .Y(n504) );
  OR2XL U615 ( .A(n534), .B(n533), .Y(n507) );
  ADDFX2 U616 ( .A(n540), .B(n539), .CI(n538), .CO(n875), .S(n887) );
  OAI2BB1XL U617 ( .A0N(n1084), .A1N(n1011), .B0(n503), .Y(n538) );
  OAI22XL U618 ( .A0(n1020), .A1(n536), .B0(n1018), .B1(n502), .Y(n539) );
  OAI22XL U619 ( .A0(n1016), .A1(n535), .B0(n877), .B1(n501), .Y(n540) );
  OAI22XL U620 ( .A0(n1074), .A1(n937), .B0(n1072), .B1(n905), .Y(n918) );
  ADDFX2 U621 ( .A(n888), .B(n887), .CI(n886), .CO(n894), .S(n926) );
  CMPR32X1 U622 ( .A(n936), .B(n935), .C(n934), .CO(n921), .S(n953) );
  OAI22XL U623 ( .A0(n11), .A1(n931), .B0(n96), .B1(n898), .Y(n936) );
  CMPR32X1 U624 ( .A(n970), .B(n969), .C(n968), .CO(n954), .S(n988) );
  OAI22XL U625 ( .A0(n11), .A1(n965), .B0(n96), .B1(n931), .Y(n970) );
  OAI22X1 U626 ( .A0(n10), .A1(n966), .B0(n1143), .B1(n932), .Y(n969) );
  OAI22X2 U627 ( .A0(n10), .A1(n1057), .B0(n1143), .B1(n1000), .Y(n1098) );
  OAI22XL U628 ( .A0(n1061), .A1(n1060), .B0(n6), .B1(n1059), .Y(n1094) );
  OAI22XL U629 ( .A0(n1020), .A1(n638), .B0(n1018), .B1(n674), .Y(n670) );
  OAI22XL U630 ( .A0(n1140), .A1(n653), .B0(n6), .B1(n666), .Y(n662) );
  INVXL U631 ( .A(n268), .Y(n297) );
  OAI22XL U632 ( .A0(n10), .A1(n264), .B0(n1143), .B1(n258), .Y(n299) );
  OAI22XL U633 ( .A0(n1140), .A1(n265), .B0(n6), .B1(n260), .Y(n302) );
  OAI22XL U634 ( .A0(n1140), .A1(n333), .B0(n6), .B1(n322), .Y(n339) );
  OAI22XL U635 ( .A0(n1016), .A1(n357), .B0(n877), .B1(n352), .Y(n366) );
  ADDFX2 U636 ( .A(n461), .B(n460), .CI(n459), .CO(n441), .S(n518) );
  NOR2BXL U637 ( .AN(A[0]), .B(n1018), .Y(n121) );
  OAI22XL U638 ( .A0(n1011), .A1(n118), .B0(n124), .B1(n1084), .Y(n122) );
  OAI22XL U639 ( .A0(n1020), .A1(n426), .B0(n1018), .B1(n127), .Y(n128) );
  NAND2BXL U640 ( .AN(A[0]), .B(B[3]), .Y(n127) );
  OAI22XL U641 ( .A0(n10), .A1(n1133), .B0(n1143), .B1(n1144), .Y(n1153) );
  NAND2XL U642 ( .A(n122), .B(n121), .Y(n1217) );
  INVXL U643 ( .A(n1223), .Y(n1219) );
  NAND2XL U644 ( .A(n1157), .B(n1156), .Y(mult_x_1_n121) );
  NAND2XL U645 ( .A(n1187), .B(n1186), .Y(n1188) );
  XOR2X1 U646 ( .A(n860), .B(n91), .Y(n1320) );
  NAND2XL U647 ( .A(n60), .B(n867), .Y(n868) );
  INVXL U648 ( .A(n856), .Y(n864) );
  NAND2XL U649 ( .A(n1172), .B(n1171), .Y(mult_x_1_n58) );
  NAND2XL U650 ( .A(n1170), .B(n1169), .Y(n1171) );
  NOR2XL U651 ( .A(n1155), .B(n1154), .Y(mult_x_1_n109) );
  NAND2XL U652 ( .A(n1155), .B(n1154), .Y(mult_x_1_n110) );
  NOR2XL U653 ( .A(n1157), .B(n1156), .Y(mult_x_1_n120) );
  NOR2XL U654 ( .A(n1131), .B(n1130), .Y(mult_x_1_n262) );
  NAND2XL U655 ( .A(n1086), .B(n845), .Y(mult_x_1_n295) );
  NAND2X1 U656 ( .A(n1093), .B(n1092), .Y(n87) );
  INVX1 U657 ( .A(n706), .Y(n80) );
  NOR2XL U658 ( .A(n482), .B(n481), .Y(mult_x_1_n183) );
  NOR2BXL U659 ( .AN(A[0]), .B(n1084), .Y(n1331) );
  XNOR2XL U660 ( .A(n1220), .B(n1219), .Y(n1329) );
  NAND2XL U661 ( .A(n1218), .B(n1217), .Y(n1220) );
  XOR2XL U662 ( .A(n1216), .B(n1215), .Y(n1328) );
  NAND2XL U663 ( .A(n1214), .B(n1213), .Y(n1216) );
  INVXL U664 ( .A(n1212), .Y(n1214) );
  NAND2XL U665 ( .A(n136), .B(n1225), .Y(n1227) );
  NAND2XL U666 ( .A(n1230), .B(n1229), .Y(n1232) );
  INVXL U667 ( .A(n1228), .Y(n1230) );
  NAND2XL U668 ( .A(n1192), .B(n1191), .Y(n1194) );
  INVXL U669 ( .A(n1190), .Y(n1192) );
  NAND2XL U670 ( .A(n1180), .B(n1181), .Y(n1182) );
  AND2X1 U671 ( .A(n611), .B(n610), .Y(n59) );
  OR2X2 U672 ( .A(n186), .B(n185), .Y(n60) );
  CMPR22X1 U673 ( .A(n939), .B(n938), .CO(n916), .S(n950) );
  CMPR22X1 U674 ( .A(n1076), .B(n1075), .CO(n1028), .S(n1101) );
  OAI22X1 U675 ( .A0(n119), .A1(n195), .B0(n194), .B1(n1084), .Y(n202) );
  XOR2X1 U676 ( .A(n90), .B(n228), .Y(n237) );
  OAI22X1 U677 ( .A0(n493), .A1(n331), .B0(n1072), .B1(n262), .Y(n306) );
  CMPR22X1 U678 ( .A(n543), .B(n542), .CO(n556), .S(n884) );
  CMPR22X1 U679 ( .A(n117), .B(n116), .CO(n111), .S(n140) );
  CMPR22X1 U680 ( .A(n161), .B(n160), .CO(n174), .S(n182) );
  OAI22X1 U681 ( .A0(n11), .A1(n325), .B0(n96), .B1(n95), .Y(n160) );
  AOI21XL U682 ( .A0(n1206), .A1(n1205), .B0(n1204), .Y(n1207) );
  AOI21XL U683 ( .A0(n1206), .A1(n1199), .B0(n1203), .Y(n1195) );
  NOR2X1 U684 ( .A(n598), .B(n581), .Y(n64) );
  NOR2X2 U685 ( .A(n605), .B(n609), .Y(n279) );
  OAI21X1 U686 ( .A0(n73), .A1(n217), .B0(n216), .Y(n72) );
  BUFX2 U687 ( .A(n707), .Y(n78) );
  OAI21X1 U688 ( .A0(n706), .A1(n78), .B0(n705), .Y(n79) );
  INVX1 U689 ( .A(n78), .Y(n81) );
  NAND3X1 U690 ( .A(n88), .B(n87), .C(n1091), .Y(mult_x_1_n309) );
  NAND2BX1 U691 ( .AN(n853), .B(n89), .Y(n1093) );
  NAND2XL U692 ( .A(n151), .B(n150), .Y(n1186) );
  XOR2X2 U693 ( .A(n1089), .B(n1088), .Y(PRODUCT[21]) );
  XNOR2X2 U694 ( .A(B[14]), .B(B[13]), .Y(n1165) );
  XNOR2X1 U695 ( .A(n807), .B(n1284), .Y(PRODUCT[15]) );
  CMPR22X1 U696 ( .A(n1008), .B(n1007), .CO(n984), .S(n1029) );
  NOR2X1 U697 ( .A(n1013), .B(n975), .Y(n1007) );
  CMPR22X1 U698 ( .A(n679), .B(n678), .CO(n1062), .S(n668) );
  NOR2X1 U699 ( .A(n1013), .B(n656), .Y(n678) );
  OAI22X1 U700 ( .A0(n11), .A1(n167), .B0(n96), .B1(n203), .Y(n200) );
  OAI22X1 U701 ( .A0(n11), .A1(n203), .B0(n96), .B1(n207), .Y(n212) );
  INVX8 U702 ( .A(n325), .Y(n964) );
  AOI21XL U703 ( .A0(n1206), .A1(n1174), .B0(n1173), .Y(n1175) );
  NOR2XL U704 ( .A(n568), .B(n283), .Y(n285) );
  XNOR2X1 U705 ( .A(n964), .B(A[3]), .Y(n203) );
  XNOR2X1 U706 ( .A(n1001), .B(A[1]), .Y(n787) );
  XNOR2XL U707 ( .A(n5), .B(A[21]), .Y(n974) );
  XNOR2XL U708 ( .A(B[3]), .B(A[0]), .Y(n125) );
  INVX1 U709 ( .A(B[0]), .Y(n940) );
  XNOR2X1 U710 ( .A(n5), .B(A[7]), .Y(n166) );
  BUFX3 U711 ( .A(n940), .Y(n1084) );
  OAI22X1 U712 ( .A0(n119), .A1(n97), .B0(n166), .B1(n1084), .Y(n161) );
  XNOR2X1 U713 ( .A(n5), .B(A[5]), .Y(n104) );
  XOR2X1 U714 ( .A(B[4]), .B(B[5]), .Y(n98) );
  XNOR2X1 U715 ( .A(B[4]), .B(B[3]), .Y(n381) );
  XNOR2X1 U716 ( .A(n979), .B(A[1]), .Y(n114) );
  XNOR2X1 U717 ( .A(n979), .B(A[2]), .Y(n102) );
  OAI22X1 U718 ( .A0(n1020), .A1(n103), .B0(n1018), .B1(n157), .Y(n173) );
  XNOR2XL U719 ( .A(n964), .B(A[0]), .Y(n101) );
  XNOR2X1 U720 ( .A(n979), .B(A[3]), .Y(n159) );
  XNOR2X1 U721 ( .A(B[3]), .B(A[3]), .Y(n113) );
  OAI22X1 U722 ( .A0(n1011), .A1(n130), .B0(n104), .B1(n1084), .Y(n117) );
  OAI22X1 U723 ( .A0(n1024), .A1(n106), .B0(n1022), .B1(n105), .Y(n116) );
  CMPR32X1 U724 ( .A(n109), .B(n108), .C(n107), .CO(n181), .S(n110) );
  CMPR32X1 U725 ( .A(n112), .B(n111), .C(n110), .CO(n150), .S(n149) );
  XNOR2X1 U726 ( .A(B[3]), .B(A[2]), .Y(n132) );
  XNOR2XL U727 ( .A(n979), .B(A[0]), .Y(n115) );
  OAI22XL U728 ( .A0(n734), .A1(n115), .B0(n1022), .B1(n114), .Y(n141) );
  NOR2XL U729 ( .A(n1185), .B(n1190), .Y(n153) );
  OR2X2 U730 ( .A(n122), .B(n121), .Y(n1218) );
  BUFX3 U731 ( .A(n119), .Y(n1011) );
  OAI22X1 U732 ( .A0(n1011), .A1(n124), .B0(n131), .B1(n1084), .Y(n135) );
  XNOR2X1 U733 ( .A(B[3]), .B(A[1]), .Y(n133) );
  OAI22X1 U734 ( .A0(n1020), .A1(n125), .B0(n1018), .B1(n133), .Y(n134) );
  BUFX3 U735 ( .A(n126), .Y(n1018) );
  OAI21XL U736 ( .A0(n1215), .A1(n1212), .B0(n1213), .Y(n1226) );
  CMPR22X1 U737 ( .A(n135), .B(n134), .CO(n137), .S(n129) );
  CMPR32X1 U738 ( .A(n142), .B(n141), .C(n140), .CO(n148), .S(n147) );
  CMPR32X1 U739 ( .A(n145), .B(n144), .C(n143), .CO(n146), .S(n138) );
  NOR2XL U740 ( .A(n147), .B(n146), .Y(n1228) );
  NAND2XL U741 ( .A(n147), .B(n146), .Y(n1229) );
  OAI21XL U742 ( .A0(n1231), .A1(n1228), .B0(n1229), .Y(n1184) );
  AOI21XL U743 ( .A0(n153), .A1(n1184), .B0(n152), .Y(n865) );
  NAND2X2 U744 ( .A(n154), .B(n155), .Y(n493) );
  XNOR2X1 U745 ( .A(n979), .B(A[4]), .Y(n158) );
  XNOR2X1 U746 ( .A(n979), .B(A[5]), .Y(n205) );
  OAI22X1 U747 ( .A0(n1020), .A1(n157), .B0(n1018), .B1(n162), .Y(n176) );
  OAI22X2 U748 ( .A0(n1024), .A1(n159), .B0(n1022), .B1(n158), .Y(n175) );
  XNOR2X1 U749 ( .A(B[3]), .B(A[7]), .Y(n206) );
  XNOR2X1 U750 ( .A(n5), .B(A[8]), .Y(n165) );
  XNOR2X1 U751 ( .A(n5), .B(A[9]), .Y(n195) );
  OAI22X1 U752 ( .A0(n1011), .A1(n165), .B0(n195), .B1(n1084), .Y(n192) );
  OAI22X1 U753 ( .A0(n493), .A1(n164), .B0(n1072), .B1(n163), .Y(n191) );
  ADDFHX1 U754 ( .A(n182), .B(n181), .CI(n180), .CO(n183), .S(n151) );
  NAND2XL U755 ( .A(n60), .B(n1180), .Y(n189) );
  NAND2XL U756 ( .A(n184), .B(n183), .Y(n1181) );
  INVXL U757 ( .A(n1181), .Y(n866) );
  NAND2XL U758 ( .A(n186), .B(n185), .Y(n867) );
  INVXL U759 ( .A(n867), .Y(n187) );
  AOI21XL U760 ( .A0(n60), .A1(n866), .B0(n187), .Y(n188) );
  XNOR2X1 U761 ( .A(n979), .B(A[6]), .Y(n204) );
  XNOR2X1 U762 ( .A(n979), .B(A[7]), .Y(n243) );
  XNOR2X1 U763 ( .A(n5), .B(A[10]), .Y(n194) );
  XNOR2X1 U764 ( .A(n5), .B(A[11]), .Y(n229) );
  BUFX3 U765 ( .A(n193), .Y(n877) );
  CMPR22X1 U766 ( .A(n192), .B(n191), .CO(n217), .S(n214) );
  OAI22X2 U767 ( .A0(n1024), .A1(n205), .B0(n1022), .B1(n204), .Y(n211) );
  XNOR2X1 U768 ( .A(B[3]), .B(A[8]), .Y(n209) );
  XNOR2X1 U769 ( .A(n964), .B(A[5]), .Y(n240) );
  CMPR32X1 U770 ( .A(n219), .B(n218), .C(n61), .CO(n225), .S(n224) );
  OAI22XL U771 ( .A0(n1074), .A1(n227), .B0(n1072), .B1(n763), .Y(n819) );
  XNOR2X1 U772 ( .A(B[12]), .B(B[11]), .Y(n256) );
  NOR2BX1 U773 ( .AN(A[0]), .B(n6), .Y(n798) );
  XNOR2X1 U774 ( .A(n5), .B(A[12]), .Y(n737) );
  OAI22X2 U775 ( .A0(n1011), .A1(n229), .B0(n737), .B1(n1084), .Y(n797) );
  XNOR2X1 U776 ( .A(n976), .B(A[2]), .Y(n790) );
  OAI22XL U777 ( .A0(n1016), .A1(n230), .B0(n193), .B1(n790), .Y(n796) );
  ADDFHX1 U778 ( .A(n236), .B(n235), .CI(n234), .CO(n828), .S(n231) );
  OAI22XL U779 ( .A0(n11), .A1(n240), .B0(n96), .B1(n786), .Y(n801) );
  XNOR2X1 U780 ( .A(n979), .B(A[8]), .Y(n767) );
  CMPR32X1 U781 ( .A(n246), .B(n245), .C(n244), .CO(n248), .S(n226) );
  NOR2X1 U782 ( .A(n249), .B(n248), .Y(n247) );
  INVX1 U783 ( .A(n247), .Y(n1090) );
  XNOR2X1 U784 ( .A(n855), .B(n250), .Y(n1319) );
  BUFX3 U785 ( .A(n1013), .Y(n1162) );
  XNOR2X1 U786 ( .A(B[16]), .B(A[20]), .Y(n251) );
  OAI22X1 U787 ( .A0(n1016), .A1(n266), .B0(n877), .B1(n253), .Y(n268) );
  XOR2X1 U788 ( .A(B[12]), .B(B[13]), .Y(n255) );
  NAND2X2 U789 ( .A(n255), .B(n256), .Y(n1061) );
  XNOR2X1 U790 ( .A(n1001), .B(A[23]), .Y(n260) );
  XNOR2X1 U791 ( .A(n1001), .B(A[24]), .Y(n272) );
  OAI22XL U792 ( .A0(n1140), .A1(n260), .B0(n6), .B1(n272), .Y(n275) );
  XOR2X1 U793 ( .A(B[14]), .B(B[15]), .Y(n257) );
  XNOR2XL U794 ( .A(B[16]), .B(A[19]), .Y(n259) );
  XNOR2XL U795 ( .A(n1001), .B(A[22]), .Y(n265) );
  XNOR2X1 U796 ( .A(B[16]), .B(A[18]), .Y(n261) );
  XNOR2XL U797 ( .A(n904), .B(A[25]), .Y(n262) );
  OAI22XL U798 ( .A0(n10), .A1(n303), .B0(n1143), .B1(n264), .Y(n310) );
  OAI22XL U799 ( .A0(n1140), .A1(n322), .B0(n6), .B1(n265), .Y(n309) );
  CMPR32X1 U800 ( .A(n269), .B(n268), .C(n267), .CO(n1150), .S(n313) );
  CLKINVX8 U801 ( .A(n739), .Y(n1001) );
  XNOR2X1 U802 ( .A(n1001), .B(A[25]), .Y(n1138) );
  OAI22X1 U803 ( .A0(n1140), .A1(n272), .B0(n6), .B1(n1138), .Y(n1147) );
  CMPR32X1 U804 ( .A(n275), .B(n274), .C(n273), .CO(n1148), .S(n312) );
  NOR2XL U805 ( .A(n277), .B(n276), .Y(mult_x_1_n129) );
  NAND2XL U806 ( .A(n277), .B(n276), .Y(mult_x_1_n130) );
  NOR2XL U807 ( .A(n1087), .B(n1273), .Y(n603) );
  NOR2X2 U808 ( .A(n1298), .B(n1299), .Y(n609) );
  NOR2X1 U809 ( .A(n1292), .B(n1293), .Y(n567) );
  NOR2XL U810 ( .A(n567), .B(n575), .Y(n281) );
  NOR2X1 U811 ( .A(n1277), .B(n1279), .Y(n622) );
  NAND2XL U812 ( .A(n1298), .B(n1299), .Y(n610) );
  NAND2X1 U813 ( .A(n1296), .B(n1297), .Y(n599) );
  NAND2X1 U814 ( .A(n1294), .B(n1295), .Y(n593) );
  OAI21XL U815 ( .A0(n592), .A1(n599), .B0(n593), .Y(n570) );
  OAI21XL U816 ( .A0(n575), .A1(n583), .B0(n576), .Y(n280) );
  AOI21XL U817 ( .A0(n281), .A1(n570), .B0(n280), .Y(n282) );
  OAI21X1 U818 ( .A0(n598), .A1(n283), .B0(n282), .Y(n284) );
  BUFX3 U819 ( .A(n483), .Y(n1246) );
  NOR2XL U820 ( .A(n1271), .B(n1269), .Y(n449) );
  NOR2XL U821 ( .A(n1267), .B(n1265), .Y(n287) );
  NAND2XL U822 ( .A(n449), .B(n287), .Y(n1235) );
  INVXL U823 ( .A(n1200), .Y(n294) );
  OAI21XL U824 ( .A0(n1269), .A1(n1272), .B0(n1270), .Y(n450) );
  OAI21XL U825 ( .A0(n1265), .A1(n1268), .B0(n1266), .Y(n286) );
  AOI21X1 U826 ( .A0(n450), .A1(n287), .B0(n286), .Y(n1242) );
  OAI21XL U827 ( .A0(n290), .A1(n1264), .B0(n289), .Y(n1239) );
  OAI21XL U828 ( .A0(n1242), .A1(n292), .B0(n291), .Y(n1206) );
  INVXL U829 ( .A(n1206), .Y(n293) );
  OAI21XL U830 ( .A0(n1246), .A1(n294), .B0(n293), .Y(n296) );
  CMPR32X1 U831 ( .A(n299), .B(n298), .C(n297), .CO(n273), .S(n342) );
  CMPR32X1 U832 ( .A(n302), .B(n301), .C(n300), .CO(n311), .S(n341) );
  OAI22XL U833 ( .A0(n10), .A1(n332), .B0(n1143), .B1(n303), .Y(n336) );
  OAI22XL U834 ( .A0(n1016), .A1(n352), .B0(n877), .B1(n304), .Y(n335) );
  INVXL U835 ( .A(n306), .Y(n334) );
  CMPR32X1 U836 ( .A(n307), .B(n306), .C(n305), .CO(n301), .S(n329) );
  CMPR32X1 U837 ( .A(n310), .B(n309), .C(n308), .CO(n300), .S(n328) );
  CMPR32X1 U838 ( .A(n313), .B(n312), .C(n311), .CO(n277), .S(n314) );
  NOR2XL U839 ( .A(n315), .B(n314), .Y(mult_x_1_n136) );
  NAND2XL U840 ( .A(n315), .B(n314), .Y(mult_x_1_n137) );
  NOR2XL U841 ( .A(n1235), .B(n1263), .Y(n345) );
  NAND2XL U842 ( .A(n345), .B(n349), .Y(n318) );
  OAI21XL U843 ( .A0(n1242), .A1(n1263), .B0(n1264), .Y(n346) );
  AOI21XL U844 ( .A0(n346), .A1(n349), .B0(n316), .Y(n317) );
  OAI21XL U845 ( .A0(n1246), .A1(n318), .B0(n317), .Y(n321) );
  XNOR2X1 U846 ( .A(n1001), .B(A[20]), .Y(n333) );
  XNOR2X1 U847 ( .A(B[16]), .B(A[17]), .Y(n323) );
  XNOR2X1 U848 ( .A(n964), .B(A[24]), .Y(n388) );
  OAI22X1 U849 ( .A0(n11), .A1(n388), .B0(n96), .B1(n326), .Y(n362) );
  CMPR32X1 U850 ( .A(n330), .B(n329), .C(n328), .CO(n340), .S(n371) );
  XNOR2X1 U851 ( .A(n1001), .B(A[19]), .Y(n353) );
  CMPR32X1 U852 ( .A(n336), .B(n335), .C(n334), .CO(n330), .S(n368) );
  CMPR32X1 U853 ( .A(n339), .B(n338), .C(n337), .CO(n372), .S(n367) );
  CMPR32X1 U854 ( .A(n342), .B(n341), .C(n340), .CO(n315), .S(n343) );
  NOR2XL U855 ( .A(n344), .B(n343), .Y(mult_x_1_n151) );
  NAND2XL U856 ( .A(n344), .B(n343), .Y(mult_x_1_n152) );
  INVXL U857 ( .A(n345), .Y(n348) );
  INVXL U858 ( .A(n346), .Y(n347) );
  XNOR2X1 U859 ( .A(n1001), .B(A[18]), .Y(n392) );
  OAI22X1 U860 ( .A0(n1140), .A1(n392), .B0(n6), .B1(n353), .Y(n387) );
  XNOR2X1 U861 ( .A(B[16]), .B(A[15]), .Y(n355) );
  CMPR32X1 U862 ( .A(n360), .B(n359), .C(n358), .CO(n369), .S(n406) );
  CMPR32X1 U863 ( .A(n369), .B(n368), .C(n367), .CO(n370), .S(n407) );
  CMPR32X1 U864 ( .A(n372), .B(n371), .C(n370), .CO(n344), .S(n373) );
  NOR2XL U865 ( .A(n374), .B(n373), .Y(mult_x_1_n160) );
  NAND2XL U866 ( .A(n374), .B(n373), .Y(mult_x_1_n161) );
  OAI21XL U867 ( .A0(n1246), .A1(n1235), .B0(n1242), .Y(n377) );
  XNOR2X1 U868 ( .A(n377), .B(n376), .Y(PRODUCT[33]) );
  XNOR2X1 U869 ( .A(B[16]), .B(A[14]), .Y(n378) );
  OAI22X1 U870 ( .A0(n1024), .A1(n429), .B0(n1022), .B1(n379), .Y(n399) );
  CMPR32X1 U871 ( .A(n384), .B(n383), .C(n382), .CO(n364), .S(n419) );
  CMPR32X1 U872 ( .A(n387), .B(n386), .C(n385), .CO(n365), .S(n418) );
  XNOR2X1 U873 ( .A(n1132), .B(A[15]), .Y(n396) );
  XNOR2X1 U874 ( .A(n1001), .B(A[17]), .Y(n394) );
  XNOR2XL U875 ( .A(B[16]), .B(A[13]), .Y(n393) );
  XNOR2X1 U876 ( .A(n1001), .B(A[16]), .Y(n433) );
  INVXL U877 ( .A(n399), .Y(n435) );
  XNOR2XL U878 ( .A(n964), .B(A[22]), .Y(n431) );
  OAI22XL U879 ( .A0(n11), .A1(n431), .B0(n96), .B1(n395), .Y(n440) );
  INVX8 U880 ( .A(n685), .Y(n1142) );
  XNOR2XL U881 ( .A(n500), .B(A[18]), .Y(n434) );
  CMPR32X1 U882 ( .A(n400), .B(n399), .C(n398), .CO(n420), .S(n460) );
  CMPR32X1 U883 ( .A(n403), .B(n402), .C(n401), .CO(n443), .S(n459) );
  CMPR32X1 U884 ( .A(n409), .B(n408), .C(n407), .CO(n374), .S(n410) );
  NOR2XL U885 ( .A(n411), .B(n410), .Y(mult_x_1_n169) );
  NAND2XL U886 ( .A(n411), .B(n410), .Y(mult_x_1_n170) );
  AOI21XL U887 ( .A0(n450), .A1(n453), .B0(n412), .Y(n413) );
  OAI21XL U888 ( .A0(n1246), .A1(n414), .B0(n413), .Y(n417) );
  XNOR2X1 U889 ( .A(n417), .B(n416), .Y(PRODUCT[32]) );
  CMPR32X1 U890 ( .A(n420), .B(n419), .C(n418), .CO(n446), .S(n458) );
  XNOR2XL U891 ( .A(B[16]), .B(A[12]), .Y(n425) );
  XNOR2X1 U892 ( .A(B[3]), .B(A[24]), .Y(n502) );
  XNOR2X1 U893 ( .A(n979), .B(A[23]), .Y(n488) );
  XNOR2X1 U894 ( .A(n1142), .B(A[13]), .Y(n471) );
  XNOR2X1 U895 ( .A(n964), .B(A[21]), .Y(n468) );
  OAI22XL U896 ( .A0(n11), .A1(n468), .B0(n96), .B1(n431), .Y(n472) );
  OAI22XL U897 ( .A0(n493), .A1(n492), .B0(n1072), .B1(n432), .Y(n477) );
  XNOR2X1 U898 ( .A(n1001), .B(A[15]), .Y(n487) );
  XNOR2XL U899 ( .A(n500), .B(A[17]), .Y(n494) );
  OAI22XL U900 ( .A0(n1016), .A1(n494), .B0(n877), .B1(n434), .Y(n475) );
  CMPR32X1 U901 ( .A(n443), .B(n442), .C(n441), .CO(n445), .S(n456) );
  ADDFHX1 U902 ( .A(n446), .B(n445), .CI(n444), .CO(n411), .S(n447) );
  NOR2XL U903 ( .A(n448), .B(n447), .Y(mult_x_1_n176) );
  NAND2XL U904 ( .A(n448), .B(n447), .Y(mult_x_1_n177) );
  INVXL U905 ( .A(n449), .Y(n452) );
  INVXL U906 ( .A(n450), .Y(n451) );
  NAND2X1 U907 ( .A(n453), .B(n1268), .Y(n454) );
  ADDFHX1 U908 ( .A(n458), .B(n457), .CI(n456), .CO(n448), .S(n482) );
  CMPR32X1 U909 ( .A(n467), .B(n466), .C(n465), .CO(n463), .S(n499) );
  XNOR2X1 U910 ( .A(B[16]), .B(A[11]), .Y(n469) );
  NOR2X1 U911 ( .A(n1013), .B(n469), .Y(n527) );
  XNOR2X1 U912 ( .A(n1142), .B(A[12]), .Y(n496) );
  ADDFHX1 U913 ( .A(n474), .B(n473), .CI(n472), .CO(n465), .S(n511) );
  CMPR32X1 U914 ( .A(n480), .B(n479), .C(n478), .CO(n462), .S(n497) );
  NAND2XL U915 ( .A(n482), .B(n481), .Y(mult_x_1_n184) );
  INVXL U916 ( .A(n1269), .Y(n484) );
  XNOR2X1 U917 ( .A(n1001), .B(A[14]), .Y(n525) );
  OAI22X1 U918 ( .A0(n1140), .A1(n525), .B0(n6), .B1(n487), .Y(n506) );
  XNOR2X1 U919 ( .A(n979), .B(A[22]), .Y(n523) );
  OAI22X1 U920 ( .A0(n1024), .A1(n523), .B0(n1022), .B1(n488), .Y(n505) );
  OAI22XL U921 ( .A0(n493), .A1(n529), .B0(n1072), .B1(n492), .Y(n509) );
  XNOR2XL U922 ( .A(n500), .B(A[16]), .Y(n501) );
  OAI22XL U923 ( .A0(n1016), .A1(n501), .B0(n877), .B1(n494), .Y(n508) );
  XNOR2XL U924 ( .A(n964), .B(A[19]), .Y(n549) );
  OAI22XL U925 ( .A0(n11), .A1(n549), .B0(n96), .B1(n495), .Y(n534) );
  XNOR2X1 U926 ( .A(n1142), .B(A[11]), .Y(n550) );
  OAI22XL U927 ( .A0(n10), .A1(n550), .B0(n1143), .B1(n496), .Y(n533) );
  XNOR2X1 U928 ( .A(B[3]), .B(A[23]), .Y(n536) );
  CMPR32X1 U929 ( .A(n509), .B(n508), .C(n507), .CO(n513), .S(n873) );
  CMPR32X1 U930 ( .A(n515), .B(n514), .C(n513), .CO(n563), .S(n558) );
  ADDFHX1 U931 ( .A(n518), .B(n517), .CI(n516), .CO(n481), .S(n519) );
  NOR2XL U932 ( .A(n520), .B(n519), .Y(mult_x_1_n194) );
  NAND2XL U933 ( .A(n520), .B(n519), .Y(mult_x_1_n195) );
  INVXL U934 ( .A(n1271), .Y(n521) );
  XNOR2X1 U935 ( .A(B[16]), .B(A[10]), .Y(n524) );
  XNOR2X1 U936 ( .A(n1001), .B(A[13]), .Y(n551) );
  OAI22XL U937 ( .A0(n1140), .A1(n551), .B0(n6), .B1(n525), .Y(n552) );
  OAI22X1 U938 ( .A0(n1011), .A1(n544), .B0(n531), .B1(n940), .Y(n543) );
  XNOR2X1 U939 ( .A(B[16]), .B(A[9]), .Y(n532) );
  XNOR2X1 U940 ( .A(n534), .B(n533), .Y(n555) );
  XNOR2X1 U941 ( .A(B[3]), .B(A[22]), .Y(n878) );
  XNOR2X1 U942 ( .A(B[16]), .B(A[8]), .Y(n545) );
  NOR2XL U943 ( .A(n1013), .B(n545), .Y(n906) );
  CMPR32X1 U944 ( .A(n548), .B(n547), .C(n546), .CO(n872), .S(n893) );
  OAI22XL U945 ( .A0(n11), .A1(n898), .B0(n96), .B1(n549), .Y(n903) );
  XNOR2X1 U946 ( .A(n1142), .B(A[10]), .Y(n899) );
  OAI22X1 U947 ( .A0(n10), .A1(n899), .B0(n1143), .B1(n550), .Y(n902) );
  XNOR2X1 U948 ( .A(n1001), .B(A[12]), .Y(n900) );
  OAI22XL U949 ( .A0(n1061), .A1(n900), .B0(n6), .B1(n551), .Y(n901) );
  CMPR32X1 U950 ( .A(n557), .B(n556), .C(n555), .CO(n546), .S(n889) );
  CMPR32X1 U951 ( .A(n560), .B(n559), .C(n558), .CO(n561), .S(n870) );
  NOR2X1 U952 ( .A(n565), .B(n564), .Y(mult_x_1_n197) );
  NAND2X1 U953 ( .A(n565), .B(n564), .Y(mult_x_1_n198) );
  INVXL U954 ( .A(n570), .Y(n580) );
  INVXL U955 ( .A(n575), .Y(n577) );
  NAND2X1 U956 ( .A(n594), .B(n593), .Y(n595) );
  NAND2XL U957 ( .A(n600), .B(n599), .Y(n601) );
  XNOR2X1 U958 ( .A(n602), .B(n601), .Y(PRODUCT[25]) );
  INVXL U959 ( .A(n603), .Y(n604) );
  NAND2XL U960 ( .A(n603), .B(n615), .Y(n608) );
  INVXL U961 ( .A(n614), .Y(n606) );
  AOI21XL U962 ( .A0(n612), .A1(n615), .B0(n606), .Y(n607) );
  INVXL U963 ( .A(n612), .Y(n613) );
  OAI21X1 U964 ( .A0(n1089), .A1(n604), .B0(n613), .Y(n617) );
  NAND2XL U965 ( .A(n615), .B(n614), .Y(n616) );
  INVXL U966 ( .A(n1273), .Y(n619) );
  OAI21XL U967 ( .A0(n630), .A1(n1275), .B0(n1276), .Y(n627) );
  INVXL U968 ( .A(n623), .Y(n625) );
  NAND2X1 U969 ( .A(n625), .B(n624), .Y(n626) );
  XNOR2X2 U970 ( .A(n627), .B(n626), .Y(PRODUCT[20]) );
  INVXL U971 ( .A(n1275), .Y(n628) );
  XOR2X1 U972 ( .A(n630), .B(n629), .Y(PRODUCT[19]) );
  XNOR2X1 U973 ( .A(B[16]), .B(A[1]), .Y(n631) );
  NOR2XL U974 ( .A(n1013), .B(n631), .Y(n643) );
  XNOR2X1 U975 ( .A(n1001), .B(A[4]), .Y(n636) );
  XNOR2X1 U976 ( .A(n1001), .B(A[5]), .Y(n653) );
  OAI22XL U977 ( .A0(n1140), .A1(n636), .B0(n6), .B1(n653), .Y(n642) );
  XNOR2X1 U978 ( .A(n976), .B(A[8]), .Y(n673) );
  OAI22X1 U979 ( .A0(n1016), .A1(n637), .B0(n193), .B1(n673), .Y(n672) );
  OAI22X1 U980 ( .A0(n10), .A1(n633), .B0(n1143), .B1(n665), .Y(n671) );
  XNOR2X1 U981 ( .A(B[3]), .B(A[15]), .Y(n638) );
  OAI22X1 U982 ( .A0(n1011), .A1(n683), .B0(n634), .B1(n1084), .Y(n687) );
  XNOR2X1 U983 ( .A(n1142), .B(A[1]), .Y(n690) );
  XNOR2X1 U984 ( .A(B[3]), .B(A[14]), .Y(n639) );
  OAI22X1 U985 ( .A0(n1020), .A1(n696), .B0(n1018), .B1(n639), .Y(n700) );
  XNOR2X1 U986 ( .A(n1001), .B(A[3]), .Y(n692) );
  OAI22X1 U987 ( .A0(n1140), .A1(n692), .B0(n6), .B1(n636), .Y(n699) );
  OAI22X1 U988 ( .A0(n1020), .A1(n639), .B0(n1018), .B1(n638), .Y(n649) );
  XNOR2X1 U989 ( .A(n979), .B(A[11]), .Y(n720) );
  XNOR2X1 U990 ( .A(n976), .B(A[5]), .Y(n697) );
  XNOR2X1 U991 ( .A(n964), .B(A[9]), .Y(n698) );
  CMPR32X1 U992 ( .A(n647), .B(n646), .C(n645), .CO(n681), .S(n717) );
  XNOR2X1 U993 ( .A(n1001), .B(A[6]), .Y(n666) );
  XNOR2XL U994 ( .A(n964), .B(A[12]), .Y(n664) );
  OAI22XL U995 ( .A0(n11), .A1(n654), .B0(n96), .B1(n664), .Y(n669) );
  OAI22X1 U996 ( .A0(n1011), .A1(n655), .B0(n676), .B1(n1084), .Y(n679) );
  XNOR2XL U997 ( .A(B[16]), .B(A[2]), .Y(n656) );
  ADDHXL U998 ( .A(n658), .B(n657), .CO(n667), .S(n645) );
  CMPR32X1 U999 ( .A(n661), .B(n660), .C(n659), .CO(n1048), .S(n705) );
  XNOR2X1 U1000 ( .A(B[7]), .B(A[13]), .Y(n1056) );
  OAI22X1 U1001 ( .A0(n11), .A1(n664), .B0(n96), .B1(n1056), .Y(n1054) );
  OAI22X1 U1002 ( .A0(n10), .A1(n665), .B0(n1143), .B1(n1058), .Y(n1053) );
  XNOR2X1 U1003 ( .A(n1001), .B(A[7]), .Y(n1060) );
  OAI22X1 U1004 ( .A0(n1140), .A1(n666), .B0(n6), .B1(n1060), .Y(n1052) );
  CMPR32X1 U1005 ( .A(n669), .B(n668), .C(n667), .CO(n1043), .S(n659) );
  XNOR2XL U1006 ( .A(n979), .B(A[15]), .Y(n1023) );
  XNOR2XL U1007 ( .A(n904), .B(A[11]), .Y(n1073) );
  XNOR2X1 U1008 ( .A(B[16]), .B(A[3]), .Y(n677) );
  NOR2XL U1009 ( .A(n1013), .B(n677), .Y(n1077) );
  CMPR32X1 U1010 ( .A(n682), .B(n681), .C(n680), .CO(n1083), .S(n716) );
  OAI22X1 U1011 ( .A0(n1011), .A1(n723), .B0(n683), .B1(n940), .Y(n722) );
  OAI22XL U1012 ( .A0(n1074), .A1(n728), .B0(n1072), .B1(n689), .Y(n732) );
  XNOR2X1 U1013 ( .A(n1142), .B(A[0]), .Y(n691) );
  XNOR2X1 U1014 ( .A(n1001), .B(A[2]), .Y(n724) );
  XNOR2X1 U1015 ( .A(n976), .B(A[4]), .Y(n729) );
  XNOR2XL U1016 ( .A(n964), .B(A[8]), .Y(n735) );
  CMPR32X1 U1017 ( .A(n704), .B(n703), .C(n702), .CO(n719), .S(n750) );
  NOR2XL U1018 ( .A(n709), .B(n708), .Y(mult_x_1_n276) );
  NAND2XL U1019 ( .A(n709), .B(n708), .Y(mult_x_1_n277) );
  INVXL U1020 ( .A(n1277), .Y(n711) );
  XOR2X1 U1021 ( .A(n713), .B(n712), .Y(PRODUCT[18]) );
  XNOR2X1 U1022 ( .A(n979), .B(A[10]), .Y(n733) );
  CMPR22X1 U1023 ( .A(n722), .B(n721), .CO(n727), .S(n757) );
  XNOR2X1 U1024 ( .A(n5), .B(A[13]), .Y(n736) );
  OAI22XL U1025 ( .A0(n1140), .A1(n787), .B0(n6), .B1(n724), .Y(n759) );
  OAI22XL U1026 ( .A0(n1074), .A1(n762), .B0(n1072), .B1(n728), .Y(n770) );
  XNOR2X1 U1027 ( .A(n976), .B(A[3]), .Y(n789) );
  OAI22X1 U1028 ( .A0(n1011), .A1(n737), .B0(n736), .B1(n1084), .Y(n795) );
  OAI22X1 U1029 ( .A0(n1140), .A1(n739), .B0(n6), .B1(n738), .Y(n794) );
  NOR2XL U1030 ( .A(n744), .B(n743), .Y(mult_x_1_n281) );
  NAND2XL U1031 ( .A(n745), .B(n1280), .Y(n746) );
  CMPR32X1 U1032 ( .A(n752), .B(n751), .C(n750), .CO(n740), .S(n781) );
  CMPR32X1 U1033 ( .A(n755), .B(n754), .C(n753), .CO(n752), .S(n804) );
  CMPR32X1 U1034 ( .A(n758), .B(n757), .C(n756), .CO(n773), .S(n803) );
  NOR2XL U1035 ( .A(n775), .B(n774), .Y(mult_x_1_n286) );
  NAND2XL U1036 ( .A(n775), .B(n774), .Y(mult_x_1_n287) );
  INVXL U1037 ( .A(n1281), .Y(n776) );
  NAND2XL U1038 ( .A(n776), .B(n1282), .Y(n777) );
  XNOR2X1 U1039 ( .A(n1001), .B(A[0]), .Y(n788) );
  OAI22X1 U1040 ( .A0(n1140), .A1(n788), .B0(n6), .B1(n787), .Y(n812) );
  CMPR32X1 U1041 ( .A(n801), .B(n800), .C(n799), .CO(n823), .S(n826) );
  OAI21XL U1042 ( .A0(n844), .A1(n1248), .B0(n1249), .Y(n807) );
  CMPR32X1 U1043 ( .A(n816), .B(n815), .C(n814), .CO(n809), .S(n830) );
  CMPR32X1 U1044 ( .A(n819), .B(n818), .C(n817), .CO(n829), .S(n851) );
  CMPR32X1 U1045 ( .A(n822), .B(n821), .C(n820), .CO(n833), .S(n835) );
  NOR2X1 U1046 ( .A(n839), .B(n838), .Y(mult_x_1_n306) );
  INVX1 U1047 ( .A(mult_x_1_n306), .Y(n845) );
  NAND2X1 U1048 ( .A(n841), .B(n840), .Y(n1085) );
  INVX1 U1049 ( .A(n1085), .Y(n842) );
  NAND2XL U1050 ( .A(n845), .B(mult_x_1_n307), .Y(mult_x_1_n84) );
  CMPR32X1 U1051 ( .A(n848), .B(n847), .C(n846), .CO(n838), .S(n853) );
  CMPR32X1 U1052 ( .A(n851), .B(n850), .C(n849), .CO(n852), .S(n249) );
  NAND2XL U1053 ( .A(n1093), .B(n1091), .Y(mult_x_1_n85) );
  AOI21XL U1054 ( .A0(n855), .A1(n1090), .B0(n1092), .Y(mult_x_1_n316) );
  INVXL U1055 ( .A(n857), .Y(n859) );
  NAND2XL U1056 ( .A(n859), .B(n858), .Y(n860) );
  NAND2XL U1057 ( .A(n7), .B(n862), .Y(n863) );
  INVXL U1058 ( .A(n865), .Y(n1183) );
  AOI21XL U1059 ( .A0(n1183), .A1(n1180), .B0(n866), .Y(n869) );
  ADDFHX1 U1060 ( .A(n875), .B(n874), .CI(n873), .CO(n560), .S(n897) );
  XNOR2X1 U1061 ( .A(n976), .B(A[13]), .Y(n910) );
  XNOR2X1 U1062 ( .A(B[3]), .B(A[21]), .Y(n911) );
  XNOR2X1 U1063 ( .A(n979), .B(A[19]), .Y(n912) );
  CMPR32X1 U1064 ( .A(n885), .B(n884), .C(n883), .CO(n886), .S(n922) );
  CMPR32X1 U1065 ( .A(n891), .B(n890), .C(n889), .CO(n892), .S(n925) );
  ADDFHX1 U1066 ( .A(n897), .B(n896), .CI(n895), .CO(mult_x_1_n521), .S(
        mult_x_1_n522) );
  XNOR2X1 U1067 ( .A(n1142), .B(A[9]), .Y(n932) );
  OAI22X2 U1068 ( .A0(n10), .A1(n932), .B0(n1143), .B1(n899), .Y(n935) );
  XNOR2XL U1069 ( .A(n1001), .B(A[11]), .Y(n933) );
  OAI22XL U1070 ( .A0(n1061), .A1(n933), .B0(n6), .B1(n900), .Y(n934) );
  ADDFHX1 U1071 ( .A(n903), .B(n902), .CI(n901), .CO(n891), .S(n920) );
  ADDHXL U1072 ( .A(n907), .B(n906), .CO(n883), .S(n917) );
  OAI22X1 U1073 ( .A0(n1011), .A1(n941), .B0(n908), .B1(n1084), .Y(n939) );
  XNOR2X1 U1074 ( .A(n976), .B(A[12]), .Y(n943) );
  XNOR2X1 U1075 ( .A(B[3]), .B(A[20]), .Y(n944) );
  XNOR2X1 U1076 ( .A(n979), .B(A[18]), .Y(n945) );
  CMPR32X1 U1077 ( .A(n918), .B(n916), .C(n917), .CO(n919), .S(n955) );
  CMPR32X1 U1078 ( .A(n921), .B(n920), .C(n919), .CO(n930), .S(n959) );
  ADDFHX1 U1079 ( .A(n927), .B(n926), .CI(n925), .CO(n896), .S(n928) );
  ADDFHX1 U1080 ( .A(n930), .B(n929), .CI(n928), .CO(mult_x_1_n537), .S(
        mult_x_1_n538) );
  XNOR2X1 U1081 ( .A(n1001), .B(A[10]), .Y(n967) );
  OAI22XL U1082 ( .A0(n1140), .A1(n967), .B0(n6), .B1(n933), .Y(n968) );
  OAI22XL U1083 ( .A0(n1074), .A1(n971), .B0(n1072), .B1(n937), .Y(n951) );
  XNOR2X1 U1084 ( .A(B[16]), .B(A[6]), .Y(n942) );
  NOR2XL U1085 ( .A(n1013), .B(n942), .Y(n972) );
  XNOR2X1 U1086 ( .A(n976), .B(A[11]), .Y(n977) );
  XNOR2X1 U1087 ( .A(B[3]), .B(A[19]), .Y(n978) );
  XNOR2XL U1088 ( .A(n979), .B(A[17]), .Y(n980) );
  CMPR32X1 U1089 ( .A(n948), .B(n947), .C(n946), .CO(n957), .S(n991) );
  CMPR32X1 U1090 ( .A(n951), .B(n950), .C(n949), .CO(n952), .S(n990) );
  ADDFHX1 U1091 ( .A(n960), .B(n959), .CI(n958), .CO(n929), .S(n961) );
  ADDFHX1 U1092 ( .A(n963), .B(n962), .CI(n961), .CO(mult_x_1_n553), .S(
        mult_x_1_n554) );
  OAI22X1 U1093 ( .A0(n11), .A1(n999), .B0(n96), .B1(n965), .Y(n1005) );
  XNOR2X1 U1094 ( .A(n1142), .B(A[7]), .Y(n1000) );
  OAI22X2 U1095 ( .A0(n10), .A1(n1000), .B0(n1143), .B1(n966), .Y(n1004) );
  XNOR2X1 U1096 ( .A(n1001), .B(A[9]), .Y(n1002) );
  OAI22X1 U1097 ( .A0(n1140), .A1(n1002), .B0(n6), .B1(n967), .Y(n1003) );
  XNOR2XL U1098 ( .A(n904), .B(A[13]), .Y(n1006) );
  OAI22XL U1099 ( .A0(n1074), .A1(n1006), .B0(n1072), .B1(n971), .Y(n986) );
  ADDHXL U1100 ( .A(n973), .B(n972), .CO(n949), .S(n985) );
  OAI22X1 U1101 ( .A0(n1011), .A1(n1009), .B0(n974), .B1(n1084), .Y(n1008) );
  XNOR2XL U1102 ( .A(B[16]), .B(A[5]), .Y(n975) );
  OAI22X1 U1103 ( .A0(n1016), .A1(n1014), .B0(n877), .B1(n977), .Y(n1027) );
  XNOR2X1 U1104 ( .A(B[3]), .B(A[18]), .Y(n1017) );
  XNOR2XL U1105 ( .A(n979), .B(A[16]), .Y(n1021) );
  OAI22XL U1106 ( .A0(n1024), .A1(n1021), .B0(n1022), .B1(n980), .Y(n1025) );
  CMPR32X1 U1107 ( .A(n983), .B(n982), .C(n981), .CO(n992), .S(n1035) );
  CMPR32X1 U1108 ( .A(n986), .B(n984), .C(n985), .CO(n987), .S(n1034) );
  ADDFHX1 U1109 ( .A(n995), .B(n994), .CI(n993), .CO(n962), .S(n996) );
  ADDFHX1 U1110 ( .A(n998), .B(n997), .CI(n996), .CO(mult_x_1_n569), .S(
        mult_x_1_n570) );
  OAI22X1 U1111 ( .A0(n11), .A1(n1055), .B0(n96), .B1(n999), .Y(n1099) );
  XNOR2X1 U1112 ( .A(n1001), .B(A[8]), .Y(n1059) );
  OAI22X1 U1113 ( .A0(n1061), .A1(n1059), .B0(n6), .B1(n1002), .Y(n1097) );
  XNOR2XL U1114 ( .A(n904), .B(A[12]), .Y(n1071) );
  OAI22XL U1115 ( .A0(n1074), .A1(n1071), .B0(n1072), .B1(n1006), .Y(n1030) );
  OAI22X1 U1116 ( .A0(n1011), .A1(n1010), .B0(n1009), .B1(n1084), .Y(n1076) );
  XNOR2XL U1117 ( .A(B[16]), .B(A[4]), .Y(n1012) );
  NOR2XL U1118 ( .A(n1013), .B(n1012), .Y(n1075) );
  OAI22XL U1119 ( .A0(n1024), .A1(n1023), .B0(n1022), .B1(n1021), .Y(n1068) );
  CMPR32X1 U1120 ( .A(n1030), .B(n1029), .C(n1028), .CO(n1031), .S(n1109) );
  CMPR32X1 U1121 ( .A(n1033), .B(n1032), .C(n1031), .CO(n1042), .S(n1113) );
  ADDFHX1 U1122 ( .A(n1039), .B(n1038), .CI(n1037), .CO(n997), .S(n1040) );
  ADDFHX1 U1123 ( .A(n1042), .B(n1041), .CI(n1040), .CO(mult_x_1_n585), .S(
        mult_x_1_n586) );
  CMPR32X1 U1124 ( .A(n1045), .B(n1044), .C(n1043), .CO(n1081), .S(n1047) );
  OAI22X1 U1125 ( .A0(n11), .A1(n1056), .B0(n96), .B1(n1055), .Y(n1096) );
  OAI22X1 U1126 ( .A0(n10), .A1(n1058), .B0(n1143), .B1(n1057), .Y(n1095) );
  CMPR32X1 U1127 ( .A(n1064), .B(n1062), .C(n1063), .CO(n1115), .S(n1049) );
  CMPR32X1 U1128 ( .A(n1070), .B(n1069), .C(n1068), .CO(n1111), .S(n1104) );
  OAI22XL U1129 ( .A0(n1074), .A1(n1073), .B0(n1072), .B1(n1071), .Y(n1102) );
  ADDHXL U1130 ( .A(n1078), .B(n1077), .CO(n1100), .S(n1063) );
  ADDFHX1 U1131 ( .A(n1081), .B(n1080), .CI(n1079), .CO(mult_x_1_n633), .S(
        mult_x_1_n634) );
  NAND2X1 U1132 ( .A(n93), .B(n618), .Y(n1088) );
  CMPR32X1 U1133 ( .A(n1102), .B(n1101), .C(n1100), .CO(n1106), .S(n1103) );
  ADDFX2 U1134 ( .A(n1108), .B(n1107), .CI(n1106), .CO(n1126), .S(n1122) );
  CMPR32X1 U1135 ( .A(n1111), .B(n1110), .C(n1109), .CO(n1114), .S(n1121) );
  ADDFX2 U1136 ( .A(n1117), .B(n1116), .CI(n1115), .CO(n1129), .S(n1119) );
  ADDFHX1 U1137 ( .A(n1126), .B(n1125), .CI(n1124), .CO(mult_x_1_n601), .S(
        n1131) );
  NAND2XL U1138 ( .A(n1131), .B(n1130), .Y(mult_x_1_n263) );
  CMPR32X1 U1139 ( .A(n1136), .B(n1135), .C(n1134), .CO(n1152), .S(n1149) );
  XNOR2X1 U1140 ( .A(B[16]), .B(A[22]), .Y(n1137) );
  XNOR2X1 U1141 ( .A(B[16]), .B(A[23]), .Y(n1141) );
  XNOR2X1 U1142 ( .A(n1142), .B(A[25]), .Y(n1163) );
  CMPR32X1 U1143 ( .A(n1147), .B(n1146), .C(n1145), .CO(n1158), .S(n1151) );
  CMPR32X1 U1144 ( .A(n1150), .B(n1149), .C(n1148), .CO(n1157), .S(n276) );
  CMPR32X1 U1145 ( .A(n1153), .B(n1152), .C(n1151), .CO(n1155), .S(n1156) );
  CMPR32X1 U1146 ( .A(n1160), .B(n1159), .C(n1158), .CO(n1170), .S(n1154) );
  OAI2BB1X1 U1147 ( .A0N(n1165), .A1N(n10), .B0(n1164), .Y(n1166) );
  XOR3X2 U1148 ( .A(n1168), .B(n1167), .C(n1166), .Y(n1169) );
  OAI21XL U1149 ( .A0(n1246), .A1(n1176), .B0(n1175), .Y(n1179) );
  OAI21XL U1150 ( .A0(n1193), .A1(n1190), .B0(n1191), .Y(n1189) );
  INVXL U1151 ( .A(n1185), .Y(n1187) );
  OAI21XL U1152 ( .A0(n1255), .A1(n1258), .B0(n1256), .Y(n1203) );
  OAI21XL U1153 ( .A0(n1246), .A1(n1196), .B0(n1195), .Y(n1198) );
  OAI21XL U1154 ( .A0(n1246), .A1(n1208), .B0(n1207), .Y(n1211) );
  XNOR2XL U1155 ( .A(n1227), .B(n1226), .Y(n1327) );
  XOR2XL U1156 ( .A(n1232), .B(n1231), .Y(n1326) );
  OAI21XL U1157 ( .A0(n1236), .A1(n1251), .B0(n1252), .Y(n1237) );
  AOI21XL U1158 ( .A0(n1239), .A1(n1238), .B0(n1237), .Y(n1240) );
  OAI21XL U1159 ( .A0(n1242), .A1(n1241), .B0(n1240), .Y(n1243) );
  OAI21XL U1160 ( .A0(n1246), .A1(n1245), .B0(n1244), .Y(n1247) );
  XNOR2XL U1161 ( .A(n1247), .B(n1250), .Y(PRODUCT[40]) );
endmodule


module FFT2048_DW02_mult_2_stage_J1_1 ( A, B, TC, CLK, PRODUCT );
  input [25:0] A;
  input [16:0] B;
  output [42:0] PRODUCT;
  input TC, CLK;
  wire   n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, mult_x_1_n649, mult_x_1_n634, mult_x_1_n633,
         mult_x_1_n618, mult_x_1_n617, mult_x_1_n602, mult_x_1_n601,
         mult_x_1_n586, mult_x_1_n585, mult_x_1_n570, mult_x_1_n569,
         mult_x_1_n554, mult_x_1_n553, mult_x_1_n538, mult_x_1_n537,
         mult_x_1_n522, mult_x_1_n521, mult_x_1_n508, mult_x_1_n507,
         mult_x_1_n494, mult_x_1_n321, mult_x_1_n316, mult_x_1_n309,
         mult_x_1_n307, mult_x_1_n306, mult_x_1_n296, mult_x_1_n295,
         mult_x_1_n293, mult_x_1_n292, mult_x_1_n287, mult_x_1_n286,
         mult_x_1_n282, mult_x_1_n281, mult_x_1_n277, mult_x_1_n276,
         mult_x_1_n195, mult_x_1_n194, mult_x_1_n184, mult_x_1_n183,
         mult_x_1_n177, mult_x_1_n176, mult_x_1_n170, mult_x_1_n169,
         mult_x_1_n161, mult_x_1_n160, mult_x_1_n152, mult_x_1_n151,
         mult_x_1_n137, mult_x_1_n136, mult_x_1_n130, mult_x_1_n129,
         mult_x_1_n121, mult_x_1_n120, mult_x_1_n110, mult_x_1_n109,
         mult_x_1_n86, mult_x_1_n85, mult_x_1_n84, mult_x_1_n83, mult_x_1_n58,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380;

  DFFHQX4 mult_x_1_clk_r_REG46_S1 ( .D(mult_x_1_n286), .CK(CLK), .Q(n1349) );
  DFFHQXL mult_x_1_clk_r_REG16_S1 ( .D(mult_x_1_n169), .CK(CLK), .Q(n1337) );
  DFFHQXL mult_x_1_clk_r_REG18_S1 ( .D(mult_x_1_n160), .CK(CLK), .Q(n1335) );
  DFFHQXL mult_x_1_clk_r_REG20_S1 ( .D(mult_x_1_n151), .CK(CLK), .Q(n1333) );
  DFFHQX4 mult_x_1_clk_r_REG40_S1 ( .D(mult_x_1_n649), .CK(CLK), .Q(n1380) );
  DFFHQX4 mult_x_1_clk_r_REG39_S1 ( .D(mult_x_1_n634), .CK(CLK), .Q(n1379) );
  DFFHQX4 mult_x_1_clk_r_REG38_S1 ( .D(mult_x_1_n633), .CK(CLK), .Q(n1378) );
  DFFHQX4 mult_x_1_clk_r_REG37_S1 ( .D(mult_x_1_n618), .CK(CLK), .Q(n1377) );
  DFFHQX4 mult_x_1_clk_r_REG34_S1 ( .D(mult_x_1_n601), .CK(CLK), .Q(n1374) );
  DFFHQX4 mult_x_1_clk_r_REG33_S1 ( .D(mult_x_1_n586), .CK(CLK), .Q(n1373) );
  DFFHQX4 mult_x_1_clk_r_REG32_S1 ( .D(mult_x_1_n585), .CK(CLK), .Q(n1372) );
  DFFHQX4 mult_x_1_clk_r_REG31_S1 ( .D(mult_x_1_n570), .CK(CLK), .Q(n1371) );
  DFFHQX4 mult_x_1_clk_r_REG7_S1 ( .D(mult_x_1_n508), .CK(CLK), .Q(n1363) );
  DFFHQX4 mult_x_1_clk_r_REG56_S1 ( .D(mult_x_1_n309), .CK(CLK), .Q(n1359) );
  DFFHQX4 mult_x_1_clk_r_REG50_S1 ( .D(mult_x_1_n296), .CK(CLK), .Q(n1358) );
  DFFHQX4 mult_x_1_clk_r_REG51_S1 ( .D(mult_x_1_n295), .CK(CLK), .Q(n1353) );
  DFFHQX4 mult_x_1_clk_r_REG48_S1 ( .D(mult_x_1_n292), .CK(CLK), .Q(n1351) );
  DFFHQX4 mult_x_1_clk_r_REG44_S1 ( .D(mult_x_1_n281), .CK(CLK), .Q(n1347) );
  DFFHQXL clk_r_REG61_S1 ( .D(n1394), .CK(CLK), .Q(PRODUCT[10]) );
  DFFHQXL mult_x_1_clk_r_REG13_S1 ( .D(mult_x_1_n177), .CK(CLK), .Q(n1340) );
  DFFHQXL mult_x_1_clk_r_REG14_S1 ( .D(mult_x_1_n176), .CK(CLK), .Q(n1339) );
  DFFHQXL mult_x_1_clk_r_REG19_S1 ( .D(mult_x_1_n152), .CK(CLK), .Q(n1334) );
  DFFHQXL mult_x_1_clk_r_REG15_S1 ( .D(mult_x_1_n170), .CK(CLK), .Q(n1338) );
  DFFHQXL clk_r_REG62_S1 ( .D(n1395), .CK(CLK), .Q(PRODUCT[9]) );
  DFFHQXL mult_x_1_clk_r_REG11_S1 ( .D(mult_x_1_n184), .CK(CLK), .Q(n1342) );
  DFFHQXL mult_x_1_clk_r_REG17_S1 ( .D(mult_x_1_n161), .CK(CLK), .Q(n1336) );
  DFFHQXL mult_x_1_clk_r_REG60_S1 ( .D(mult_x_1_n321), .CK(CLK), .Q(n1323) );
  DFFHQXL mult_x_1_clk_r_REG12_S1 ( .D(mult_x_1_n183), .CK(CLK), .Q(n1341) );
  DFFHQXL clk_r_REG59_S1 ( .D(n1393), .CK(CLK), .Q(PRODUCT[11]) );
  DFFHQXL mult_x_1_clk_r_REG9_S1 ( .D(mult_x_1_n195), .CK(CLK), .Q(n1344) );
  DFFHQXL clk_r_REG63_S1 ( .D(n1396), .CK(CLK), .Q(PRODUCT[8]) );
  DFFHQXL clk_r_REG64_S1 ( .D(n1397), .CK(CLK), .Q(PRODUCT[7]) );
  DFFHQXL clk_r_REG65_S1 ( .D(n1398), .CK(CLK), .Q(PRODUCT[6]) );
  DFFHQXL clk_r_REG66_S1 ( .D(n1399), .CK(CLK), .Q(PRODUCT[5]) );
  DFFHQXL clk_r_REG67_S1 ( .D(n1400), .CK(CLK), .Q(PRODUCT[4]) );
  DFFHQXL clk_r_REG68_S1 ( .D(n1401), .CK(CLK), .Q(PRODUCT[3]) );
  DFFHQXL clk_r_REG69_S1 ( .D(n1402), .CK(CLK), .Q(PRODUCT[2]) );
  DFFHQXL clk_r_REG70_S1 ( .D(n1403), .CK(CLK), .Q(PRODUCT[1]) );
  DFFHQXL clk_r_REG71_S1 ( .D(n1404), .CK(CLK), .Q(PRODUCT[0]) );
  DFFHQXL mult_x_1_clk_r_REG57_S1 ( .D(mult_x_1_n86), .CK(CLK), .Q(n1357) );
  DFFHQX1 mult_x_1_clk_r_REG55_S1 ( .D(mult_x_1_n85), .CK(CLK), .Q(n1356) );
  DFFHQXL mult_x_1_clk_r_REG52_S1 ( .D(mult_x_1_n84), .CK(CLK), .Q(n1355) );
  DFFHQXL mult_x_1_clk_r_REG49_S1 ( .D(mult_x_1_n83), .CK(CLK), .Q(n1354) );
  DFFHQX1 mult_x_1_clk_r_REG47_S1 ( .D(mult_x_1_n293), .CK(CLK), .Q(n1352) );
  DFFHQXL mult_x_1_clk_r_REG10_S1 ( .D(mult_x_1_n194), .CK(CLK), .Q(n1343) );
  DFFHQXL mult_x_1_clk_r_REG21_S1 ( .D(mult_x_1_n137), .CK(CLK), .Q(n1332) );
  DFFHQXL mult_x_1_clk_r_REG23_S1 ( .D(mult_x_1_n130), .CK(CLK), .Q(n1330) );
  DFFHQXL mult_x_1_clk_r_REG24_S1 ( .D(mult_x_1_n129), .CK(CLK), .Q(n1329) );
  DFFHQXL mult_x_1_clk_r_REG25_S1 ( .D(mult_x_1_n121), .CK(CLK), .Q(n1328) );
  DFFHQXL mult_x_1_clk_r_REG26_S1 ( .D(mult_x_1_n120), .CK(CLK), .Q(n1327) );
  DFFHQXL mult_x_1_clk_r_REG27_S1 ( .D(mult_x_1_n110), .CK(CLK), .Q(n1326) );
  DFFHQXL mult_x_1_clk_r_REG28_S1 ( .D(mult_x_1_n109), .CK(CLK), .Q(n1325) );
  DFFHQXL mult_x_1_clk_r_REG29_S1 ( .D(mult_x_1_n58), .CK(CLK), .Q(n1324) );
  DFFHQXL mult_x_1_clk_r_REG53_S1 ( .D(mult_x_1_n307), .CK(CLK), .Q(n1322) );
  DFFHQXL mult_x_1_clk_r_REG54_S1 ( .D(mult_x_1_n306), .CK(CLK), .Q(n1321) );
  DFFHQXL mult_x_1_clk_r_REG58_S1 ( .D(mult_x_1_n316), .CK(CLK), .Q(n1360) );
  DFFHQXL mult_x_1_clk_r_REG22_S1 ( .D(mult_x_1_n136), .CK(CLK), .Q(n1331) );
  DFFHQX2 mult_x_1_clk_r_REG42_S1 ( .D(mult_x_1_n276), .CK(CLK), .Q(n1345) );
  DFFHQX4 mult_x_1_clk_r_REG45_S1 ( .D(mult_x_1_n287), .CK(CLK), .Q(n1350) );
  DFFHQX1 mult_x_1_clk_r_REG3_S1 ( .D(mult_x_1_n538), .CK(CLK), .Q(n1367) );
  DFFHQXL mult_x_1_clk_r_REG8_S1 ( .D(mult_x_1_n494), .CK(CLK), .Q(n1361) );
  DFFHQX1 mult_x_1_clk_r_REG43_S1 ( .D(mult_x_1_n282), .CK(CLK), .Q(n1348) );
  DFFHQX1 mult_x_1_clk_r_REG41_S1 ( .D(mult_x_1_n277), .CK(CLK), .Q(n1346) );
  DFFHQX1 mult_x_1_clk_r_REG4_S1 ( .D(mult_x_1_n521), .CK(CLK), .Q(n1364) );
  DFFHQX1 mult_x_1_clk_r_REG30_S1 ( .D(mult_x_1_n569), .CK(CLK), .Q(n1370) );
  DFFHQX1 mult_x_1_clk_r_REG1_S1 ( .D(mult_x_1_n554), .CK(CLK), .Q(n1369) );
  DFFHQX1 mult_x_1_clk_r_REG0_S1 ( .D(mult_x_1_n553), .CK(CLK), .Q(n1368) );
  DFFHQX2 mult_x_1_clk_r_REG36_S1 ( .D(mult_x_1_n617), .CK(CLK), .Q(n1376) );
  DFFHQX2 mult_x_1_clk_r_REG2_S1 ( .D(mult_x_1_n537), .CK(CLK), .Q(n1366) );
  DFFHQX2 mult_x_1_clk_r_REG5_S1 ( .D(mult_x_1_n522), .CK(CLK), .Q(n1365) );
  DFFHQX2 mult_x_1_clk_r_REG35_S1 ( .D(mult_x_1_n602), .CK(CLK), .Q(n1375) );
  DFFHQX1 mult_x_1_clk_r_REG6_S1 ( .D(mult_x_1_n507), .CK(CLK), .Q(n1362) );
  CMPR32X1 U1 ( .A(n361), .B(n360), .C(n359), .CO(n337), .S(n362) );
  OAI2BB1X1 U2 ( .A0N(n1005), .A1N(n1006), .B0(n91), .Y(n966) );
  OAI2BB1X1 U3 ( .A0N(n79), .A1N(n1144), .B0(n78), .Y(n1121) );
  ADDFHX1 U4 ( .A(n805), .B(n804), .CI(n803), .CO(n502), .S(mult_x_1_n494) );
  ADDFHX1 U5 ( .A(n667), .B(n666), .CI(n665), .CO(n660), .S(n691) );
  ADDFHX1 U6 ( .A(n1152), .B(n1151), .CI(n1150), .CO(n1153), .S(n661) );
  NAND2X1 U7 ( .A(n88), .B(n87), .Y(n1148) );
  ADDFHX1 U8 ( .A(n1095), .B(n1094), .CI(n1093), .CO(n1057), .S(n1096) );
  ADDFHX1 U9 ( .A(n689), .B(n688), .CI(n687), .CO(n666), .S(n695) );
  ADDFHX1 U10 ( .A(n1119), .B(n1118), .CI(n1117), .CO(n1097), .S(n1120) );
  OAI21XL U11 ( .A0(n1142), .A1(n1143), .B0(n18), .Y(n88) );
  ADDFX2 U12 ( .A(n494), .B(n493), .CI(n492), .CO(n483), .S(n843) );
  ADDFHX1 U13 ( .A(n1049), .B(n1048), .CI(n1047), .CO(n1058), .S(n1094) );
  ADDFHX1 U14 ( .A(n762), .B(n761), .CI(n760), .CO(n765), .S(n764) );
  ADDFHX1 U15 ( .A(n759), .B(n758), .CI(n757), .CO(n723), .S(n766) );
  ADDFX2 U16 ( .A(n635), .B(n634), .CI(n633), .CO(n1142), .S(n667) );
  ADDFX2 U17 ( .A(n1130), .B(n1129), .CI(n1128), .CO(n1131), .S(n787) );
  ADDFX2 U18 ( .A(n464), .B(n463), .CI(n462), .CO(n467), .S(n492) );
  ADDFX2 U19 ( .A(n1080), .B(n1079), .CI(n1078), .CO(n1116), .S(n1139) );
  ADDFX2 U20 ( .A(n743), .B(n742), .CI(n741), .CO(n758), .S(n760) );
  CMPR32X1 U21 ( .A(n907), .B(n906), .C(n905), .CO(n892), .S(n922) );
  NAND2BXL U22 ( .AN(n1110), .B(n62), .Y(n61) );
  OAI21X1 U23 ( .A0(n89), .A1(n75), .B0(n73), .Y(n1043) );
  ADDFHX1 U24 ( .A(n728), .B(n727), .CI(n726), .CO(n720), .S(n762) );
  ADDFHX1 U25 ( .A(n1104), .B(n1103), .CI(n1102), .CO(n1089), .S(n1112) );
  ADDFHX1 U26 ( .A(n783), .B(n782), .CI(n781), .CO(n1126), .S(n1128) );
  NOR2X1 U27 ( .A(n202), .B(n201), .Y(n1258) );
  XOR2X1 U28 ( .A(n986), .B(n76), .Y(n75) );
  XOR2XL U29 ( .A(n986), .B(n28), .Y(n27) );
  NAND2BXL U30 ( .AN(n987), .B(n74), .Y(n73) );
  OAI21XL U31 ( .A0(n749), .A1(n750), .B0(n31), .Y(n29) );
  OAI22X1 U32 ( .A0(n1033), .A1(n605), .B0(n1031), .B1(n597), .Y(n623) );
  OAI22X1 U33 ( .A0(n6), .A1(n485), .B0(n1035), .B1(n414), .Y(n476) );
  ADDFHX1 U34 ( .A(n231), .B(n230), .CI(n229), .CO(n237), .S(n236) );
  ADDFHX1 U35 ( .A(n1101), .B(n1100), .CI(n1099), .CO(n1113), .S(n1109) );
  CLKBUFX3 U36 ( .A(n380), .Y(n1030) );
  INVXL U37 ( .A(n1162), .Y(n5) );
  NOR2XL U38 ( .A(n1062), .B(n1065), .Y(n54) );
  BUFX3 U39 ( .A(n457), .Y(n1063) );
  BUFX3 U40 ( .A(n580), .Y(n1206) );
  CLKBUFX8 U41 ( .A(B[16]), .Y(n1224) );
  OAI21X2 U42 ( .A0(n1031), .A1(n714), .B0(n102), .Y(n90) );
  CLKBUFX3 U43 ( .A(n652), .Y(n1040) );
  NAND2X1 U44 ( .A(n149), .B(n155), .Y(n652) );
  BUFX4 U45 ( .A(n628), .Y(n1061) );
  OAI21X1 U46 ( .A0(n1072), .A1(n251), .B0(n43), .Y(n42) );
  NAND2X4 U47 ( .A(n205), .B(n206), .Y(n214) );
  XNOR2X1 U48 ( .A(n529), .B(n528), .Y(PRODUCT[27]) );
  XOR2X1 U49 ( .A(n568), .B(n567), .Y(PRODUCT[21]) );
  NOR2X2 U50 ( .A(n1379), .B(n1380), .Y(n571) );
  XNOR2X2 U51 ( .A(B[2]), .B(B[1]), .Y(n819) );
  OAI22X1 U52 ( .A0(n6), .A1(n851), .B0(n819), .B1(n818), .Y(n854) );
  OAI22X1 U53 ( .A0(n6), .A1(n989), .B0(n1035), .B1(n948), .Y(n994) );
  OAI22X1 U54 ( .A0(n6), .A1(n914), .B0(n1035), .B1(n882), .Y(n917) );
  BUFX3 U55 ( .A(n177), .Y(n6) );
  OAI22X1 U56 ( .A0(n170), .A1(n261), .B0(n712), .B1(n1123), .Y(n737) );
  OAI22X1 U57 ( .A0(n1040), .A1(n915), .B0(n1038), .B1(n883), .Y(n916) );
  ADDFX2 U58 ( .A(n247), .B(n246), .CI(n245), .CO(n276), .S(n254) );
  OAI22X1 U59 ( .A0(n6), .A1(n213), .B0(n1035), .B1(n244), .Y(n247) );
  AOI21XL U60 ( .A0(n294), .A1(n436), .B0(n122), .Y(n1310) );
  AOI21XL U61 ( .A0(n338), .A1(n124), .B0(n339), .Y(n127) );
  OAI21XL U62 ( .A0(n1310), .A1(n1245), .B0(n1244), .Y(n1279) );
  XNOR2XL U63 ( .A(n991), .B(n1012), .Y(n243) );
  XNOR2XL U64 ( .A(B[1]), .B(n977), .Y(n711) );
  XNOR2XL U65 ( .A(n991), .B(n1124), .Y(n166) );
  XNOR2XL U66 ( .A(n1187), .B(n949), .Y(n420) );
  XNOR2XL U67 ( .A(B[1]), .B(n1212), .Y(n879) );
  XNOR2XL U68 ( .A(n681), .B(n1158), .Y(n914) );
  XNOR2XL U69 ( .A(n681), .B(n947), .Y(n989) );
  XNOR2XL U70 ( .A(n1021), .B(A[25]), .Y(n309) );
  XNOR2XL U71 ( .A(B[9]), .B(n1201), .Y(n376) );
  XNOR2XL U72 ( .A(n681), .B(n968), .Y(n599) );
  XOR2XL U73 ( .A(n302), .B(n985), .Y(n608) );
  XNOR2XL U74 ( .A(B[9]), .B(n947), .Y(n812) );
  XNOR2XL U75 ( .A(n1214), .B(n945), .Y(n871) );
  BUFX3 U76 ( .A(n819), .Y(n1035) );
  XNOR2XL U77 ( .A(B[1]), .B(n640), .Y(n169) );
  OAI2BB1X1 U78 ( .A0N(n61), .A1N(n1108), .B0(n60), .Y(n1146) );
  ADDFX2 U79 ( .A(n477), .B(n476), .CI(n475), .CO(n452), .S(n496) );
  XOR2XL U80 ( .A(n1267), .B(n1266), .Y(n1398) );
  XOR2XL U81 ( .A(n792), .B(n791), .Y(n1394) );
  INVX4 U82 ( .A(B[7]), .Y(n302) );
  NAND2X1 U83 ( .A(n279), .B(n278), .Y(n771) );
  NAND2X1 U84 ( .A(n37), .B(n59), .Y(n36) );
  NAND2XL U85 ( .A(n661), .B(n660), .Y(mult_x_1_n282) );
  NAND2BX1 U86 ( .AN(n77), .B(n80), .Y(n79) );
  NAND2X1 U87 ( .A(n238), .B(n237), .Y(n795) );
  INVX1 U88 ( .A(n1131), .Y(n84) );
  INVX1 U89 ( .A(n787), .Y(n83) );
  NAND2XL U90 ( .A(n39), .B(n252), .Y(n38) );
  OAI2BB1X1 U91 ( .A0N(n353), .A1N(n116), .B0(n115), .Y(n395) );
  OAI2BB1X1 U92 ( .A0N(n1069), .A1N(n138), .B0(n137), .Y(n1049) );
  NAND2XL U93 ( .A(n23), .B(n22), .Y(n21) );
  NAND2XL U94 ( .A(n64), .B(n994), .Y(n63) );
  OAI2BB1XL U95 ( .A0N(n951), .A1N(n93), .B0(n92), .Y(n961) );
  NAND2X1 U96 ( .A(n1110), .B(n1109), .Y(n60) );
  XOR3X2 U97 ( .A(n1109), .B(n1110), .C(n1108), .Y(n18) );
  NAND2XL U98 ( .A(n106), .B(n778), .Y(n105) );
  NAND2BXL U99 ( .AN(n94), .B(n952), .Y(n92) );
  NAND2BXL U100 ( .AN(n952), .B(n94), .Y(n93) );
  INVX1 U101 ( .A(n750), .Y(n32) );
  OAI22X2 U102 ( .A0(n913), .A1(n89), .B0(n1031), .B1(n881), .Y(n17) );
  INVX1 U103 ( .A(n19), .Y(n12) );
  NOR2X1 U104 ( .A(n1013), .B(n1063), .Y(n53) );
  NOR2X1 U105 ( .A(n1226), .B(n324), .Y(n1167) );
  NOR2X1 U106 ( .A(n1226), .B(n300), .Y(n321) );
  NOR2X1 U107 ( .A(n1226), .B(n301), .Y(n352) );
  NOR2X1 U108 ( .A(n1226), .B(n1213), .Y(n1223) );
  NOR2X1 U109 ( .A(n1226), .B(n1202), .Y(n1217) );
  NOR2X1 U110 ( .A(n1226), .B(n308), .Y(n329) );
  NOR2X1 U111 ( .A(n1226), .B(n365), .Y(n386) );
  INVXL U112 ( .A(n854), .Y(n8) );
  NOR2X1 U113 ( .A(n1226), .B(n581), .Y(n631) );
  NOR2BX1 U114 ( .AN(n1124), .B(n1072), .Y(n222) );
  NOR2X1 U115 ( .A(n1226), .B(n344), .Y(n370) );
  INVX1 U116 ( .A(n1163), .Y(n74) );
  NOR2X1 U117 ( .A(n1030), .B(n630), .Y(n1076) );
  XNOR2X1 U118 ( .A(n1284), .B(n1283), .Y(PRODUCT[39]) );
  NAND2XL U119 ( .A(n132), .B(n546), .Y(n131) );
  NAND2XL U120 ( .A(n70), .B(n553), .Y(n558) );
  INVX4 U121 ( .A(n413), .Y(n681) );
  XOR2X1 U122 ( .A(n578), .B(n577), .Y(PRODUCT[19]) );
  XNOR2X1 U123 ( .A(n664), .B(n663), .Y(PRODUCT[17]) );
  NAND2X1 U124 ( .A(n144), .B(n664), .Y(n72) );
  NAND2X1 U125 ( .A(n517), .B(n516), .Y(n518) );
  INVX1 U126 ( .A(n544), .Y(n556) );
  BUFX2 U127 ( .A(A[15]), .Y(n990) );
  BUFX2 U128 ( .A(A[16]), .Y(n949) );
  BUFX2 U129 ( .A(A[8]), .Y(n972) );
  BUFX3 U130 ( .A(A[7]), .Y(n1014) );
  NAND2X1 U131 ( .A(n787), .B(n786), .Y(n1174) );
  XNOR2X1 U132 ( .A(n784), .B(n35), .Y(n279) );
  OR2X2 U133 ( .A(n36), .B(n785), .Y(n34) );
  NAND2X1 U134 ( .A(n36), .B(n785), .Y(n33) );
  INVXL U135 ( .A(n1137), .Y(n767) );
  NAND2XL U136 ( .A(n48), .B(n487), .Y(n47) );
  NAND2XL U137 ( .A(n429), .B(n430), .Y(n55) );
  XOR2X1 U138 ( .A(n252), .B(n42), .Y(n41) );
  NOR2X1 U139 ( .A(n200), .B(n199), .Y(n1263) );
  NAND2X1 U140 ( .A(n200), .B(n199), .Y(n1264) );
  INVX1 U141 ( .A(n894), .Y(n22) );
  NAND2BX1 U142 ( .AN(n854), .B(n9), .Y(n7) );
  XOR2X1 U143 ( .A(n487), .B(n51), .Y(n50) );
  OAI2BB1XL U144 ( .A0N(n1163), .A1N(n1162), .B0(n1161), .Y(n1181) );
  INVX1 U145 ( .A(n17), .Y(n16) );
  AND2X2 U146 ( .A(n96), .B(n737), .Y(n119) );
  OAI22X1 U147 ( .A0(n1162), .A1(n346), .B0(n1163), .B1(n341), .Y(n355) );
  NOR2X1 U148 ( .A(n1226), .B(n1186), .Y(n1199) );
  NOR2X1 U149 ( .A(n1226), .B(n1159), .Y(n1183) );
  INVXL U150 ( .A(n917), .Y(n15) );
  NOR2X1 U151 ( .A(n1030), .B(n984), .Y(n1023) );
  OR2XL U152 ( .A(n173), .B(n172), .Y(n1291) );
  XNOR2X1 U153 ( .A(n1249), .B(n1248), .Y(PRODUCT[36]) );
  XNOR2X1 U154 ( .A(n1256), .B(n1255), .Y(PRODUCT[37]) );
  XNOR2X1 U155 ( .A(n1271), .B(n1270), .Y(PRODUCT[38]) );
  AND2X2 U156 ( .A(n532), .B(n69), .Y(n68) );
  NAND3BX1 U157 ( .AN(n508), .B(n541), .C(n509), .Y(n69) );
  NAND2BX1 U158 ( .AN(n554), .B(n509), .Y(n70) );
  NOR2X1 U159 ( .A(n1303), .B(n1245), .Y(n1273) );
  NAND2X1 U160 ( .A(n566), .B(n565), .Y(n567) );
  XNOR2X1 U161 ( .A(n694), .B(n693), .Y(PRODUCT[16]) );
  INVX1 U162 ( .A(n949), .Y(n28) );
  INVX1 U163 ( .A(n539), .Y(n541) );
  NOR2X1 U164 ( .A(n571), .B(n1345), .Y(n287) );
  NAND2XL U165 ( .A(n1238), .B(n1336), .Y(n340) );
  AND2X1 U166 ( .A(n364), .B(n1338), .Y(n118) );
  BUFX2 U167 ( .A(A[18]), .Y(n947) );
  BUFX2 U168 ( .A(A[20]), .Y(n1158) );
  INVX1 U169 ( .A(n1335), .Y(n1238) );
  INVXL U170 ( .A(n1174), .Y(n1133) );
  INVXL U171 ( .A(n786), .Y(n82) );
  OAI2BB1X1 U172 ( .A0N(n34), .A1N(n784), .B0(n33), .Y(n786) );
  NAND2X1 U173 ( .A(n25), .B(n24), .Y(n868) );
  XNOR2X1 U174 ( .A(n1262), .B(n1261), .Y(n1397) );
  NAND2X1 U175 ( .A(n897), .B(n898), .Y(n24) );
  NOR2X1 U176 ( .A(n691), .B(n690), .Y(mult_x_1_n286) );
  NAND2X1 U177 ( .A(n766), .B(n765), .Y(n1137) );
  ADDFHX2 U178 ( .A(n844), .B(n843), .CI(n842), .CO(n803), .S(n845) );
  NOR2X1 U179 ( .A(n764), .B(n763), .Y(mult_x_1_n306) );
  ADDFHX2 U180 ( .A(n1055), .B(n1054), .CI(n1053), .CO(n1008), .S(n1056) );
  XNOR3X2 U181 ( .A(n898), .B(n897), .C(n26), .Y(n899) );
  INVXL U182 ( .A(n114), .Y(n113) );
  ADDFHX1 U183 ( .A(n866), .B(n865), .CI(n864), .CO(n846), .S(n867) );
  ADDFHX2 U184 ( .A(n256), .B(n255), .CI(n254), .CO(n257), .S(n238) );
  OAI2BB1X1 U185 ( .A0N(n993), .A1N(n65), .B0(n63), .Y(n1003) );
  OR2XL U186 ( .A(n1235), .B(n1234), .Y(n1237) );
  ADDFHX2 U187 ( .A(n484), .B(n483), .CI(n482), .CO(n498), .S(n804) );
  XOR2X1 U188 ( .A(n429), .B(n58), .Y(n57) );
  OAI2BB2X1 U189 ( .B0(n9), .B1(n8), .A0N(n7), .A1N(n853), .Y(n860) );
  NAND2X1 U190 ( .A(n895), .B(n894), .Y(n20) );
  XOR2X1 U191 ( .A(n488), .B(n50), .Y(n849) );
  INVX1 U192 ( .A(n430), .Y(n58) );
  INVX1 U193 ( .A(n42), .Y(n40) );
  ADDFHX1 U194 ( .A(n746), .B(n745), .CI(n744), .CO(n741), .S(n1127) );
  INVX1 U195 ( .A(n1109), .Y(n62) );
  NAND2XL U196 ( .A(n779), .B(n780), .Y(n104) );
  OAI21XL U197 ( .A0(n16), .A1(n15), .B0(n14), .Y(n926) );
  OAI2BB1XL U198 ( .A0N(n1072), .A1N(n214), .B0(n310), .Y(n327) );
  NAND2BX2 U199 ( .AN(n207), .B(n44), .Y(n43) );
  XOR2X1 U200 ( .A(n96), .B(n737), .Y(n31) );
  NAND2BXL U201 ( .AN(n719), .B(n110), .Y(n109) );
  INVXL U202 ( .A(n946), .Y(n95) );
  OR2X2 U203 ( .A(n189), .B(n188), .Y(n187) );
  NAND2XL U204 ( .A(B[7]), .B(n98), .Y(n146) );
  AND2XL U205 ( .A(n1297), .B(n1296), .Y(n1403) );
  XNOR2XL U206 ( .A(n1224), .B(n981), .Y(n324) );
  OR2XL U207 ( .A(n1295), .B(n1294), .Y(n1297) );
  XNOR2XL U208 ( .A(n1224), .B(A[24]), .Y(n1225) );
  XNOR2XL U209 ( .A(n1224), .B(n1212), .Y(n1213) );
  XNOR2XL U210 ( .A(n1224), .B(n1201), .Y(n1202) );
  XOR2X1 U211 ( .A(n127), .B(n340), .Y(PRODUCT[34]) );
  INVXL U212 ( .A(n1038), .Y(n110) );
  BUFX3 U213 ( .A(n155), .Y(n1038) );
  INVXL U214 ( .A(n1314), .Y(n124) );
  NAND2X1 U215 ( .A(B[1]), .B(n827), .Y(n170) );
  AND2X2 U216 ( .A(n535), .B(n534), .Y(n536) );
  INVXL U217 ( .A(n990), .Y(n11) );
  NAND2XL U218 ( .A(n123), .B(n1340), .Y(n122) );
  INVXL U219 ( .A(n1124), .Y(n98) );
  INVX1 U220 ( .A(n985), .Y(n76) );
  BUFX2 U221 ( .A(A[12]), .Y(n977) );
  BUFX2 U222 ( .A(A[10]), .Y(n945) );
  BUFX2 U223 ( .A(A[3]), .Y(n1028) );
  BUFX2 U224 ( .A(A[2]), .Y(n704) );
  BUFX2 U225 ( .A(A[1]), .Y(n640) );
  BUFX2 U226 ( .A(A[6]), .Y(n970) );
  BUFX2 U227 ( .A(A[4]), .Y(n983) );
  BUFX2 U228 ( .A(A[17]), .Y(n988) );
  BUFX2 U229 ( .A(A[23]), .Y(n1212) );
  BUFX2 U230 ( .A(A[22]), .Y(n1201) );
  BUFX2 U231 ( .A(A[19]), .Y(n981) );
  OAI22X1 U232 ( .A0(n89), .A1(n606), .B0(n605), .B1(n1163), .Y(n613) );
  INVX1 U233 ( .A(n476), .Y(n487) );
  INVX1 U234 ( .A(B[3]), .Y(n413) );
  OAI21XL U235 ( .A0(n1136), .A1(n1135), .B0(n1134), .Y(mult_x_1_n309) );
  OAI22X1 U236 ( .A0(n214), .A1(n260), .B0(n1072), .B1(n736), .Y(n749) );
  XOR2X2 U237 ( .A(B[8]), .B(B[9]), .Y(n205) );
  BUFX8 U238 ( .A(n456), .Y(n1065) );
  XNOR2X1 U239 ( .A(n986), .B(A[13]), .Y(n881) );
  NOR2BX1 U240 ( .AN(n1124), .B(n1067), .Y(n740) );
  OAI22X1 U241 ( .A0(n1033), .A1(n597), .B0(n1031), .B1(n1032), .Y(n1080) );
  OAI22X1 U242 ( .A0(n881), .A1(n1162), .B0(n19), .B1(n1163), .Y(n886) );
  XOR2X1 U243 ( .A(n1360), .B(n1356), .Y(PRODUCT[13]) );
  OAI22X1 U244 ( .A0(n214), .A1(n594), .B0(n1072), .B1(n593), .Y(n603) );
  XOR2X2 U245 ( .A(B[12]), .B(n1187), .Y(n299) );
  OAI22X1 U246 ( .A0(n1205), .A1(n626), .B0(n1067), .B1(n1068), .Y(n1099) );
  OAI22X1 U247 ( .A0(n214), .A1(n307), .B0(n1072), .B1(n215), .Y(n248) );
  NOR2X1 U248 ( .A(n258), .B(n257), .Y(n788) );
  BUFX3 U249 ( .A(n1033), .Y(n89) );
  XNOR3X2 U250 ( .A(n854), .B(n9), .C(n853), .Y(n894) );
  AOI21X2 U251 ( .A0(n5), .A1(n12), .B0(n10), .Y(n9) );
  NOR2X1 U252 ( .A(n817), .B(n1163), .Y(n10) );
  XOR2X1 U253 ( .A(n986), .B(n11), .Y(n817) );
  NAND2X4 U254 ( .A(n13), .B(n1031), .Y(n1033) );
  XNOR2X4 U255 ( .A(B[10]), .B(B[9]), .Y(n1031) );
  XOR2X2 U256 ( .A(B[11]), .B(B[10]), .Y(n13) );
  OAI21XL U257 ( .A0(n917), .A1(n17), .B0(n916), .Y(n14) );
  XOR3X2 U258 ( .A(n917), .B(n17), .C(n916), .Y(n960) );
  XOR3X2 U259 ( .A(n18), .B(n1143), .C(n1142), .Y(n1150) );
  XOR2X1 U260 ( .A(n986), .B(n97), .Y(n19) );
  OAI2BB1X1 U261 ( .A0N(n893), .A1N(n21), .B0(n20), .Y(n898) );
  INVX1 U262 ( .A(n895), .Y(n23) );
  XOR3X2 U263 ( .A(n895), .B(n894), .C(n893), .Y(n927) );
  INVX1 U264 ( .A(n896), .Y(n26) );
  OAI21XL U265 ( .A0(n897), .A1(n898), .B0(n896), .Y(n25) );
  OAI22X1 U266 ( .A0(n817), .A1(n1162), .B0(n1163), .B1(n27), .Y(n823) );
  OAI22X1 U267 ( .A0(n1163), .A1(n479), .B0(n1162), .B1(n27), .Y(n490) );
  NAND2X1 U268 ( .A(n764), .B(n763), .Y(mult_x_1_n307) );
  OAI22X1 U269 ( .A0(n1162), .A1(n306), .B0(n1163), .B1(n262), .Y(n96) );
  OAI21X2 U270 ( .A0(n32), .A1(n30), .B0(n29), .Y(n782) );
  INVX1 U271 ( .A(n749), .Y(n30) );
  XNOR3X2 U272 ( .A(n749), .B(n32), .C(n31), .Y(n785) );
  XNOR2X1 U273 ( .A(n36), .B(n785), .Y(n35) );
  OR2X2 U274 ( .A(n85), .B(n86), .Y(n37) );
  OAI2BB1X1 U275 ( .A0N(n253), .A1N(n42), .B0(n38), .Y(n263) );
  NAND2BX1 U276 ( .AN(n253), .B(n40), .Y(n39) );
  XOR2X1 U277 ( .A(n253), .B(n41), .Y(n256) );
  INVX1 U278 ( .A(n214), .Y(n44) );
  XOR2X1 U279 ( .A(n45), .B(n263), .Y(n275) );
  XNOR2X1 U280 ( .A(n264), .B(n86), .Y(n45) );
  XOR2X1 U281 ( .A(n46), .B(n1097), .Y(mult_x_1_n618) );
  XOR2X1 U282 ( .A(n1096), .B(n1098), .Y(n46) );
  OAI2BB1X1 U283 ( .A0N(n488), .A1N(n51), .B0(n47), .Y(n497) );
  NAND2BX1 U284 ( .AN(n488), .B(n49), .Y(n48) );
  INVXL U285 ( .A(n51), .Y(n49) );
  OAI22X4 U286 ( .A0(n1205), .A1(n808), .B0(n1206), .B1(n473), .Y(n51) );
  NAND2X1 U287 ( .A(n52), .B(n1070), .Y(n137) );
  INVX1 U288 ( .A(n139), .Y(n52) );
  XNOR2X2 U289 ( .A(n1070), .B(n139), .Y(n140) );
  NOR2X2 U290 ( .A(n54), .B(n53), .Y(n139) );
  OAI21XL U291 ( .A0(n1097), .A1(n1098), .B0(n1096), .Y(n136) );
  OAI2BB1X1 U292 ( .A0N(n56), .A1N(n428), .B0(n55), .Y(n432) );
  NAND2BX1 U293 ( .AN(n429), .B(n58), .Y(n56) );
  XNOR2X1 U294 ( .A(n428), .B(n57), .Y(n442) );
  CLKINVX3 U295 ( .A(B[5]), .Y(n157) );
  OAI21XL U296 ( .A0(n264), .A1(n265), .B0(n263), .Y(n59) );
  NOR2X1 U297 ( .A(n279), .B(n278), .Y(n772) );
  INVX1 U298 ( .A(n66), .Y(n64) );
  NAND2BX1 U299 ( .AN(n994), .B(n66), .Y(n65) );
  XNOR3X2 U300 ( .A(n994), .B(n66), .C(n993), .Y(n1051) );
  AOI2BB1X2 U301 ( .A0N(n89), .A1N(n987), .B0(n67), .Y(n66) );
  NOR2X1 U302 ( .A(n946), .B(n1031), .Y(n67) );
  NOR3BX2 U303 ( .AN(n570), .B(n571), .C(n1345), .Y(n144) );
  NOR2X2 U304 ( .A(n1349), .B(n1347), .Y(n570) );
  NOR2X1 U305 ( .A(n559), .B(n564), .Y(n551) );
  NOR2X4 U306 ( .A(n1378), .B(n1377), .Y(n564) );
  NOR2X2 U307 ( .A(n1376), .B(n1375), .Y(n559) );
  INVX1 U308 ( .A(n508), .Y(n537) );
  CLKINVX3 U309 ( .A(n509), .Y(n568) );
  XNOR2X2 U310 ( .A(n68), .B(n536), .Y(PRODUCT[26]) );
  NAND2X4 U311 ( .A(n72), .B(n71), .Y(n509) );
  AOI21X2 U312 ( .A0(n287), .A1(n569), .B0(n99), .Y(n71) );
  INVX4 U313 ( .A(B[11]), .Y(n306) );
  OAI22X1 U314 ( .A0(n1032), .A1(n89), .B0(n1163), .B1(n75), .Y(n1083) );
  XNOR2X2 U315 ( .A(B[6]), .B(B[5]), .Y(n147) );
  INVX4 U316 ( .A(n1353), .Y(n129) );
  OAI21XL U317 ( .A0(n929), .A1(n928), .B0(n927), .Y(n142) );
  BUFX2 U318 ( .A(n1146), .Y(n77) );
  NAND2X1 U319 ( .A(n77), .B(n1145), .Y(n78) );
  INVX1 U320 ( .A(n1145), .Y(n80) );
  XNOR3X2 U321 ( .A(n1145), .B(n81), .C(n1144), .Y(n1147) );
  INVX1 U322 ( .A(n1146), .Y(n81) );
  NAND2XL U323 ( .A(n1173), .B(n1175), .Y(n1135) );
  NAND2X1 U324 ( .A(n83), .B(n82), .Y(n1175) );
  NAND2BX2 U325 ( .AN(n1132), .B(n84), .Y(n1173) );
  INVX1 U326 ( .A(n264), .Y(n85) );
  INVX1 U327 ( .A(n265), .Y(n86) );
  NAND2X1 U328 ( .A(n1142), .B(n1143), .Y(n87) );
  INVX1 U329 ( .A(n1033), .Y(n103) );
  NAND2X1 U330 ( .A(n90), .B(n748), .Y(n100) );
  OAI21XL U331 ( .A0(n90), .A1(n748), .B0(n747), .Y(n101) );
  XOR3X2 U332 ( .A(n747), .B(n90), .C(n748), .Y(n778) );
  OAI21XL U333 ( .A0(n1006), .A1(n1005), .B0(n1004), .Y(n91) );
  XOR3X2 U334 ( .A(n1004), .B(n1005), .C(n1006), .Y(n1007) );
  XNOR3X2 U335 ( .A(n952), .B(n94), .C(n951), .Y(n1002) );
  AOI2BB2X2 U336 ( .B0(n95), .B1(n5), .A0N(n913), .A1N(n1031), .Y(n94) );
  NAND2X1 U337 ( .A(n1172), .B(n1174), .Y(n108) );
  NAND2X1 U338 ( .A(n1132), .B(n1131), .Y(n1172) );
  INVX1 U339 ( .A(n968), .Y(n97) );
  XOR3X2 U340 ( .A(n927), .B(n928), .C(n929), .Y(n930) );
  XOR2X1 U341 ( .A(n302), .B(A[13]), .Y(n1059) );
  XOR2X1 U342 ( .A(n302), .B(n977), .Y(n1060) );
  XOR2X1 U343 ( .A(n302), .B(n640), .Y(n219) );
  XOR2X1 U344 ( .A(n302), .B(n1028), .Y(n242) );
  XOR2X1 U345 ( .A(n302), .B(n1124), .Y(n151) );
  XOR2X1 U346 ( .A(n302), .B(n1185), .Y(n454) );
  XOR2X1 U347 ( .A(n302), .B(n704), .Y(n218) );
  XOR2X1 U348 ( .A(n302), .B(n988), .Y(n902) );
  XOR2X1 U349 ( .A(n302), .B(n968), .Y(n1010) );
  XOR2X1 U350 ( .A(n302), .B(n1020), .Y(n627) );
  XOR2X1 U351 ( .A(n302), .B(n981), .Y(n833) );
  XOR2X1 U352 ( .A(n302), .B(n949), .Y(n933) );
  XOR2X1 U353 ( .A(n302), .B(n1158), .Y(n480) );
  XOR2X1 U354 ( .A(n302), .B(n983), .Y(n272) );
  XOR2X1 U355 ( .A(n302), .B(n990), .Y(n969) );
  XOR2X1 U356 ( .A(n302), .B(n1012), .Y(n716) );
  XOR2X1 U357 ( .A(n302), .B(n1212), .Y(n382) );
  XOR2X1 U358 ( .A(n302), .B(n947), .Y(n870) );
  XOR2X1 U359 ( .A(n302), .B(n972), .Y(n653) );
  XOR2X1 U360 ( .A(n302), .B(A[25]), .Y(n303) );
  XOR2X1 U361 ( .A(n302), .B(n1201), .Y(n418) );
  XOR2X1 U362 ( .A(n302), .B(n970), .Y(n715) );
  XOR2X1 U363 ( .A(n302), .B(A[24]), .Y(n374) );
  XOR2X1 U364 ( .A(n302), .B(n1014), .Y(n701) );
  XOR2X1 U365 ( .A(n302), .B(n945), .Y(n607) );
  XNOR2X1 U366 ( .A(B[15]), .B(B[16]), .Y(n380) );
  OAI21X1 U367 ( .A0(n571), .A1(n1346), .B0(n572), .Y(n99) );
  NAND2X1 U368 ( .A(n1379), .B(n1380), .Y(n572) );
  OAI21X1 U369 ( .A0(n1350), .A1(n1347), .B0(n1348), .Y(n569) );
  NAND2X1 U370 ( .A(n101), .B(n100), .Y(n783) );
  NAND2BX2 U371 ( .AN(n273), .B(n103), .Y(n102) );
  NAND2X1 U372 ( .A(n105), .B(n104), .Y(n1129) );
  OR2X2 U373 ( .A(n779), .B(n780), .Y(n106) );
  XOR2X1 U374 ( .A(n779), .B(n107), .Y(n784) );
  XOR2X1 U375 ( .A(n778), .B(n780), .Y(n107) );
  XNOR2X1 U376 ( .A(B[4]), .B(B[3]), .Y(n155) );
  NAND2X1 U377 ( .A(n108), .B(n1173), .Y(n1134) );
  OAI22X1 U378 ( .A0(n259), .A1(n1040), .B0(n155), .B1(n111), .Y(n750) );
  OAI21XL U379 ( .A0(n1040), .A1(n111), .B0(n109), .Y(n751) );
  XNOR2X1 U380 ( .A(n991), .B(n1014), .Y(n111) );
  NAND2X1 U381 ( .A(n691), .B(n690), .Y(mult_x_1_n287) );
  OAI2BB1X2 U382 ( .A0N(n657), .A1N(n113), .B0(n112), .Y(n1151) );
  NAND2X1 U383 ( .A(n658), .B(n659), .Y(n112) );
  NOR2X1 U384 ( .A(n658), .B(n659), .Y(n114) );
  XOR3X2 U385 ( .A(n659), .B(n658), .C(n657), .Y(n665) );
  NAND2XL U386 ( .A(n354), .B(n355), .Y(n115) );
  OR2X1 U387 ( .A(n354), .B(n355), .Y(n116) );
  XOR3X2 U388 ( .A(n355), .B(n354), .C(n353), .Y(n390) );
  OAI22X2 U389 ( .A0(n1040), .A1(n625), .B0(n1038), .B1(n1039), .Y(n1100) );
  OAI22X1 U390 ( .A0(n1061), .A1(n1060), .B0(n1011), .B1(n1059), .Y(n1104) );
  OAI22X1 U391 ( .A0(n1205), .A1(n1068), .B0(n1067), .B1(n1066), .Y(n1102) );
  OAI21X2 U392 ( .A0(n565), .A1(n559), .B0(n560), .Y(n552) );
  NAND2X4 U393 ( .A(n1378), .B(n1377), .Y(n565) );
  NAND2X1 U394 ( .A(n1376), .B(n1375), .Y(n560) );
  OAI22X1 U395 ( .A0(n1205), .A1(n378), .B0(n1206), .B1(n342), .Y(n373) );
  XNOR2X1 U396 ( .A(n681), .B(n1201), .Y(n851) );
  XNOR2X1 U397 ( .A(n681), .B(n945), .Y(n717) );
  OAI22X2 U398 ( .A0(n1065), .A1(n1064), .B0(n1063), .B1(n1062), .Y(n1103) );
  INVX8 U399 ( .A(n584), .Y(n1214) );
  INVX4 U400 ( .A(B[15]), .Y(n584) );
  BUFX3 U401 ( .A(n380), .Y(n1226) );
  XNOR2XL U402 ( .A(n991), .B(A[25]), .Y(n366) );
  OAI21XL U403 ( .A0(n1343), .A1(n504), .B0(n1344), .Y(n436) );
  NAND2XL U404 ( .A(n1238), .B(n1240), .Y(n1243) );
  AOI21XL U405 ( .A0(n1279), .A1(n1251), .B0(n1250), .Y(n1252) );
  INVXL U406 ( .A(n1332), .Y(n1250) );
  INVX1 U407 ( .A(n1359), .Y(n769) );
  XNOR2XL U408 ( .A(n991), .B(A[24]), .Y(n416) );
  BUFX3 U409 ( .A(A[14]), .Y(n968) );
  XNOR2XL U410 ( .A(n1214), .B(n981), .Y(n311) );
  BUFX3 U411 ( .A(A[5]), .Y(n1012) );
  BUFX3 U412 ( .A(A[9]), .Y(n985) );
  XNOR2XL U413 ( .A(n991), .B(n985), .Y(n683) );
  XNOR2XL U414 ( .A(n1021), .B(n1012), .Y(n680) );
  BUFX3 U415 ( .A(A[11]), .Y(n1020) );
  NAND2XL U416 ( .A(n1251), .B(n1332), .Y(n1248) );
  NAND2XL U417 ( .A(n1240), .B(n1334), .Y(n297) );
  OAI21XL U418 ( .A0(n1314), .A1(n296), .B0(n295), .Y(n298) );
  OR2XL U419 ( .A(n1339), .B(n1342), .Y(n123) );
  NOR2X1 U420 ( .A(n1339), .B(n1341), .Y(n294) );
  NOR2XL U421 ( .A(n1243), .B(n1337), .Y(n1302) );
  NOR2XL U422 ( .A(n1301), .B(n1325), .Y(n1306) );
  OAI21XL U423 ( .A0(n548), .A1(n555), .B0(n549), .Y(n288) );
  XNOR2X1 U424 ( .A(n575), .B(n574), .Y(PRODUCT[20]) );
  NAND2XL U425 ( .A(n573), .B(n572), .Y(n574) );
  OAI21XL U426 ( .A0(n578), .A1(n1345), .B0(n1346), .Y(n575) );
  AOI21X1 U427 ( .A0(n664), .A1(n662), .B0(n283), .Y(n286) );
  BUFX3 U428 ( .A(n580), .Y(n1067) );
  XNOR2XL U429 ( .A(n1214), .B(n1185), .Y(n1165) );
  XNOR2XL U430 ( .A(n1214), .B(n1158), .Y(n323) );
  CMPR32X1 U431 ( .A(n679), .B(n678), .C(n677), .CO(n674), .S(n728) );
  OAI22XL U432 ( .A0(n1027), .A1(n654), .B0(n639), .B1(n827), .Y(n678) );
  NOR2BX1 U433 ( .AN(n1124), .B(n1063), .Y(n679) );
  OAI22XL U434 ( .A0(n1205), .A1(n702), .B0(n1067), .B1(n641), .Y(n677) );
  INVX4 U435 ( .A(n157), .Y(n991) );
  NAND2XL U436 ( .A(n1275), .B(n1328), .Y(n1270) );
  XNOR2XL U437 ( .A(n1214), .B(A[24]), .Y(n1215) );
  XNOR2XL U438 ( .A(n1214), .B(n1212), .Y(n1197) );
  OAI22XL U439 ( .A0(n1229), .A1(n1215), .B0(n1230), .B1(n1227), .Y(n1233) );
  INVXL U440 ( .A(n1331), .Y(n1251) );
  INVXL U441 ( .A(n1337), .Y(n364) );
  INVXL U442 ( .A(n1342), .Y(n399) );
  NAND2XL U443 ( .A(n398), .B(n439), .Y(n401) );
  INVXL U444 ( .A(n1339), .Y(n402) );
  INVXL U445 ( .A(n398), .Y(n438) );
  INVXL U446 ( .A(n436), .Y(n437) );
  INVXL U447 ( .A(n1341), .Y(n439) );
  INVXL U448 ( .A(n1336), .Y(n1241) );
  INVXL U449 ( .A(n1333), .Y(n1240) );
  NAND2XL U450 ( .A(n1273), .B(n1251), .Y(n1253) );
  INVXL U451 ( .A(n1329), .Y(n1254) );
  INVXL U452 ( .A(n1343), .Y(n470) );
  NOR2XL U453 ( .A(n1362), .B(n1361), .Y(n503) );
  NAND2X1 U454 ( .A(n1361), .B(n1362), .Y(n504) );
  NAND2BX1 U455 ( .AN(n547), .B(n509), .Y(n132) );
  AOI21XL U456 ( .A0(n552), .A1(n556), .B0(n545), .Y(n546) );
  XNOR2XL U457 ( .A(n1021), .B(n640), .Y(n251) );
  NAND2BX1 U458 ( .AN(n1124), .B(n986), .Y(n262) );
  XNOR2X1 U459 ( .A(n1021), .B(n1028), .Y(n736) );
  OR2X2 U460 ( .A(n375), .B(n1230), .Y(n120) );
  INVXL U461 ( .A(n366), .Y(n367) );
  XNOR2XL U462 ( .A(n1214), .B(n949), .Y(n375) );
  XNOR2XL U463 ( .A(n1214), .B(n988), .Y(n345) );
  XNOR2XL U464 ( .A(n1214), .B(n947), .Y(n315) );
  XNOR2XL U465 ( .A(n1021), .B(n970), .Y(n645) );
  XNOR2XL U466 ( .A(n1187), .B(n640), .Y(n702) );
  XNOR2X1 U467 ( .A(n1021), .B(n1014), .Y(n594) );
  XNOR2X1 U468 ( .A(n986), .B(n970), .Y(n605) );
  INVXL U469 ( .A(n1307), .Y(n1244) );
  INVXL U470 ( .A(n1301), .Y(n1278) );
  XOR2X1 U471 ( .A(n769), .B(n1355), .Y(PRODUCT[14]) );
  OAI22XL U472 ( .A0(n1027), .A1(n711), .B0(n654), .B1(n1123), .Y(n710) );
  OAI22XL U473 ( .A0(n1205), .A1(n656), .B0(n1206), .B1(n655), .Y(n709) );
  INVXL U474 ( .A(n1187), .Y(n656) );
  OAI22XL U475 ( .A0(n1033), .A1(n714), .B0(n1031), .B1(n713), .Y(n738) );
  OAI22XL U476 ( .A0(n170), .A1(n712), .B0(n711), .B1(n1123), .Y(n739) );
  OAI22XL U477 ( .A0(n1061), .A1(n716), .B0(n1011), .B1(n715), .Y(n753) );
  OAI22XL U478 ( .A0(n6), .A1(n718), .B0(n1035), .B1(n717), .Y(n752) );
  INVXL U479 ( .A(n1160), .Y(n1161) );
  CMPR32X1 U480 ( .A(n424), .B(n423), .C(n422), .CO(n408), .S(n466) );
  NOR2XL U481 ( .A(n1030), .B(n381), .Y(n423) );
  OAI22X1 U482 ( .A0(n1205), .A1(n420), .B0(n1206), .B1(n379), .Y(n424) );
  OAI22XL U483 ( .A0(n1061), .A1(n833), .B0(n1011), .B1(n480), .Y(n816) );
  INVXL U484 ( .A(n813), .Y(n486) );
  XNOR2X1 U485 ( .A(n1214), .B(n1020), .Y(n834) );
  XNOR2X1 U486 ( .A(n1187), .B(A[13]), .Y(n835) );
  OAI22XL U487 ( .A0(n1027), .A1(n1026), .B0(n1025), .B1(n1123), .Y(n1075) );
  XNOR2XL U488 ( .A(n1021), .B(n945), .Y(n1073) );
  XNOR2XL U489 ( .A(n1021), .B(n985), .Y(n624) );
  XNOR2X1 U490 ( .A(n1021), .B(n972), .Y(n593) );
  XNOR2XL U491 ( .A(n986), .B(n972), .Y(n1032) );
  OAI22XL U492 ( .A0(n1162), .A1(n313), .B0(n1163), .B1(n325), .Y(n330) );
  OAI22XL U493 ( .A0(n1229), .A1(n311), .B0(n1230), .B1(n323), .Y(n332) );
  OAI22XL U494 ( .A0(n1205), .A1(n312), .B0(n1206), .B1(n326), .Y(n331) );
  INVXL U495 ( .A(n309), .Y(n310) );
  BUFX8 U496 ( .A(n1033), .Y(n1162) );
  INVXL U497 ( .A(n303), .Y(n304) );
  OAI22XL U498 ( .A0(n1040), .A1(n719), .B0(n1038), .B1(n683), .Y(n732) );
  OAI22XL U499 ( .A0(n214), .A1(n735), .B0(n1072), .B1(n680), .Y(n734) );
  AOI21XL U500 ( .A0(n1307), .A1(n1306), .B0(n1305), .Y(n1308) );
  NAND2XL U501 ( .A(n1302), .B(n1306), .Y(n1309) );
  AOI21XL U502 ( .A0(n1279), .A1(n1278), .B0(n1277), .Y(n1280) );
  INVXL U503 ( .A(n1304), .Y(n1277) );
  NAND2XL U504 ( .A(n1273), .B(n1278), .Y(n1281) );
  INVXL U505 ( .A(n1325), .Y(n1282) );
  NOR2X2 U506 ( .A(n293), .B(n508), .Y(n126) );
  NAND2X1 U507 ( .A(n507), .B(n291), .Y(n293) );
  OAI22XL U508 ( .A0(n1229), .A1(n1184), .B0(n1230), .B1(n1197), .Y(n1200) );
  INVXL U509 ( .A(n1218), .Y(n1198) );
  OAI22XL U510 ( .A0(n1229), .A1(n1165), .B0(n1230), .B1(n1184), .Y(n1190) );
  OAI22XL U511 ( .A0(n1205), .A1(n1164), .B0(n1206), .B1(n1188), .Y(n1191) );
  AOI21XL U512 ( .A0(n796), .A1(n794), .B0(n239), .Y(n240) );
  NAND2X1 U513 ( .A(n796), .B(n800), .Y(n241) );
  OAI22XL U514 ( .A0(n214), .A1(n419), .B0(n1072), .B1(n411), .Y(n453) );
  OAI22XL U515 ( .A0(n214), .A1(n908), .B0(n1072), .B1(n876), .Y(n889) );
  ADDFX2 U516 ( .A(n886), .B(n885), .CI(n884), .CO(n895), .S(n925) );
  OAI22XL U517 ( .A0(n1040), .A1(n883), .B0(n1038), .B1(n852), .Y(n884) );
  OAI22XL U518 ( .A0(n6), .A1(n882), .B0(n1035), .B1(n851), .Y(n885) );
  OAI22X1 U519 ( .A0(n1065), .A1(n1013), .B0(n1063), .B1(n971), .Y(n1018) );
  OAI22XL U520 ( .A0(n1061), .A1(n653), .B0(n1011), .B1(n608), .Y(n671) );
  OAI22XL U521 ( .A0(n6), .A1(n647), .B0(n1035), .B1(n600), .Y(n673) );
  OAI22XL U522 ( .A0(n89), .A1(n646), .B0(n1163), .B1(n606), .Y(n672) );
  OAI22XL U523 ( .A0(n1040), .A1(n651), .B0(n1038), .B1(n636), .Y(n676) );
  NOR2BXL U524 ( .AN(n1124), .B(n1035), .Y(n172) );
  OAI22XL U525 ( .A0(n1027), .A1(n169), .B0(n175), .B1(n1123), .Y(n173) );
  OAI22XL U526 ( .A0(n6), .A1(n184), .B0(n1035), .B1(n183), .Y(n194) );
  OAI22XL U527 ( .A0(n1027), .A1(n182), .B0(n181), .B1(n1123), .Y(n195) );
  NOR2BXL U528 ( .AN(n1124), .B(n1038), .Y(n196) );
  OAI22XL U529 ( .A0(n6), .A1(n183), .B0(n1035), .B1(n164), .Y(n193) );
  OAI22XL U530 ( .A0(n6), .A1(n164), .B0(n1035), .B1(n153), .Y(n163) );
  OR2X2 U531 ( .A(n238), .B(n237), .Y(n796) );
  NAND2X1 U532 ( .A(n257), .B(n258), .Y(n789) );
  OAI2BB1XL U533 ( .A0N(n1230), .A1N(n1229), .B0(n1228), .Y(n1231) );
  INVXL U534 ( .A(n1227), .Y(n1228) );
  NOR2XL U535 ( .A(n1226), .B(n1225), .Y(n1232) );
  INVXL U536 ( .A(n1233), .Y(n1222) );
  ADDFX2 U537 ( .A(n926), .B(n925), .CI(n924), .CO(n929), .S(n962) );
  OAI22XL U538 ( .A0(n1027), .A1(n1124), .B0(n169), .B1(n1123), .Y(n1295) );
  NAND2XL U539 ( .A(n171), .B(n1027), .Y(n1294) );
  NAND2BXL U540 ( .AN(n1124), .B(B[1]), .Y(n171) );
  NAND2XL U541 ( .A(n1295), .B(n1294), .Y(n1296) );
  NAND2XL U542 ( .A(n173), .B(n172), .Y(n1290) );
  INVXL U543 ( .A(n1296), .Y(n1292) );
  NOR2XL U544 ( .A(n180), .B(n179), .Y(n1285) );
  NAND2XL U545 ( .A(n180), .B(n179), .Y(n1286) );
  AOI21XL U546 ( .A0(n1291), .A1(n1292), .B0(n174), .Y(n1288) );
  INVXL U547 ( .A(n1290), .Y(n174) );
  NAND2XL U548 ( .A(n198), .B(n197), .Y(n1317) );
  INVXL U549 ( .A(n1257), .Y(n1266) );
  INVXL U550 ( .A(n507), .Y(n520) );
  NOR2X1 U551 ( .A(n520), .B(n525), .Y(n512) );
  INVXL U552 ( .A(n1279), .Y(n1246) );
  INVXL U553 ( .A(n1273), .Y(n1247) );
  OAI21XL U554 ( .A0(n1310), .A1(n1337), .B0(n1338), .Y(n339) );
  NOR2XL U555 ( .A(n1331), .B(n1329), .Y(n1272) );
  INVXL U556 ( .A(n1302), .Y(n1245) );
  NAND2XL U557 ( .A(n1272), .B(n1275), .Y(n1301) );
  AOI21XL U558 ( .A0(n531), .A1(n512), .B0(n511), .Y(n513) );
  OAI21XL U559 ( .A0(n521), .A1(n525), .B0(n526), .Y(n511) );
  INVXL U560 ( .A(n510), .Y(n521) );
  INVXL U561 ( .A(n515), .Y(n517) );
  NAND2XL U562 ( .A(n537), .B(n522), .Y(n524) );
  AOI21XL U563 ( .A0(n531), .A1(n522), .B0(n510), .Y(n523) );
  AOI21XL U564 ( .A0(n531), .A1(n541), .B0(n530), .Y(n532) );
  INVXL U565 ( .A(n533), .Y(n535) );
  INVXL U566 ( .A(n1350), .Y(n283) );
  INVX1 U567 ( .A(n1349), .Y(n662) );
  XNOR2XL U568 ( .A(n1323), .B(n1357), .Y(PRODUCT[12]) );
  XNOR2XL U569 ( .A(n986), .B(n1124), .Y(n273) );
  NAND2BXL U570 ( .AN(n1124), .B(n1187), .Y(n655) );
  XNOR2XL U571 ( .A(n681), .B(n985), .Y(n718) );
  XNOR2XL U572 ( .A(n1214), .B(n1124), .Y(n589) );
  NAND2BX1 U573 ( .AN(n1124), .B(n1021), .Y(n215) );
  OAI22XL U574 ( .A0(n214), .A1(n251), .B0(n1072), .B1(n260), .Y(n266) );
  XNOR2XL U575 ( .A(n1224), .B(n947), .Y(n308) );
  XNOR2XL U576 ( .A(n1224), .B(n949), .Y(n301) );
  XNOR2XL U577 ( .A(n991), .B(n972), .Y(n719) );
  XNOR2XL U578 ( .A(n991), .B(n704), .Y(n152) );
  XNOR2XL U579 ( .A(n681), .B(n1012), .Y(n208) );
  XNOR2XL U580 ( .A(n681), .B(n970), .Y(n213) );
  XNOR2XL U581 ( .A(n991), .B(n1028), .Y(n210) );
  XNOR2XL U582 ( .A(n991), .B(n983), .Y(n209) );
  XNOR2X1 U583 ( .A(n404), .B(n403), .Y(PRODUCT[32]) );
  NAND2XL U584 ( .A(n402), .B(n1340), .Y(n403) );
  OAI21XL U585 ( .A0(n1314), .A1(n401), .B0(n400), .Y(n404) );
  XNOR2X1 U586 ( .A(n441), .B(n440), .Y(PRODUCT[31]) );
  NAND2XL U587 ( .A(n439), .B(n1342), .Y(n440) );
  OAI21XL U588 ( .A0(n1314), .A1(n438), .B0(n437), .Y(n441) );
  AOI21XL U589 ( .A0(n1241), .A1(n1240), .B0(n1239), .Y(n1242) );
  INVXL U590 ( .A(n1334), .Y(n1239) );
  AOI21XL U591 ( .A0(n1279), .A1(n1272), .B0(n1276), .Y(n1268) );
  NAND2XL U592 ( .A(n1273), .B(n1272), .Y(n1269) );
  INVXL U593 ( .A(n1327), .Y(n1275) );
  AOI21XL U594 ( .A0(n1276), .A1(n1275), .B0(n1274), .Y(n1304) );
  INVXL U595 ( .A(n1328), .Y(n1274) );
  NOR2XL U596 ( .A(n539), .B(n533), .Y(n507) );
  AOI21X1 U597 ( .A0(n291), .A1(n510), .B0(n290), .Y(n292) );
  NAND2XL U598 ( .A(n1254), .B(n1330), .Y(n1255) );
  XNOR2X1 U599 ( .A(n472), .B(n471), .Y(PRODUCT[30]) );
  NAND2XL U600 ( .A(n470), .B(n1344), .Y(n471) );
  XOR2X1 U601 ( .A(n1314), .B(n506), .Y(PRODUCT[29]) );
  NAND2XL U602 ( .A(n505), .B(n504), .Y(n506) );
  INVXL U603 ( .A(n503), .Y(n505) );
  XNOR2X1 U604 ( .A(n543), .B(n542), .Y(PRODUCT[25]) );
  NAND2XL U605 ( .A(n541), .B(n540), .Y(n542) );
  XOR2X1 U606 ( .A(n131), .B(n117), .Y(PRODUCT[24]) );
  AND2XL U607 ( .A(n550), .B(n549), .Y(n117) );
  NAND2XL U608 ( .A(n662), .B(n1350), .Y(n663) );
  OAI22XL U609 ( .A0(n6), .A1(n244), .B0(n1035), .B1(n274), .Y(n269) );
  OAI22XL U610 ( .A0(n1061), .A1(n242), .B0(n1011), .B1(n272), .Y(n271) );
  OAI22XL U611 ( .A0(n652), .A1(n243), .B0(n1038), .B1(n259), .Y(n270) );
  OAI22XL U612 ( .A0(n652), .A1(n209), .B0(n1038), .B1(n243), .Y(n252) );
  OAI22XL U613 ( .A0(n1061), .A1(n218), .B0(n1011), .B1(n242), .Y(n253) );
  INVXL U614 ( .A(n1203), .Y(n1204) );
  XNOR2XL U615 ( .A(n1224), .B(n1185), .Y(n1186) );
  XNOR2XL U616 ( .A(n1214), .B(n1201), .Y(n1184) );
  OAI22XL U617 ( .A0(n1033), .A1(n713), .B0(n1031), .B1(n705), .Y(n729) );
  OAI22XL U618 ( .A0(n1061), .A1(n715), .B0(n1011), .B1(n701), .Y(n731) );
  OAI22XL U619 ( .A0(n1205), .A1(n703), .B0(n1067), .B1(n702), .Y(n730) );
  OAI22XL U620 ( .A0(n652), .A1(n683), .B0(n1038), .B1(n651), .Y(n708) );
  OAI22XL U621 ( .A0(n1061), .A1(n701), .B0(n1011), .B1(n653), .Y(n707) );
  CMPR32X1 U622 ( .A(n650), .B(n649), .C(n648), .CO(n642), .S(n699) );
  OAI22XL U623 ( .A0(n214), .A1(n645), .B0(n1072), .B1(n594), .Y(n650) );
  OAI22XL U624 ( .A0(n1205), .A1(n641), .B0(n1067), .B1(n596), .Y(n648) );
  OAI22XL U625 ( .A0(n1065), .A1(n589), .B0(n1063), .B1(n588), .Y(n649) );
  ADDFX2 U626 ( .A(n777), .B(n119), .CI(n776), .CO(n754), .S(n1130) );
  XNOR2XL U627 ( .A(n1021), .B(n1158), .Y(n419) );
  ADDFX2 U628 ( .A(n427), .B(n426), .CI(n425), .CO(n447), .S(n465) );
  OAI22XL U629 ( .A0(n1061), .A1(n418), .B0(n1011), .B1(n382), .Y(n427) );
  OAI22XL U630 ( .A0(n1061), .A1(n454), .B0(n1011), .B1(n418), .Y(n459) );
  XNOR2XL U631 ( .A(n986), .B(n977), .Y(n913) );
  XNOR2XL U632 ( .A(n991), .B(n947), .Y(n915) );
  XNOR2XL U633 ( .A(n681), .B(n1185), .Y(n882) );
  XNOR2XL U634 ( .A(n991), .B(n981), .Y(n883) );
  XNOR2XL U635 ( .A(n991), .B(n1158), .Y(n852) );
  OAI22XL U636 ( .A0(n1027), .A1(n911), .B0(n879), .B1(n1123), .Y(n910) );
  XNOR2XL U637 ( .A(n1224), .B(n1014), .Y(n880) );
  XNOR2XL U638 ( .A(n1021), .B(n968), .Y(n939) );
  OAI22XL U639 ( .A0(n1027), .A1(n982), .B0(n943), .B1(n1123), .Y(n980) );
  XNOR2XL U640 ( .A(n1224), .B(n983), .Y(n984) );
  OAI22XL U641 ( .A0(n1040), .A1(n950), .B0(n1038), .B1(n915), .Y(n951) );
  OAI22X1 U642 ( .A0(n6), .A1(n948), .B0(n1035), .B1(n914), .Y(n952) );
  OAI22XL U643 ( .A0(n1040), .A1(n992), .B0(n1038), .B1(n950), .Y(n993) );
  ADDFX2 U644 ( .A(n1043), .B(n1042), .CI(n1041), .CO(n1052), .S(n1091) );
  OAI22XL U645 ( .A0(n1040), .A1(n1037), .B0(n1038), .B1(n992), .Y(n1041) );
  OAI22XL U646 ( .A0(n6), .A1(n1034), .B0(n1035), .B1(n989), .Y(n1042) );
  XNOR2XL U647 ( .A(n1224), .B(n704), .Y(n630) );
  OAI22XL U648 ( .A0(n1027), .A1(n586), .B0(n585), .B1(n1123), .Y(n591) );
  NOR2BXL U649 ( .AN(n1124), .B(n1030), .Y(n592) );
  OAI22XL U650 ( .A0(n1065), .A1(n588), .B0(n1063), .B1(n587), .Y(n590) );
  OAI22XL U651 ( .A0(n1027), .A1(n585), .B0(n629), .B1(n1123), .Y(n632) );
  NAND2BXL U652 ( .AN(n1124), .B(n1224), .Y(n581) );
  ADDFX2 U653 ( .A(n623), .B(n622), .CI(n621), .CO(n1110), .S(n609) );
  OAI22XL U654 ( .A0(n1040), .A1(n604), .B0(n1038), .B1(n625), .Y(n621) );
  OAI22XL U655 ( .A0(n6), .A1(n599), .B0(n1035), .B1(n598), .Y(n622) );
  OAI22XL U656 ( .A0(n1040), .A1(n1039), .B0(n1038), .B1(n1037), .Y(n1081) );
  OAI22XL U657 ( .A0(n6), .A1(n1036), .B0(n1035), .B1(n1034), .Y(n1082) );
  OAI22XL U658 ( .A0(n214), .A1(n411), .B0(n1072), .B1(n376), .Y(n387) );
  OAI22XL U659 ( .A0(n1061), .A1(n382), .B0(n1011), .B1(n374), .Y(n389) );
  OAI21XL U660 ( .A0(n1229), .A1(n121), .B0(n120), .Y(n388) );
  OAI22XL U661 ( .A0(n1162), .A1(n383), .B0(n1163), .B1(n377), .Y(n410) );
  OAI2BB1XL U662 ( .A0N(n1038), .A1N(n1040), .B0(n367), .Y(n384) );
  XNOR2XL U663 ( .A(n1224), .B(n968), .Y(n365) );
  ADDFX2 U664 ( .A(n373), .B(n372), .CI(n371), .CO(n354), .S(n405) );
  INVXL U665 ( .A(n351), .Y(n371) );
  OAI22XL U666 ( .A0(n214), .A1(n376), .B0(n1072), .B1(n343), .Y(n372) );
  OAI22XL U667 ( .A0(n1162), .A1(n377), .B0(n1163), .B1(n346), .Y(n368) );
  OAI22XL U668 ( .A0(n214), .A1(n343), .B0(n1072), .B1(n314), .Y(n349) );
  OAI22XL U669 ( .A0(n1205), .A1(n342), .B0(n1206), .B1(n316), .Y(n347) );
  INVXL U670 ( .A(n328), .Y(n317) );
  OAI22XL U671 ( .A0(n1229), .A1(n315), .B0(n1230), .B1(n311), .Y(n319) );
  OAI22XL U672 ( .A0(n1162), .A1(n341), .B0(n1163), .B1(n313), .Y(n318) );
  ADDFX2 U673 ( .A(n686), .B(n685), .CI(n684), .CO(n700), .S(n726) );
  OAI22XL U674 ( .A0(n214), .A1(n680), .B0(n1072), .B1(n645), .Y(n686) );
  OAI22XL U675 ( .A0(n89), .A1(n705), .B0(n1163), .B1(n646), .Y(n685) );
  XNOR2XL U676 ( .A(n991), .B(n945), .Y(n651) );
  XNOR2XL U677 ( .A(n991), .B(n1020), .Y(n636) );
  NAND2BXL U678 ( .AN(n1124), .B(n1214), .Y(n583) );
  ADDFX2 U679 ( .A(n603), .B(n602), .CI(n601), .CO(n610), .S(n669) );
  OAI22X1 U680 ( .A0(n6), .A1(n600), .B0(n1035), .B1(n599), .Y(n602) );
  ADDFX2 U681 ( .A(n644), .B(n643), .CI(n642), .CO(n659), .S(n688) );
  XNOR2XL U682 ( .A(n681), .B(n640), .Y(n184) );
  XNOR2XL U683 ( .A(n991), .B(n640), .Y(n165) );
  XNOR2XL U684 ( .A(n681), .B(n704), .Y(n183) );
  XNOR2XL U685 ( .A(n681), .B(n983), .Y(n153) );
  XNOR2XL U686 ( .A(n681), .B(n1028), .Y(n164) );
  NAND2BXL U687 ( .AN(n1124), .B(n991), .Y(n156) );
  ADDFX2 U688 ( .A(n160), .B(n159), .CI(n158), .CO(n233), .S(n161) );
  OAI22X1 U689 ( .A0(n1027), .A1(n154), .B0(n148), .B1(n1123), .Y(n159) );
  OAI22XL U690 ( .A0(n1040), .A1(n165), .B0(n1038), .B1(n152), .Y(n158) );
  NOR2BXL U691 ( .AN(n1124), .B(n1011), .Y(n160) );
  ADDFX2 U692 ( .A(n225), .B(n224), .CI(n223), .CO(n230), .S(n232) );
  OAI22XL U693 ( .A0(n652), .A1(n152), .B0(n1038), .B1(n210), .Y(n223) );
  OAI22X1 U694 ( .A0(n1061), .A1(n151), .B0(n1011), .B1(n219), .Y(n224) );
  OAI22XL U695 ( .A0(n6), .A1(n153), .B0(n1035), .B1(n208), .Y(n225) );
  ADDFX2 U696 ( .A(n228), .B(n227), .CI(n226), .CO(n255), .S(n229) );
  OAI22X1 U697 ( .A0(n1040), .A1(n210), .B0(n1038), .B1(n209), .Y(n227) );
  OAI22XL U698 ( .A0(n6), .A1(n208), .B0(n1035), .B1(n213), .Y(n228) );
  ADDFX2 U699 ( .A(n222), .B(n221), .CI(n220), .CO(n245), .S(n231) );
  OAI22XL U700 ( .A0(n1027), .A1(n217), .B0(n216), .B1(n1123), .Y(n221) );
  ADDFX2 U701 ( .A(n756), .B(n755), .CI(n754), .CO(n761), .S(n1125) );
  XNOR2XL U702 ( .A(n1224), .B(n1158), .Y(n1159) );
  OAI2BB1XL U703 ( .A0N(n819), .A1N(n6), .B0(n415), .Y(n475) );
  INVXL U704 ( .A(n414), .Y(n415) );
  CMPR32X1 U705 ( .A(n811), .B(n810), .C(n809), .CO(n494), .S(n831) );
  OAI22XL U706 ( .A0(n1061), .A1(n480), .B0(n1011), .B1(n454), .Y(n811) );
  NOR2XL U707 ( .A(n1030), .B(n807), .Y(n837) );
  OAI22XL U708 ( .A0(n1205), .A1(n835), .B0(n1206), .B1(n808), .Y(n836) );
  OAI22XL U709 ( .A0(n214), .A1(n824), .B0(n1072), .B1(n812), .Y(n841) );
  OAI22XL U710 ( .A0(n1040), .A1(n806), .B0(n1038), .B1(n474), .Y(n488) );
  OAI22XL U711 ( .A0(n214), .A1(n812), .B0(n1072), .B1(n478), .Y(n491) );
  OR2XL U712 ( .A(n816), .B(n815), .Y(n489) );
  OAI2BB1XL U713 ( .A0N(n827), .A1N(n1027), .B0(n486), .Y(n821) );
  OAI22XL U714 ( .A0(n6), .A1(n818), .B0(n819), .B1(n485), .Y(n822) );
  OAI22X1 U715 ( .A0(n1065), .A1(n871), .B0(n1063), .B1(n834), .Y(n874) );
  OAI22XL U716 ( .A0(n214), .A1(n876), .B0(n1072), .B1(n824), .Y(n857) );
  OAI22XL U717 ( .A0(n1040), .A1(n852), .B0(n1038), .B1(n820), .Y(n853) );
  ADDFX2 U718 ( .A(n938), .B(n937), .CI(n936), .CO(n923), .S(n957) );
  OAI22XL U719 ( .A0(n1061), .A1(n933), .B0(n1011), .B1(n902), .Y(n938) );
  OAI22X1 U720 ( .A0(n1065), .A1(n934), .B0(n1063), .B1(n903), .Y(n937) );
  OAI22XL U721 ( .A0(n1061), .A1(n969), .B0(n1011), .B1(n933), .Y(n976) );
  OAI22X1 U722 ( .A0(n1065), .A1(n971), .B0(n1063), .B1(n934), .Y(n975) );
  ADDFX2 U723 ( .A(n1052), .B(n1051), .CI(n1050), .CO(n1055), .S(n1093) );
  OAI22X1 U724 ( .A0(n214), .A1(n624), .B0(n1072), .B1(n1073), .Y(n1101) );
  ADDFX2 U725 ( .A(n611), .B(n610), .CI(n609), .CO(n1143), .S(n658) );
  NOR2XL U726 ( .A(n1030), .B(n579), .Y(n616) );
  OAI22XL U727 ( .A0(n1205), .A1(n595), .B0(n1067), .B1(n626), .Y(n615) );
  OAI22XL U728 ( .A0(n6), .A1(n598), .B0(n1035), .B1(n1036), .Y(n1078) );
  INVXL U729 ( .A(n1182), .Y(n1166) );
  OAI22XL U730 ( .A0(n1229), .A1(n323), .B0(n1230), .B1(n1165), .Y(n1168) );
  OAI22XL U731 ( .A0(n1205), .A1(n326), .B0(n1206), .B1(n1164), .Y(n1171) );
  OAI22XL U732 ( .A0(n1205), .A1(n316), .B0(n1206), .B1(n312), .Y(n322) );
  XNOR2XL U733 ( .A(n1224), .B(n988), .Y(n300) );
  ADDFX2 U734 ( .A(n392), .B(n391), .CI(n390), .CO(n394), .S(n431) );
  CMPR32X1 U735 ( .A(n358), .B(n357), .C(n356), .CO(n359), .S(n393) );
  OAI22XL U736 ( .A0(n6), .A1(n413), .B0(n819), .B1(n178), .Y(n179) );
  NAND2BXL U737 ( .AN(n1124), .B(n681), .Y(n178) );
  OR2XL U738 ( .A(n1303), .B(n1309), .Y(n1313) );
  INVXL U739 ( .A(n1311), .Y(n1312) );
  NAND2XL U740 ( .A(n1282), .B(n1326), .Y(n1283) );
  OAI22XL U741 ( .A0(n1229), .A1(n1197), .B0(n1230), .B1(n1215), .Y(n1211) );
  CMPR32X1 U742 ( .A(n1180), .B(n1179), .C(n1178), .CO(n1193), .S(n1176) );
  INVXL U743 ( .A(mult_x_1_n306), .Y(n770) );
  ADDFX2 U744 ( .A(n850), .B(n849), .CI(n848), .CO(n844), .S(n869) );
  CMPR32X1 U745 ( .A(n958), .B(n957), .C(n956), .CO(n967), .S(n1005) );
  NAND2BXL U746 ( .AN(n1070), .B(n139), .Y(n138) );
  CMPR32X1 U747 ( .A(n1089), .B(n1088), .C(n1087), .CO(n1098), .S(n1118) );
  XOR2X1 U748 ( .A(n1069), .B(n140), .Y(n1088) );
  ADDFX2 U749 ( .A(n1113), .B(n1112), .CI(n1111), .CO(n1122), .S(n1145) );
  ADDFX2 U750 ( .A(n1157), .B(n1156), .CI(n1155), .CO(n1177), .S(n336) );
  OAI2BB1X1 U751 ( .A0N(n722), .A1N(n721), .B0(n133), .Y(n696) );
  OAI21XL U752 ( .A0(n721), .A1(n722), .B0(n720), .Y(n133) );
  NAND2XL U753 ( .A(n796), .B(n795), .Y(n797) );
  NAND2XL U754 ( .A(n397), .B(n396), .Y(mult_x_1_n170) );
  NOR2XL U755 ( .A(n1177), .B(n1176), .Y(mult_x_1_n136) );
  NAND2XL U756 ( .A(n1237), .B(n1236), .Y(mult_x_1_n58) );
  NAND2XL U757 ( .A(n1235), .B(n1234), .Y(n1236) );
  NOR2XL U758 ( .A(n1220), .B(n1219), .Y(mult_x_1_n109) );
  NAND2XL U759 ( .A(n1220), .B(n1219), .Y(mult_x_1_n110) );
  NOR2XL U760 ( .A(n1208), .B(n1207), .Y(mult_x_1_n120) );
  NAND2XL U761 ( .A(n1208), .B(n1207), .Y(mult_x_1_n121) );
  NOR2XL U762 ( .A(n1193), .B(n1192), .Y(mult_x_1_n129) );
  NAND2XL U763 ( .A(n1193), .B(n1192), .Y(mult_x_1_n130) );
  NAND2XL U764 ( .A(n1177), .B(n1176), .Y(mult_x_1_n137) );
  NAND2X1 U765 ( .A(n142), .B(n141), .Y(n900) );
  NAND2XL U766 ( .A(n928), .B(n929), .Y(n141) );
  NAND2XL U767 ( .A(n136), .B(n135), .Y(mult_x_1_n617) );
  NAND2XL U768 ( .A(n1097), .B(n1098), .Y(n135) );
  NOR2BXL U769 ( .AN(n1124), .B(n1123), .Y(n1404) );
  NAND2XL U770 ( .A(n1291), .B(n1290), .Y(n1293) );
  XOR2XL U771 ( .A(n1289), .B(n1288), .Y(n1401) );
  NAND2XL U772 ( .A(n1287), .B(n1286), .Y(n1289) );
  INVXL U773 ( .A(n1285), .Y(n1287) );
  NAND2XL U774 ( .A(n187), .B(n1298), .Y(n1300) );
  NAND2XL U775 ( .A(n1318), .B(n1317), .Y(n1320) );
  INVXL U776 ( .A(n1316), .Y(n1318) );
  NAND2XL U777 ( .A(n1265), .B(n1264), .Y(n1267) );
  INVXL U778 ( .A(n1263), .Y(n1265) );
  NAND2XL U779 ( .A(n1260), .B(n1259), .Y(n1261) );
  INVX8 U780 ( .A(n307), .Y(n1021) );
  NAND2X1 U781 ( .A(n551), .B(n289), .Y(n508) );
  INVX4 U782 ( .A(B[9]), .Y(n307) );
  ADDFX2 U783 ( .A(n1127), .B(n1126), .CI(n1125), .CO(n763), .S(n1132) );
  XOR2X1 U784 ( .A(n143), .B(n118), .Y(PRODUCT[33]) );
  CMPR22X1 U785 ( .A(n878), .B(n877), .CO(n855), .S(n888) );
  CMPR22X1 U786 ( .A(n942), .B(n941), .CO(n918), .S(n954) );
  CMPR22X1 U787 ( .A(n1024), .B(n1023), .CO(n995), .S(n1045) );
  CMPR22X1 U788 ( .A(n186), .B(n185), .CO(n188), .S(n180) );
  OAI22X1 U789 ( .A0(n6), .A1(n176), .B0(n1035), .B1(n184), .Y(n185) );
  CMPR22X1 U790 ( .A(n826), .B(n825), .CO(n840), .S(n856) );
  CMPR22X1 U791 ( .A(n168), .B(n167), .CO(n162), .S(n191) );
  OAI22X1 U792 ( .A0(n1061), .A1(n902), .B0(n1011), .B1(n870), .Y(n907) );
  CMPR22X1 U793 ( .A(n212), .B(n211), .CO(n226), .S(n234) );
  OAI22X1 U794 ( .A0(n1061), .A1(n302), .B0(n1011), .B1(n146), .Y(n211) );
  OAI22X1 U795 ( .A0(n214), .A1(n314), .B0(n1072), .B1(n309), .Y(n328) );
  NAND2X1 U796 ( .A(n561), .B(n560), .Y(n562) );
  XNOR2X1 U797 ( .A(n1214), .B(n990), .Y(n121) );
  ADDFX2 U798 ( .A(n268), .B(n267), .CI(n266), .CO(n780), .S(n264) );
  OAI21XL U799 ( .A0(n1314), .A1(n1303), .B0(n1310), .Y(n143) );
  NOR2X1 U800 ( .A(n1303), .B(n1337), .Y(n338) );
  OAI22X1 U801 ( .A0(n417), .A1(n1229), .B0(n1230), .B1(n121), .Y(n426) );
  AOI21X4 U802 ( .A0(n126), .A1(n509), .B0(n125), .Y(n1314) );
  OAI21X2 U803 ( .A0(n293), .A1(n538), .B0(n292), .Y(n125) );
  NOR2X1 U804 ( .A(n1365), .B(n1366), .Y(n525) );
  NAND3BX4 U805 ( .AN(n130), .B(n128), .C(n1352), .Y(n664) );
  NAND3BX4 U806 ( .AN(n1351), .B(n129), .C(n1359), .Y(n128) );
  NOR2X1 U807 ( .A(n1351), .B(n1358), .Y(n130) );
  XOR2X1 U808 ( .A(n134), .B(n720), .Y(n757) );
  XOR2X1 U809 ( .A(n721), .B(n722), .Y(n134) );
  XOR2X1 U810 ( .A(B[14]), .B(B[15]), .Y(n305) );
  XNOR2X2 U811 ( .A(B[7]), .B(B[8]), .Y(n206) );
  OAI22X1 U812 ( .A0(n1229), .A1(n584), .B0(n1230), .B1(n583), .Y(n637) );
  OAI22X2 U813 ( .A0(n1065), .A1(n903), .B0(n1063), .B1(n871), .Y(n906) );
  BUFX12 U814 ( .A(B[13]), .Y(n1187) );
  OAI21X1 U815 ( .A0(n793), .A1(n241), .B0(n240), .Y(n775) );
  NAND2X1 U816 ( .A(n1374), .B(n1373), .Y(n555) );
  NOR2X1 U817 ( .A(n1372), .B(n1371), .Y(n548) );
  ADDFX2 U818 ( .A(n1000), .B(n999), .CI(n998), .CO(n1009), .S(n1054) );
  OAI22X1 U819 ( .A0(n1229), .A1(n458), .B0(n1230), .B1(n417), .Y(n460) );
  NAND2X2 U820 ( .A(n305), .B(n457), .Y(n456) );
  OAI21XL U821 ( .A0(n568), .A1(n508), .B0(n538), .Y(n543) );
  OAI22X1 U822 ( .A0(n1065), .A1(n582), .B0(n1063), .B1(n1064), .Y(n1079) );
  CMPR22X1 U823 ( .A(n1077), .B(n1076), .CO(n1084), .S(n1106) );
  XNOR2X1 U824 ( .A(n1214), .B(n985), .Y(n903) );
  XNOR2X1 U825 ( .A(n1187), .B(n981), .Y(n342) );
  XNOR2X1 U826 ( .A(n1187), .B(n990), .Y(n473) );
  XNOR2X1 U827 ( .A(n1187), .B(n983), .Y(n595) );
  XNOR2X1 U828 ( .A(n1187), .B(n704), .Y(n641) );
  XNOR2X1 U829 ( .A(n1187), .B(n977), .Y(n872) );
  XNOR2X1 U830 ( .A(n1187), .B(n988), .Y(n379) );
  XNOR2X1 U831 ( .A(n1187), .B(n972), .Y(n1015) );
  OAI21XL U832 ( .A0(n1314), .A1(n503), .B0(n504), .Y(n472) );
  ADDHXL U833 ( .A(n710), .B(n709), .CO(n706), .S(n746) );
  XNOR2X1 U834 ( .A(n1021), .B(n704), .Y(n260) );
  XNOR2XL U835 ( .A(B[1]), .B(n1185), .Y(n943) );
  NOR2X1 U836 ( .A(n772), .B(n788), .Y(n774) );
  XNOR2XL U837 ( .A(n1293), .B(n1292), .Y(n1402) );
  INVX1 U838 ( .A(B[0]), .Y(n827) );
  XNOR2X1 U839 ( .A(B[1]), .B(n970), .Y(n148) );
  XNOR2X1 U840 ( .A(B[1]), .B(n1014), .Y(n217) );
  BUFX3 U841 ( .A(n827), .Y(n1123) );
  OAI22X1 U842 ( .A0(n1027), .A1(n148), .B0(n217), .B1(n1123), .Y(n212) );
  XOR2X1 U843 ( .A(B[6]), .B(B[7]), .Y(n145) );
  NAND2X2 U844 ( .A(n145), .B(n147), .Y(n628) );
  BUFX3 U845 ( .A(n147), .Y(n1011) );
  BUFX3 U846 ( .A(A[0]), .Y(n1124) );
  XNOR2X1 U847 ( .A(B[1]), .B(n1012), .Y(n154) );
  XOR2X1 U848 ( .A(B[4]), .B(B[5]), .Y(n149) );
  XOR2X1 U849 ( .A(B[2]), .B(B[3]), .Y(n150) );
  NAND2X1 U850 ( .A(n150), .B(n819), .Y(n177) );
  XNOR2X1 U851 ( .A(B[1]), .B(n983), .Y(n181) );
  OAI22X1 U852 ( .A0(n1027), .A1(n181), .B0(n154), .B1(n1123), .Y(n168) );
  OAI22X1 U853 ( .A0(n1040), .A1(n157), .B0(n1038), .B1(n156), .Y(n167) );
  CMPR32X1 U854 ( .A(n163), .B(n162), .C(n161), .CO(n201), .S(n200) );
  OAI22XL U855 ( .A0(n1040), .A1(n166), .B0(n1038), .B1(n165), .Y(n192) );
  NOR2XL U856 ( .A(n1258), .B(n1263), .Y(n204) );
  XNOR2X1 U857 ( .A(B[1]), .B(n704), .Y(n175) );
  BUFX3 U858 ( .A(n170), .Y(n1027) );
  XNOR2X1 U859 ( .A(B[1]), .B(n1028), .Y(n182) );
  OAI22X1 U860 ( .A0(n1027), .A1(n175), .B0(n182), .B1(n1123), .Y(n186) );
  XNOR2X1 U861 ( .A(n681), .B(n1124), .Y(n176) );
  OAI21XL U862 ( .A0(n1288), .A1(n1285), .B0(n1286), .Y(n1299) );
  NAND2XL U863 ( .A(n189), .B(n188), .Y(n1298) );
  INVXL U864 ( .A(n1298), .Y(n190) );
  AOI21XL U865 ( .A0(n1299), .A1(n187), .B0(n190), .Y(n1319) );
  CMPR32X1 U866 ( .A(n193), .B(n192), .C(n191), .CO(n199), .S(n198) );
  CMPR32X1 U867 ( .A(n196), .B(n195), .C(n194), .CO(n197), .S(n189) );
  NOR2XL U868 ( .A(n198), .B(n197), .Y(n1316) );
  OAI21XL U869 ( .A0(n1319), .A1(n1316), .B0(n1317), .Y(n1257) );
  NAND2XL U870 ( .A(n202), .B(n201), .Y(n1259) );
  OAI21XL U871 ( .A0(n1258), .A1(n1264), .B0(n1259), .Y(n203) );
  AOI21XL U872 ( .A0(n204), .A1(n1257), .B0(n203), .Y(n793) );
  XNOR2XL U873 ( .A(n1021), .B(n1124), .Y(n207) );
  BUFX8 U874 ( .A(n206), .Y(n1072) );
  XNOR2X1 U875 ( .A(n681), .B(n1014), .Y(n244) );
  XNOR2X1 U876 ( .A(B[1]), .B(n972), .Y(n216) );
  XNOR2X1 U877 ( .A(B[1]), .B(n985), .Y(n250) );
  OAI22X1 U878 ( .A0(n1027), .A1(n216), .B0(n250), .B1(n1123), .Y(n249) );
  OAI22XL U879 ( .A0(n628), .A1(n219), .B0(n1011), .B1(n218), .Y(n220) );
  CMPR32X1 U880 ( .A(n234), .B(n233), .C(n232), .CO(n235), .S(n202) );
  OR2X2 U881 ( .A(n236), .B(n235), .Y(n800) );
  NAND2XL U882 ( .A(n236), .B(n235), .Y(n799) );
  INVXL U883 ( .A(n799), .Y(n794) );
  INVXL U884 ( .A(n795), .Y(n239) );
  INVX1 U885 ( .A(n775), .Y(n792) );
  XNOR2X1 U886 ( .A(n991), .B(n970), .Y(n259) );
  XNOR2X1 U887 ( .A(n681), .B(n972), .Y(n274) );
  CMPR22X1 U888 ( .A(n249), .B(n248), .CO(n265), .S(n246) );
  NOR2BX1 U889 ( .AN(n1124), .B(n1031), .Y(n268) );
  XNOR2X1 U890 ( .A(B[1]), .B(n945), .Y(n261) );
  OAI22XL U891 ( .A0(n170), .A1(n250), .B0(n261), .B1(n1123), .Y(n267) );
  OAI21XL U892 ( .A0(n792), .A1(n788), .B0(n789), .Y(n282) );
  XNOR2X1 U893 ( .A(B[1]), .B(n1020), .Y(n712) );
  BUFX3 U894 ( .A(n1031), .Y(n1163) );
  INVX8 U895 ( .A(n306), .Y(n986) );
  CMPR32X1 U896 ( .A(n271), .B(n270), .C(n269), .CO(n779), .S(n277) );
  OAI22X1 U897 ( .A0(n1061), .A1(n272), .B0(n1011), .B1(n716), .Y(n748) );
  XNOR2X1 U898 ( .A(n986), .B(n640), .Y(n714) );
  OAI22X1 U899 ( .A0(n6), .A1(n274), .B0(n1035), .B1(n718), .Y(n747) );
  CMPR32X1 U900 ( .A(n277), .B(n276), .C(n275), .CO(n278), .S(n258) );
  INVXL U901 ( .A(n772), .Y(n280) );
  NAND2XL U902 ( .A(n280), .B(n771), .Y(n281) );
  XNOR2X1 U903 ( .A(n282), .B(n281), .Y(n1393) );
  INVXL U904 ( .A(n1347), .Y(n284) );
  NAND2XL U905 ( .A(n284), .B(n1348), .Y(n285) );
  XOR2X1 U906 ( .A(n286), .B(n285), .Y(PRODUCT[18]) );
  NOR2X1 U907 ( .A(n1373), .B(n1374), .Y(n544) );
  NOR2X1 U908 ( .A(n544), .B(n548), .Y(n289) );
  NOR2X1 U909 ( .A(n1369), .B(n1370), .Y(n539) );
  NOR2X2 U910 ( .A(n1367), .B(n1368), .Y(n533) );
  NOR2X1 U911 ( .A(n1363), .B(n1364), .Y(n515) );
  NOR2X1 U912 ( .A(n525), .B(n515), .Y(n291) );
  NAND2X1 U913 ( .A(n1371), .B(n1372), .Y(n549) );
  AOI21X2 U914 ( .A0(n289), .A1(n552), .B0(n288), .Y(n538) );
  NAND2X1 U915 ( .A(n1369), .B(n1370), .Y(n540) );
  NAND2X1 U916 ( .A(n1367), .B(n1368), .Y(n534) );
  OAI21X1 U917 ( .A0(n533), .A1(n540), .B0(n534), .Y(n510) );
  NAND2X1 U918 ( .A(n1365), .B(n1366), .Y(n526) );
  NAND2X1 U919 ( .A(n1363), .B(n1364), .Y(n516) );
  OAI21XL U920 ( .A0(n515), .A1(n526), .B0(n516), .Y(n290) );
  NOR2XL U921 ( .A(n503), .B(n1343), .Y(n398) );
  NAND2XL U922 ( .A(n398), .B(n294), .Y(n1303) );
  NAND2XL U923 ( .A(n338), .B(n1238), .Y(n296) );
  AOI21XL U924 ( .A0(n339), .A1(n1238), .B0(n1241), .Y(n295) );
  XNOR2X1 U925 ( .A(n298), .B(n297), .Y(PRODUCT[35]) );
  XNOR2X2 U926 ( .A(B[12]), .B(B[11]), .Y(n580) );
  NAND2X2 U927 ( .A(n299), .B(n580), .Y(n1016) );
  BUFX8 U928 ( .A(n1016), .Y(n1205) );
  XNOR2X1 U929 ( .A(n1187), .B(n1158), .Y(n316) );
  BUFX1 U930 ( .A(A[21]), .Y(n1185) );
  XNOR2X1 U931 ( .A(n1187), .B(n1185), .Y(n312) );
  OAI22X1 U932 ( .A0(n1061), .A1(n374), .B0(n1011), .B1(n303), .Y(n351) );
  OAI2BB1X1 U933 ( .A0N(n1011), .A1N(n1061), .B0(n304), .Y(n350) );
  XNOR2X2 U934 ( .A(B[14]), .B(B[13]), .Y(n457) );
  BUFX4 U935 ( .A(n456), .Y(n1229) );
  BUFX3 U936 ( .A(n457), .Y(n1230) );
  XNOR2X1 U937 ( .A(n986), .B(n1201), .Y(n341) );
  XNOR2X1 U938 ( .A(n986), .B(n1212), .Y(n313) );
  XNOR2XL U939 ( .A(B[9]), .B(A[24]), .Y(n314) );
  XNOR2X1 U940 ( .A(n1187), .B(n1201), .Y(n326) );
  XNOR2X1 U941 ( .A(n986), .B(A[24]), .Y(n325) );
  XNOR2XL U942 ( .A(n1021), .B(n1212), .Y(n343) );
  OAI22XL U943 ( .A0(n1229), .A1(n345), .B0(n1230), .B1(n315), .Y(n348) );
  CMPR32X1 U944 ( .A(n319), .B(n318), .C(n317), .CO(n335), .S(n357) );
  CMPR32X1 U945 ( .A(n322), .B(n321), .C(n320), .CO(n361), .S(n356) );
  XNOR2X1 U946 ( .A(n986), .B(A[25]), .Y(n1160) );
  OAI22X1 U947 ( .A0(n1162), .A1(n325), .B0(n1163), .B1(n1160), .Y(n1182) );
  XNOR2X1 U948 ( .A(n1187), .B(n1212), .Y(n1164) );
  CMPR32X1 U949 ( .A(n329), .B(n328), .C(n327), .CO(n1170), .S(n334) );
  CMPR32X1 U950 ( .A(n332), .B(n331), .C(n330), .CO(n1169), .S(n333) );
  CMPR32X1 U951 ( .A(n335), .B(n334), .C(n333), .CO(n1155), .S(n360) );
  NOR2XL U952 ( .A(n337), .B(n336), .Y(mult_x_1_n151) );
  NAND2XL U953 ( .A(n337), .B(n336), .Y(mult_x_1_n152) );
  XNOR2X1 U954 ( .A(n986), .B(n1185), .Y(n346) );
  XNOR2X1 U955 ( .A(n1187), .B(n947), .Y(n378) );
  XNOR2X1 U956 ( .A(n1224), .B(n990), .Y(n344) );
  OAI22XL U957 ( .A0(n1229), .A1(n375), .B0(n1230), .B1(n345), .Y(n369) );
  XNOR2X1 U958 ( .A(n986), .B(n1158), .Y(n377) );
  CMPR32X1 U959 ( .A(n349), .B(n348), .C(n347), .CO(n358), .S(n392) );
  CMPR32X1 U960 ( .A(n352), .B(n351), .C(n350), .CO(n320), .S(n391) );
  NOR2XL U961 ( .A(n363), .B(n362), .Y(mult_x_1_n160) );
  NAND2XL U962 ( .A(n363), .B(n362), .Y(mult_x_1_n161) );
  OAI22X1 U963 ( .A0(n1040), .A1(n416), .B0(n1038), .B1(n366), .Y(n385) );
  CMPR32X1 U964 ( .A(n370), .B(n369), .C(n368), .CO(n353), .S(n406) );
  XNOR2X1 U965 ( .A(B[9]), .B(n1185), .Y(n411) );
  XNOR2XL U966 ( .A(n986), .B(n981), .Y(n383) );
  OAI22XL U967 ( .A0(n1205), .A1(n379), .B0(n1206), .B1(n378), .Y(n409) );
  XNOR2XL U968 ( .A(n1224), .B(A[13]), .Y(n381) );
  INVXL U969 ( .A(n385), .Y(n422) );
  XNOR2X1 U970 ( .A(n1214), .B(n968), .Y(n417) );
  XNOR2XL U971 ( .A(n986), .B(n947), .Y(n421) );
  OAI22XL U972 ( .A0(n1162), .A1(n421), .B0(n1163), .B1(n383), .Y(n425) );
  CMPR32X1 U973 ( .A(n386), .B(n385), .C(n384), .CO(n407), .S(n446) );
  CMPR32X1 U974 ( .A(n389), .B(n388), .C(n387), .CO(n430), .S(n445) );
  CMPR32X1 U975 ( .A(n395), .B(n394), .C(n393), .CO(n363), .S(n396) );
  NOR2XL U976 ( .A(n397), .B(n396), .Y(mult_x_1_n169) );
  AOI21XL U977 ( .A0(n436), .A1(n439), .B0(n399), .Y(n400) );
  CMPR32X1 U978 ( .A(n407), .B(n406), .C(n405), .CO(n433), .S(n444) );
  CMPR32X1 U979 ( .A(n410), .B(n409), .C(n408), .CO(n429), .S(n450) );
  XNOR2XL U980 ( .A(n1224), .B(n977), .Y(n412) );
  NOR2XL U981 ( .A(n1030), .B(n412), .Y(n477) );
  XNOR2X1 U982 ( .A(n681), .B(A[24]), .Y(n485) );
  XNOR2X1 U983 ( .A(n681), .B(A[25]), .Y(n414) );
  XNOR2X1 U984 ( .A(n991), .B(n1212), .Y(n474) );
  OAI22XL U985 ( .A0(n1040), .A1(n474), .B0(n1038), .B1(n416), .Y(n461) );
  XNOR2X1 U986 ( .A(n1214), .B(A[13]), .Y(n458) );
  XNOR2X1 U987 ( .A(n1021), .B(n981), .Y(n478) );
  OAI22X1 U988 ( .A0(n214), .A1(n478), .B0(n1072), .B1(n419), .Y(n464) );
  OAI22X1 U989 ( .A0(n1205), .A1(n473), .B0(n1206), .B1(n420), .Y(n463) );
  XNOR2X1 U990 ( .A(n986), .B(n988), .Y(n479) );
  OAI22XL U991 ( .A0(n1162), .A1(n479), .B0(n1163), .B1(n421), .Y(n462) );
  CMPR32X1 U992 ( .A(n433), .B(n432), .C(n431), .CO(n397), .S(n434) );
  NOR2XL U993 ( .A(n435), .B(n434), .Y(mult_x_1_n176) );
  NAND2XL U994 ( .A(n435), .B(n434), .Y(mult_x_1_n177) );
  ADDFHX1 U995 ( .A(n444), .B(n443), .CI(n442), .CO(n435), .S(n469) );
  CMPR32X1 U996 ( .A(n447), .B(n446), .C(n445), .CO(n428), .S(n500) );
  ADDFHX1 U997 ( .A(n450), .B(n449), .CI(n448), .CO(n443), .S(n499) );
  CMPR32X1 U998 ( .A(n453), .B(n452), .C(n451), .CO(n449), .S(n484) );
  XNOR2XL U999 ( .A(n1224), .B(n1020), .Y(n455) );
  NOR2XL U1000 ( .A(n1030), .B(n455), .Y(n810) );
  XNOR2X1 U1001 ( .A(n1214), .B(n977), .Y(n481) );
  OAI22XL U1002 ( .A0(n1065), .A1(n481), .B0(n1063), .B1(n458), .Y(n809) );
  CMPR32X1 U1003 ( .A(n461), .B(n460), .C(n459), .CO(n451), .S(n493) );
  CMPR32X1 U1004 ( .A(n467), .B(n466), .C(n465), .CO(n448), .S(n482) );
  NOR2XL U1005 ( .A(n469), .B(n468), .Y(mult_x_1_n183) );
  NAND2XL U1006 ( .A(n469), .B(n468), .Y(mult_x_1_n184) );
  XNOR2X1 U1007 ( .A(n1187), .B(n968), .Y(n808) );
  XNOR2X1 U1008 ( .A(n991), .B(n1201), .Y(n806) );
  OAI22XL U1009 ( .A0(n1065), .A1(n834), .B0(n1063), .B1(n481), .Y(n815) );
  XNOR2X1 U1010 ( .A(B[3]), .B(n1212), .Y(n818) );
  XNOR2X1 U1011 ( .A(B[1]), .B(A[25]), .Y(n813) );
  CMPR32X1 U1012 ( .A(n491), .B(n490), .C(n489), .CO(n495), .S(n848) );
  CMPR32X1 U1013 ( .A(n497), .B(n496), .C(n495), .CO(n805), .S(n842) );
  ADDFHX1 U1014 ( .A(n500), .B(n499), .CI(n498), .CO(n468), .S(n501) );
  NOR2XL U1015 ( .A(n502), .B(n501), .Y(mult_x_1_n194) );
  NAND2XL U1016 ( .A(n502), .B(n501), .Y(mult_x_1_n195) );
  NAND2XL U1017 ( .A(n512), .B(n537), .Y(n514) );
  INVX1 U1018 ( .A(n538), .Y(n531) );
  OAI21XL U1019 ( .A0(n514), .A1(n568), .B0(n513), .Y(n519) );
  XNOR2X1 U1020 ( .A(n519), .B(n518), .Y(PRODUCT[28]) );
  INVXL U1021 ( .A(n520), .Y(n522) );
  OAI21XL U1022 ( .A0(n568), .A1(n524), .B0(n523), .Y(n529) );
  INVXL U1023 ( .A(n525), .Y(n527) );
  NAND2X1 U1024 ( .A(n527), .B(n526), .Y(n528) );
  INVXL U1025 ( .A(n540), .Y(n530) );
  NAND2XL U1026 ( .A(n551), .B(n556), .Y(n547) );
  INVXL U1027 ( .A(n555), .Y(n545) );
  INVXL U1028 ( .A(n548), .Y(n550) );
  INVXL U1029 ( .A(n551), .Y(n554) );
  INVXL U1030 ( .A(n552), .Y(n553) );
  NAND2XL U1031 ( .A(n556), .B(n555), .Y(n557) );
  XNOR2X1 U1032 ( .A(n558), .B(n557), .Y(PRODUCT[23]) );
  OAI21X1 U1033 ( .A0(n568), .A1(n564), .B0(n565), .Y(n563) );
  INVXL U1034 ( .A(n559), .Y(n561) );
  XNOR2X1 U1035 ( .A(n563), .B(n562), .Y(PRODUCT[22]) );
  INVXL U1036 ( .A(n564), .Y(n566) );
  AOI21X1 U1037 ( .A0(n664), .A1(n570), .B0(n569), .Y(n578) );
  INVXL U1038 ( .A(n571), .Y(n573) );
  INVXL U1039 ( .A(n1345), .Y(n576) );
  NAND2XL U1040 ( .A(n576), .B(n1346), .Y(n577) );
  XNOR2X1 U1041 ( .A(n1214), .B(n704), .Y(n587) );
  XNOR2X1 U1042 ( .A(n1214), .B(n1028), .Y(n582) );
  OAI22XL U1043 ( .A0(n1065), .A1(n587), .B0(n1063), .B1(n582), .Y(n617) );
  XNOR2X1 U1044 ( .A(n1224), .B(n640), .Y(n579) );
  XNOR2X1 U1045 ( .A(n1187), .B(n1012), .Y(n626) );
  OAI22XL U1046 ( .A0(n628), .A1(n607), .B0(n147), .B1(n627), .Y(n620) );
  OAI22XL U1047 ( .A0(n214), .A1(n593), .B0(n1072), .B1(n624), .Y(n619) );
  XNOR2X1 U1048 ( .A(B[1]), .B(n949), .Y(n585) );
  XNOR2X1 U1049 ( .A(B[1]), .B(n988), .Y(n629) );
  XNOR2X1 U1050 ( .A(n986), .B(n1014), .Y(n597) );
  XNOR2X1 U1051 ( .A(n1214), .B(n983), .Y(n1064) );
  XNOR2X1 U1052 ( .A(B[3]), .B(n990), .Y(n598) );
  XNOR2X1 U1053 ( .A(n681), .B(n949), .Y(n1036) );
  XNOR2X1 U1054 ( .A(B[1]), .B(n968), .Y(n639) );
  XNOR2X1 U1055 ( .A(B[1]), .B(n990), .Y(n586) );
  OAI22X1 U1056 ( .A0(n1027), .A1(n639), .B0(n586), .B1(n1123), .Y(n638) );
  XNOR2X1 U1057 ( .A(n1214), .B(n640), .Y(n588) );
  XNOR2X1 U1058 ( .A(n1187), .B(n1028), .Y(n596) );
  CMPR32X1 U1059 ( .A(n592), .B(n591), .C(n590), .CO(n611), .S(n643) );
  XNOR2X1 U1060 ( .A(n681), .B(A[13]), .Y(n600) );
  OAI22XL U1061 ( .A0(n1205), .A1(n596), .B0(n1067), .B1(n595), .Y(n601) );
  XNOR2X1 U1062 ( .A(n991), .B(n977), .Y(n604) );
  XNOR2X1 U1063 ( .A(n991), .B(A[13]), .Y(n625) );
  XNOR2X1 U1064 ( .A(n681), .B(n977), .Y(n647) );
  XNOR2X1 U1065 ( .A(n986), .B(n983), .Y(n646) );
  XNOR2X1 U1066 ( .A(n986), .B(n1012), .Y(n606) );
  OAI22X1 U1067 ( .A0(n1040), .A1(n636), .B0(n1038), .B1(n604), .Y(n614) );
  OAI22XL U1068 ( .A0(n628), .A1(n608), .B0(n147), .B1(n607), .Y(n612) );
  CMPR32X1 U1069 ( .A(n614), .B(n613), .C(n612), .CO(n635), .S(n668) );
  CMPR32X1 U1070 ( .A(n617), .B(n616), .C(n615), .CO(n1141), .S(n634) );
  CMPR32X1 U1071 ( .A(n620), .B(n619), .C(n618), .CO(n1140), .S(n633) );
  XNOR2X1 U1072 ( .A(n991), .B(n968), .Y(n1039) );
  XNOR2X1 U1073 ( .A(n1187), .B(n970), .Y(n1068) );
  OAI22XL U1074 ( .A0(n628), .A1(n627), .B0(n1011), .B1(n1060), .Y(n1107) );
  XNOR2X1 U1075 ( .A(B[1]), .B(n947), .Y(n1026) );
  OAI22X1 U1076 ( .A0(n1027), .A1(n629), .B0(n1026), .B1(n1123), .Y(n1077) );
  ADDHXL U1077 ( .A(n632), .B(n631), .CO(n1105), .S(n618) );
  CMPR22X1 U1078 ( .A(n638), .B(n637), .CO(n644), .S(n675) );
  XNOR2X1 U1079 ( .A(B[1]), .B(A[13]), .Y(n654) );
  XNOR2X1 U1080 ( .A(n986), .B(n1028), .Y(n705) );
  XNOR2X1 U1081 ( .A(n681), .B(n1020), .Y(n682) );
  OAI22XL U1082 ( .A0(n6), .A1(n682), .B0(n1035), .B1(n647), .Y(n684) );
  NOR2XL U1083 ( .A(n661), .B(n660), .Y(mult_x_1_n281) );
  CMPR32X1 U1084 ( .A(n670), .B(n669), .C(n668), .CO(n657), .S(n697) );
  CMPR32X1 U1085 ( .A(n673), .B(n672), .C(n671), .CO(n670), .S(n722) );
  CMPR32X1 U1086 ( .A(n676), .B(n675), .C(n674), .CO(n689), .S(n721) );
  XNOR2X1 U1087 ( .A(n1021), .B(n983), .Y(n735) );
  OAI22XL U1088 ( .A0(n6), .A1(n717), .B0(n1035), .B1(n682), .Y(n733) );
  OAI21XL U1089 ( .A0(n769), .A1(n1353), .B0(n1358), .Y(n694) );
  INVXL U1090 ( .A(n1351), .Y(n692) );
  NAND2XL U1091 ( .A(n692), .B(n1352), .Y(n693) );
  CMPR32X1 U1092 ( .A(n697), .B(n696), .C(n695), .CO(n690), .S(n724) );
  ADDFHX1 U1093 ( .A(n700), .B(n699), .CI(n698), .CO(n687), .S(n759) );
  XNOR2X1 U1094 ( .A(n1187), .B(n1124), .Y(n703) );
  XNOR2X1 U1095 ( .A(n986), .B(n704), .Y(n713) );
  CMPR32X1 U1096 ( .A(n708), .B(n707), .C(n706), .CO(n698), .S(n742) );
  NOR2XL U1097 ( .A(n724), .B(n723), .Y(mult_x_1_n292) );
  NAND2XL U1098 ( .A(n724), .B(n723), .Y(mult_x_1_n293) );
  OAI21XL U1099 ( .A0(n769), .A1(n1321), .B0(n1322), .Y(n725) );
  XNOR2X1 U1100 ( .A(n725), .B(n1354), .Y(PRODUCT[15]) );
  CMPR32X1 U1101 ( .A(n731), .B(n730), .C(n729), .CO(n743), .S(n756) );
  CMPR32X1 U1102 ( .A(n734), .B(n733), .C(n732), .CO(n727), .S(n755) );
  OAI22XL U1103 ( .A0(n214), .A1(n736), .B0(n1072), .B1(n735), .Y(n777) );
  CMPR32X1 U1104 ( .A(n740), .B(n739), .C(n738), .CO(n745), .S(n776) );
  CMPR32X1 U1105 ( .A(n753), .B(n752), .C(n751), .CO(n744), .S(n781) );
  OR2X2 U1106 ( .A(n766), .B(n765), .Y(n1138) );
  NAND2XL U1107 ( .A(n1138), .B(n770), .Y(mult_x_1_n295) );
  INVXL U1108 ( .A(mult_x_1_n307), .Y(n768) );
  AOI21XL U1109 ( .A0(n1138), .A1(n768), .B0(n767), .Y(mult_x_1_n296) );
  NAND2XL U1110 ( .A(n770), .B(mult_x_1_n307), .Y(mult_x_1_n84) );
  OAI21XL U1111 ( .A0(n772), .A1(n789), .B0(n771), .Y(n773) );
  AOI21XL U1112 ( .A0(n775), .A1(n774), .B0(n773), .Y(n1136) );
  INVXL U1113 ( .A(n1136), .Y(mult_x_1_n321) );
  AOI21XL U1114 ( .A0(mult_x_1_n321), .A1(n1175), .B0(n1133), .Y(mult_x_1_n316) );
  INVXL U1115 ( .A(n788), .Y(n790) );
  NAND2XL U1116 ( .A(n790), .B(n789), .Y(n791) );
  INVXL U1117 ( .A(n793), .Y(n802) );
  AOI21XL U1118 ( .A0(n802), .A1(n800), .B0(n794), .Y(n798) );
  XOR2X1 U1119 ( .A(n798), .B(n797), .Y(n1395) );
  NAND2XL U1120 ( .A(n800), .B(n799), .Y(n801) );
  XNOR2X1 U1121 ( .A(n802), .B(n801), .Y(n1396) );
  XNOR2XL U1122 ( .A(n991), .B(n1185), .Y(n820) );
  OAI22XL U1123 ( .A0(n1040), .A1(n820), .B0(n1038), .B1(n806), .Y(n838) );
  XNOR2X1 U1124 ( .A(n1224), .B(n945), .Y(n807) );
  XNOR2X1 U1125 ( .A(n1021), .B(n988), .Y(n824) );
  XNOR2X1 U1126 ( .A(B[1]), .B(A[24]), .Y(n828) );
  OAI22X1 U1127 ( .A0(n1027), .A1(n828), .B0(n813), .B1(n827), .Y(n826) );
  XNOR2X1 U1128 ( .A(n1224), .B(n985), .Y(n814) );
  NOR2XL U1129 ( .A(n1030), .B(n814), .Y(n825) );
  XNOR2X1 U1130 ( .A(n816), .B(n815), .Y(n839) );
  CMPR32X1 U1131 ( .A(n823), .B(n822), .C(n821), .CO(n850), .S(n859) );
  XNOR2X1 U1132 ( .A(n1021), .B(n949), .Y(n876) );
  OAI22X1 U1133 ( .A0(n1027), .A1(n879), .B0(n828), .B1(n827), .Y(n878) );
  XNOR2X1 U1134 ( .A(n1224), .B(n972), .Y(n829) );
  NOR2XL U1135 ( .A(n1030), .B(n829), .Y(n877) );
  CMPR32X1 U1136 ( .A(n832), .B(n831), .C(n830), .CO(n847), .S(n865) );
  OAI22XL U1137 ( .A0(n1061), .A1(n870), .B0(n1011), .B1(n833), .Y(n875) );
  OAI22XL U1138 ( .A0(n1205), .A1(n872), .B0(n1067), .B1(n835), .Y(n873) );
  CMPR32X1 U1139 ( .A(n838), .B(n837), .C(n836), .CO(n832), .S(n862) );
  CMPR32X1 U1140 ( .A(n841), .B(n840), .C(n839), .CO(n830), .S(n861) );
  ADDFHX1 U1141 ( .A(n847), .B(n846), .CI(n845), .CO(mult_x_1_n507), .S(
        mult_x_1_n508) );
  CMPR32X1 U1142 ( .A(n857), .B(n856), .C(n855), .CO(n858), .S(n893) );
  ADDFHX1 U1143 ( .A(n860), .B(n859), .CI(n858), .CO(n866), .S(n897) );
  CMPR32X1 U1144 ( .A(n863), .B(n862), .C(n861), .CO(n864), .S(n896) );
  ADDFHX1 U1145 ( .A(n869), .B(n868), .CI(n867), .CO(mult_x_1_n521), .S(
        mult_x_1_n522) );
  XNOR2X1 U1146 ( .A(n1187), .B(n1020), .Y(n904) );
  OAI22XL U1147 ( .A0(n1205), .A1(n904), .B0(n1067), .B1(n872), .Y(n905) );
  CMPR32X1 U1148 ( .A(n875), .B(n874), .C(n873), .CO(n863), .S(n891) );
  XNOR2X1 U1149 ( .A(B[9]), .B(n990), .Y(n908) );
  XNOR2X1 U1150 ( .A(B[1]), .B(n1201), .Y(n911) );
  NOR2XL U1151 ( .A(n1030), .B(n880), .Y(n909) );
  CMPR32X1 U1152 ( .A(n889), .B(n888), .C(n887), .CO(n890), .S(n924) );
  CMPR32X1 U1153 ( .A(n892), .B(n891), .C(n890), .CO(n901), .S(n928) );
  ADDFHX1 U1154 ( .A(n901), .B(n900), .CI(n899), .CO(mult_x_1_n537), .S(
        mult_x_1_n538) );
  XNOR2X1 U1155 ( .A(n1214), .B(n972), .Y(n934) );
  XNOR2X1 U1156 ( .A(n1187), .B(n945), .Y(n935) );
  OAI22XL U1157 ( .A0(n1016), .A1(n935), .B0(n1067), .B1(n904), .Y(n936) );
  OAI22XL U1158 ( .A0(n214), .A1(n939), .B0(n1072), .B1(n908), .Y(n920) );
  ADDHXL U1159 ( .A(n910), .B(n909), .CO(n887), .S(n919) );
  OAI22X1 U1160 ( .A0(n1027), .A1(n943), .B0(n911), .B1(n1123), .Y(n942) );
  XNOR2XL U1161 ( .A(n1224), .B(n970), .Y(n912) );
  NOR2XL U1162 ( .A(n1030), .B(n912), .Y(n941) );
  XNOR2X1 U1163 ( .A(n986), .B(n1020), .Y(n946) );
  XNOR2X1 U1164 ( .A(n681), .B(n981), .Y(n948) );
  XNOR2X1 U1165 ( .A(n991), .B(n988), .Y(n950) );
  CMPR32X1 U1166 ( .A(n920), .B(n918), .C(n919), .CO(n921), .S(n959) );
  CMPR32X1 U1167 ( .A(n923), .B(n922), .C(n921), .CO(n932), .S(n963) );
  ADDFHX1 U1168 ( .A(n932), .B(n931), .CI(n930), .CO(mult_x_1_n553), .S(
        mult_x_1_n554) );
  XNOR2X1 U1169 ( .A(n1214), .B(n1014), .Y(n971) );
  XNOR2X1 U1170 ( .A(n1187), .B(n985), .Y(n973) );
  OAI22XL U1171 ( .A0(n1016), .A1(n973), .B0(n1067), .B1(n935), .Y(n974) );
  XNOR2X1 U1172 ( .A(n1021), .B(A[13]), .Y(n978) );
  OAI22XL U1173 ( .A0(n214), .A1(n978), .B0(n1072), .B1(n939), .Y(n955) );
  XNOR2X1 U1174 ( .A(B[1]), .B(n1158), .Y(n982) );
  XNOR2XL U1175 ( .A(n1224), .B(n1012), .Y(n944) );
  NOR2XL U1176 ( .A(n1030), .B(n944), .Y(n979) );
  XNOR2X1 U1177 ( .A(n986), .B(n945), .Y(n987) );
  XNOR2X1 U1178 ( .A(n991), .B(n949), .Y(n992) );
  CMPR32X1 U1179 ( .A(n955), .B(n954), .C(n953), .CO(n956), .S(n1001) );
  ADDFHX1 U1180 ( .A(n961), .B(n960), .CI(n959), .CO(n964), .S(n1004) );
  ADDFHX1 U1181 ( .A(n964), .B(n963), .CI(n962), .CO(n931), .S(n965) );
  ADDFHX1 U1182 ( .A(n967), .B(n966), .CI(n965), .CO(mult_x_1_n569), .S(
        mult_x_1_n570) );
  OAI22XL U1183 ( .A0(n1061), .A1(n1010), .B0(n1011), .B1(n969), .Y(n1019) );
  XNOR2X1 U1184 ( .A(n1214), .B(n970), .Y(n1013) );
  OAI22XL U1185 ( .A0(n1016), .A1(n1015), .B0(n1067), .B1(n973), .Y(n1017) );
  CMPR32X1 U1186 ( .A(n976), .B(n975), .C(n974), .CO(n958), .S(n999) );
  XNOR2XL U1187 ( .A(n1021), .B(n977), .Y(n1022) );
  OAI22XL U1188 ( .A0(n214), .A1(n1022), .B0(n1072), .B1(n978), .Y(n997) );
  ADDHXL U1189 ( .A(n980), .B(n979), .CO(n953), .S(n996) );
  XNOR2X1 U1190 ( .A(B[1]), .B(n981), .Y(n1025) );
  OAI22X1 U1191 ( .A0(n1027), .A1(n1025), .B0(n982), .B1(n1123), .Y(n1024) );
  XNOR2X1 U1192 ( .A(n681), .B(n988), .Y(n1034) );
  XNOR2X1 U1193 ( .A(n991), .B(n990), .Y(n1037) );
  CMPR32X1 U1194 ( .A(n997), .B(n995), .C(n996), .CO(n998), .S(n1050) );
  CMPR32X1 U1195 ( .A(n1003), .B(n1002), .C(n1001), .CO(n1006), .S(n1053) );
  ADDFHX1 U1196 ( .A(n1009), .B(n1008), .CI(n1007), .CO(mult_x_1_n585), .S(
        mult_x_1_n586) );
  OAI22X1 U1197 ( .A0(n1061), .A1(n1059), .B0(n1011), .B1(n1010), .Y(n1070) );
  XNOR2X1 U1198 ( .A(n1214), .B(n1012), .Y(n1062) );
  XNOR2X1 U1199 ( .A(n1187), .B(n1014), .Y(n1066) );
  OAI22XL U1200 ( .A0(n1016), .A1(n1066), .B0(n1067), .B1(n1015), .Y(n1069) );
  CMPR32X1 U1201 ( .A(n1019), .B(n1018), .C(n1017), .CO(n1000), .S(n1048) );
  XNOR2XL U1202 ( .A(n1021), .B(n1020), .Y(n1071) );
  OAI22XL U1203 ( .A0(n214), .A1(n1071), .B0(n1072), .B1(n1022), .Y(n1046) );
  XNOR2XL U1204 ( .A(n1224), .B(n1028), .Y(n1029) );
  NOR2XL U1205 ( .A(n1030), .B(n1029), .Y(n1074) );
  CMPR32X1 U1206 ( .A(n1046), .B(n1045), .C(n1044), .CO(n1047), .S(n1090) );
  ADDFHX1 U1207 ( .A(n1058), .B(n1057), .CI(n1056), .CO(mult_x_1_n601), .S(
        mult_x_1_n602) );
  OAI22XL U1208 ( .A0(n214), .A1(n1073), .B0(n1072), .B1(n1071), .Y(n1086) );
  ADDHXL U1209 ( .A(n1075), .B(n1074), .CO(n1044), .S(n1085) );
  CMPR32X1 U1210 ( .A(n1083), .B(n1082), .C(n1081), .CO(n1092), .S(n1115) );
  CMPR32X1 U1211 ( .A(n1086), .B(n1084), .C(n1085), .CO(n1087), .S(n1114) );
  ADDFHX1 U1212 ( .A(n1092), .B(n1091), .CI(n1090), .CO(n1095), .S(n1117) );
  CMPR32X1 U1213 ( .A(n1107), .B(n1106), .C(n1105), .CO(n1111), .S(n1108) );
  CMPR32X1 U1214 ( .A(n1116), .B(n1115), .C(n1114), .CO(n1119), .S(n1144) );
  ADDFHX1 U1215 ( .A(n1122), .B(n1121), .CI(n1120), .CO(mult_x_1_n633), .S(
        mult_x_1_n634) );
  NAND2XL U1216 ( .A(n1138), .B(n1137), .Y(mult_x_1_n83) );
  CMPR32X1 U1217 ( .A(n1141), .B(n1140), .C(n1139), .CO(n1149), .S(n1152) );
  ADDFHX1 U1218 ( .A(n1149), .B(n1148), .CI(n1147), .CO(mult_x_1_n649), .S(
        n1154) );
  NOR2XL U1219 ( .A(n1154), .B(n1153), .Y(mult_x_1_n276) );
  NAND2XL U1220 ( .A(n1154), .B(n1153), .Y(mult_x_1_n277) );
  XNOR2X1 U1221 ( .A(n1187), .B(A[24]), .Y(n1188) );
  CMPR32X1 U1222 ( .A(n1168), .B(n1167), .C(n1166), .CO(n1189), .S(n1157) );
  CMPR32X1 U1223 ( .A(n1171), .B(n1170), .C(n1169), .CO(n1178), .S(n1156) );
  NAND2XL U1224 ( .A(n1173), .B(n1172), .Y(mult_x_1_n85) );
  NAND2XL U1225 ( .A(n1175), .B(n1174), .Y(mult_x_1_n86) );
  CMPR32X1 U1226 ( .A(n1183), .B(n1182), .C(n1181), .CO(n1196), .S(n1180) );
  XNOR2X1 U1227 ( .A(n1187), .B(A[25]), .Y(n1203) );
  OAI22X1 U1228 ( .A0(n1205), .A1(n1188), .B0(n1206), .B1(n1203), .Y(n1218) );
  CMPR32X1 U1229 ( .A(n1191), .B(n1190), .C(n1189), .CO(n1194), .S(n1179) );
  CMPR32X1 U1230 ( .A(n1196), .B(n1195), .C(n1194), .CO(n1208), .S(n1192) );
  CMPR32X1 U1231 ( .A(n1200), .B(n1199), .C(n1198), .CO(n1210), .S(n1195) );
  OAI2BB1X1 U1232 ( .A0N(n1206), .A1N(n1205), .B0(n1204), .Y(n1216) );
  CMPR32X1 U1233 ( .A(n1211), .B(n1210), .C(n1209), .CO(n1220), .S(n1207) );
  XNOR2X1 U1234 ( .A(n1214), .B(A[25]), .Y(n1227) );
  CMPR32X1 U1235 ( .A(n1218), .B(n1217), .C(n1216), .CO(n1221), .S(n1209) );
  CMPR32X1 U1236 ( .A(n1223), .B(n1222), .C(n1221), .CO(n1235), .S(n1219) );
  XOR3X2 U1237 ( .A(n1233), .B(n1232), .C(n1231), .Y(n1234) );
  OAI21XL U1238 ( .A0(n1243), .A1(n1338), .B0(n1242), .Y(n1307) );
  OAI21XL U1239 ( .A0(n1314), .A1(n1247), .B0(n1246), .Y(n1249) );
  OAI21XL U1240 ( .A0(n1314), .A1(n1253), .B0(n1252), .Y(n1256) );
  OAI21XL U1241 ( .A0(n1266), .A1(n1263), .B0(n1264), .Y(n1262) );
  INVXL U1242 ( .A(n1258), .Y(n1260) );
  OAI21XL U1243 ( .A0(n1329), .A1(n1332), .B0(n1330), .Y(n1276) );
  OAI21XL U1244 ( .A0(n1314), .A1(n1269), .B0(n1268), .Y(n1271) );
  OAI21XL U1245 ( .A0(n1314), .A1(n1281), .B0(n1280), .Y(n1284) );
  XNOR2XL U1246 ( .A(n1300), .B(n1299), .Y(n1400) );
  OAI21XL U1247 ( .A0(n1304), .A1(n1325), .B0(n1326), .Y(n1305) );
  OAI21XL U1248 ( .A0(n1310), .A1(n1309), .B0(n1308), .Y(n1311) );
  OAI21XL U1249 ( .A0(n1314), .A1(n1313), .B0(n1312), .Y(n1315) );
  XNOR2XL U1250 ( .A(n1315), .B(n1324), .Y(PRODUCT[40]) );
  XOR2XL U1251 ( .A(n1320), .B(n1319), .Y(n1399) );
endmodule


module FFT2048_DW02_mult_2_stage_J1_0 ( A, B, TC, CLK, PRODUCT );
  input [25:0] A;
  input [16:0] B;
  output [42:0] PRODUCT;
  input TC, CLK;
  wire   n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, mult_x_1_n309, mult_x_1_n308,
         mult_x_1_n301, mult_x_1_n294, mult_x_1_n291, mult_x_1_n290,
         mult_x_1_n287, mult_x_1_n286, mult_x_1_n282, mult_x_1_n281,
         mult_x_1_n277, mult_x_1_n276, mult_x_1_n274, mult_x_1_n273,
         mult_x_1_n266, mult_x_1_n265, mult_x_1_n263, mult_x_1_n262,
         mult_x_1_n252, mult_x_1_n251, mult_x_1_n245, mult_x_1_n244,
         mult_x_1_n234, mult_x_1_n233, mult_x_1_n227, mult_x_1_n226,
         mult_x_1_n216, mult_x_1_n215, mult_x_1_n207, mult_x_1_n206,
         mult_x_1_n198, mult_x_1_n197, mult_x_1_n195, mult_x_1_n194,
         mult_x_1_n184, mult_x_1_n183, mult_x_1_n177, mult_x_1_n176,
         mult_x_1_n170, mult_x_1_n169, mult_x_1_n161, mult_x_1_n160,
         mult_x_1_n152, mult_x_1_n151, mult_x_1_n137, mult_x_1_n136,
         mult_x_1_n130, mult_x_1_n129, mult_x_1_n121, mult_x_1_n120,
         mult_x_1_n110, mult_x_1_n109, mult_x_1_n84, mult_x_1_n83,
         mult_x_1_n82, mult_x_1_n58, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303;

  DFFHQXL mult_x_1_clk_r_REG9_S1 ( .D(mult_x_1_n197), .CK(CLK), .Q(n1270) );
  DFFHQXL mult_x_1_clk_r_REG17_S1 ( .D(mult_x_1_n169), .CK(CLK), .Q(n1262) );
  DFFHQX4 mult_x_1_clk_r_REG48_S1 ( .D(mult_x_1_n291), .CK(CLK), .Q(n1300) );
  DFFHQX4 mult_x_1_clk_r_REG49_S1 ( .D(mult_x_1_n290), .CK(CLK), .Q(n1296) );
  DFFHQX4 mult_x_1_clk_r_REG45_S1 ( .D(mult_x_1_n287), .CK(CLK), .Q(n1295) );
  DFFHQX4 mult_x_1_clk_r_REG44_S1 ( .D(mult_x_1_n281), .CK(CLK), .Q(n1292) );
  DFFHQX4 mult_x_1_clk_r_REG42_S1 ( .D(mult_x_1_n276), .CK(CLK), .Q(n1290) );
  DFFHQX4 mult_x_1_clk_r_REG40_S1 ( .D(mult_x_1_n273), .CK(CLK), .Q(n1288) );
  DFFHQX4 mult_x_1_clk_r_REG37_S1 ( .D(mult_x_1_n266), .CK(CLK), .Q(n1287) );
  DFFHQX4 mult_x_1_clk_r_REG38_S1 ( .D(mult_x_1_n265), .CK(CLK), .Q(n1286) );
  DFFHQX4 mult_x_1_clk_r_REG36_S1 ( .D(mult_x_1_n262), .CK(CLK), .Q(n1284) );
  DFFHQX4 mult_x_1_clk_r_REG33_S1 ( .D(mult_x_1_n252), .CK(CLK), .Q(n1283) );
  DFFHQX4 mult_x_1_clk_r_REG34_S1 ( .D(mult_x_1_n251), .CK(CLK), .Q(n1282) );
  DFFHQX2 mult_x_1_clk_r_REG31_S1 ( .D(mult_x_1_n245), .CK(CLK), .Q(n1281) );
  DFFHQX4 mult_x_1_clk_r_REG0_S1 ( .D(mult_x_1_n234), .CK(CLK), .Q(n1279) );
  DFFHQX4 mult_x_1_clk_r_REG3_S1 ( .D(mult_x_1_n226), .CK(CLK), .Q(n1276) );
  DFFHQX4 mult_x_1_clk_r_REG5_S1 ( .D(mult_x_1_n215), .CK(CLK), .Q(n1274) );
  DFFHQXL mult_x_1_clk_r_REG6_S1 ( .D(mult_x_1_n207), .CK(CLK), .Q(n1273) );
  DFFHQX4 mult_x_1_clk_r_REG7_S1 ( .D(mult_x_1_n206), .CK(CLK), .Q(n1272) );
  DFFHQXL clk_r_REG54_S1 ( .D(n1318), .CK(CLK), .Q(PRODUCT[13]) );
  DFFHQX4 mult_x_1_clk_r_REG55_S1 ( .D(mult_x_1_n309), .CK(CLK), .Q(n1303) );
  DFFHQXL mult_x_1_clk_r_REG51_S1 ( .D(mult_x_1_n294), .CK(CLK), .Q(n1301) );
  DFFHQXL mult_x_1_clk_r_REG10_S1 ( .D(mult_x_1_n195), .CK(CLK), .Q(n1269) );
  DFFHQXL mult_x_1_clk_r_REG14_S1 ( .D(mult_x_1_n177), .CK(CLK), .Q(n1265) );
  DFFHQXL clk_r_REG58_S1 ( .D(n1320), .CK(CLK), .Q(PRODUCT[11]) );
  DFFHQX4 mult_x_1_clk_r_REG35_S1 ( .D(mult_x_1_n263), .CK(CLK), .Q(n1285) );
  DFFHQXL mult_x_1_clk_r_REG50_S1 ( .D(mult_x_1_n83), .CK(CLK), .Q(n1298) );
  DFFHQXL mult_x_1_clk_r_REG15_S1 ( .D(mult_x_1_n176), .CK(CLK), .Q(n1264) );
  DFFHQXL clk_r_REG57_S1 ( .D(n1319), .CK(CLK), .Q(PRODUCT[12]) );
  DFFHQXL mult_x_1_clk_r_REG16_S1 ( .D(mult_x_1_n170), .CK(CLK), .Q(n1263) );
  DFFHQXL mult_x_1_clk_r_REG47_S1 ( .D(mult_x_1_n82), .CK(CLK), .Q(n1297) );
  DFFHQXL clk_r_REG67_S1 ( .D(n1329), .CK(CLK), .Q(PRODUCT[2]) );
  DFFHQXL mult_x_1_clk_r_REG18_S1 ( .D(mult_x_1_n161), .CK(CLK), .Q(n1261) );
  DFFHQX4 mult_x_1_clk_r_REG2_S1 ( .D(mult_x_1_n227), .CK(CLK), .Q(n1277) );
  DFFHQX1 mult_x_1_clk_r_REG4_S1 ( .D(mult_x_1_n216), .CK(CLK), .Q(n1275) );
  DFFHQXL mult_x_1_clk_r_REG53_S1 ( .D(mult_x_1_n301), .CK(CLK), .Q(n1302) );
  DFFHQX2 mult_x_1_clk_r_REG46_S1 ( .D(mult_x_1_n286), .CK(CLK), .Q(n1294) );
  DFFHQXL clk_r_REG59_S1 ( .D(n1321), .CK(CLK), .Q(PRODUCT[10]) );
  DFFHQXL clk_r_REG60_S1 ( .D(n1322), .CK(CLK), .Q(PRODUCT[9]) );
  DFFHQXL clk_r_REG61_S1 ( .D(n1323), .CK(CLK), .Q(PRODUCT[8]) );
  DFFHQXL clk_r_REG62_S1 ( .D(n1324), .CK(CLK), .Q(PRODUCT[7]) );
  DFFHQXL clk_r_REG63_S1 ( .D(n1325), .CK(CLK), .Q(PRODUCT[6]) );
  DFFHQXL clk_r_REG64_S1 ( .D(n1326), .CK(CLK), .Q(PRODUCT[5]) );
  DFFHQXL clk_r_REG65_S1 ( .D(n1327), .CK(CLK), .Q(PRODUCT[4]) );
  DFFHQXL clk_r_REG66_S1 ( .D(n1328), .CK(CLK), .Q(PRODUCT[3]) );
  DFFHQXL clk_r_REG68_S1 ( .D(n1330), .CK(CLK), .Q(PRODUCT[1]) );
  DFFHQXL clk_r_REG69_S1 ( .D(n1331), .CK(CLK), .Q(PRODUCT[0]) );
  DFFHQXL mult_x_1_clk_r_REG13_S1 ( .D(mult_x_1_n183), .CK(CLK), .Q(n1266) );
  DFFHQX1 mult_x_1_clk_r_REG52_S1 ( .D(mult_x_1_n84), .CK(CLK), .Q(n1299) );
  DFFHQX1 mult_x_1_clk_r_REG8_S1 ( .D(mult_x_1_n198), .CK(CLK), .Q(n1271) );
  DFFHQXL mult_x_1_clk_r_REG12_S1 ( .D(mult_x_1_n184), .CK(CLK), .Q(n1267) );
  DFFHQXL mult_x_1_clk_r_REG20_S1 ( .D(mult_x_1_n152), .CK(CLK), .Q(n1259) );
  DFFHQXL mult_x_1_clk_r_REG22_S1 ( .D(mult_x_1_n137), .CK(CLK), .Q(n1257) );
  DFFHQXL mult_x_1_clk_r_REG23_S1 ( .D(mult_x_1_n136), .CK(CLK), .Q(n1256) );
  DFFHQXL mult_x_1_clk_r_REG24_S1 ( .D(mult_x_1_n130), .CK(CLK), .Q(n1255) );
  DFFHQXL mult_x_1_clk_r_REG25_S1 ( .D(mult_x_1_n129), .CK(CLK), .Q(n1254) );
  DFFHQXL mult_x_1_clk_r_REG26_S1 ( .D(mult_x_1_n121), .CK(CLK), .Q(n1253) );
  DFFHQXL mult_x_1_clk_r_REG27_S1 ( .D(mult_x_1_n120), .CK(CLK), .Q(n1252) );
  DFFHQXL mult_x_1_clk_r_REG28_S1 ( .D(mult_x_1_n110), .CK(CLK), .Q(n1251) );
  DFFHQXL mult_x_1_clk_r_REG29_S1 ( .D(mult_x_1_n109), .CK(CLK), .Q(n1250) );
  DFFHQXL mult_x_1_clk_r_REG30_S1 ( .D(mult_x_1_n58), .CK(CLK), .Q(n1249) );
  DFFHQXL mult_x_1_clk_r_REG56_S1 ( .D(mult_x_1_n308), .CK(CLK), .Q(n1248) );
  DFFHQXL mult_x_1_clk_r_REG21_S1 ( .D(mult_x_1_n151), .CK(CLK), .Q(n1258) );
  DFFHQXL mult_x_1_clk_r_REG19_S1 ( .D(mult_x_1_n160), .CK(CLK), .Q(n1260) );
  DFFHQXL mult_x_1_clk_r_REG11_S1 ( .D(mult_x_1_n194), .CK(CLK), .Q(n1268) );
  DFFHQX2 mult_x_1_clk_r_REG41_S1 ( .D(mult_x_1_n277), .CK(CLK), .Q(n1291) );
  DFFHQX1 mult_x_1_clk_r_REG39_S1 ( .D(mult_x_1_n274), .CK(CLK), .Q(n1289) );
  DFFHQX2 mult_x_1_clk_r_REG43_S1 ( .D(mult_x_1_n282), .CK(CLK), .Q(n1293) );
  DFFHQX1 mult_x_1_clk_r_REG1_S1 ( .D(mult_x_1_n233), .CK(CLK), .Q(n1278) );
  DFFHQX2 mult_x_1_clk_r_REG32_S1 ( .D(mult_x_1_n244), .CK(CLK), .Q(n1280) );
  ADDFX2 U1 ( .A(n796), .B(n795), .CI(n794), .CO(n783), .S(n825) );
  ADDFHX1 U2 ( .A(n676), .B(n675), .CI(n674), .CO(n672), .S(n706) );
  ADDFHX1 U3 ( .A(n634), .B(n633), .CI(n632), .CO(n591), .S(n635) );
  ADDFHX2 U4 ( .A(n704), .B(n703), .CI(n702), .CO(n675), .S(n715) );
  OAI21XL U5 ( .A0(n1095), .A1(n248), .B0(n247), .Y(mult_x_1_n309) );
  ADDFHX1 U6 ( .A(n1008), .B(n1007), .CI(n1006), .CO(n964), .S(n1014) );
  ADDFHX1 U7 ( .A(n1050), .B(n1049), .CI(n1048), .CO(n1040), .S(n1055) );
  ADDFHX2 U8 ( .A(n1005), .B(n1004), .CI(n1003), .CO(n1008), .S(n1029) );
  ADDFHX2 U9 ( .A(n948), .B(n947), .CI(n946), .CO(n965), .S(n1007) );
  ADDFX2 U10 ( .A(n899), .B(n898), .CI(n897), .CO(n910), .S(n953) );
  ADDFX2 U11 ( .A(n652), .B(n651), .CI(n650), .CO(n631), .S(n676) );
  OAI21XL U12 ( .A0(n905), .A1(n904), .B0(n903), .Y(n32) );
  ADDFX2 U13 ( .A(n701), .B(n700), .CI(n699), .CO(n704), .S(n744) );
  ADDFHX1 U14 ( .A(n538), .B(n537), .CI(n536), .CO(n531), .S(n588) );
  CMPR32X1 U15 ( .A(n817), .B(n816), .C(n815), .CO(n832), .S(n863) );
  CMPR32X1 U16 ( .A(n896), .B(n895), .C(n894), .CO(n897), .S(n949) );
  ADDFHX1 U17 ( .A(n1047), .B(n1046), .CI(n1045), .CO(n1056), .S(n1058) );
  ADDFX2 U18 ( .A(n516), .B(n515), .CI(n514), .CO(n535), .S(n551) );
  ADDFHX1 U19 ( .A(n331), .B(n330), .CI(n329), .CO(n1059), .S(n346) );
  ADDFHX1 U20 ( .A(n802), .B(n801), .CI(n800), .CO(n776), .S(n816) );
  CMPR32X1 U21 ( .A(n987), .B(n986), .C(n985), .CO(n1025), .S(n1021) );
  OAI22X1 U22 ( .A0(n1146), .A1(n837), .B0(n1147), .B1(n798), .Y(n840) );
  ADDFHX1 U23 ( .A(n302), .B(n301), .CI(n300), .CO(n329), .S(n311) );
  ADDFHX1 U24 ( .A(n314), .B(n313), .CI(n312), .CO(n1065), .S(n245) );
  ADDFHX1 U25 ( .A(n334), .B(n333), .CI(n332), .CO(n1047), .S(n330) );
  OAI22X2 U26 ( .A0(n1146), .A1(n9), .B0(n621), .B1(n1147), .Y(n680) );
  ADDFHX1 U27 ( .A(n233), .B(n232), .CI(n231), .CO(n313), .S(n234) );
  BUFX8 U28 ( .A(n266), .Y(n1147) );
  BUFX8 U29 ( .A(n265), .Y(n1146) );
  BUFX4 U30 ( .A(n337), .Y(n1143) );
  ADDFHX1 U31 ( .A(n193), .B(n192), .CI(n191), .CO(n194), .S(n155) );
  ADDFHX1 U32 ( .A(n224), .B(n223), .CI(n222), .CO(n279), .S(n225) );
  ADDFHX1 U33 ( .A(n181), .B(n180), .CI(n179), .CO(n229), .S(n190) );
  ADDFHX2 U34 ( .A(n143), .B(n142), .CI(n141), .CO(n192), .S(n145) );
  NAND2X1 U35 ( .A(n264), .B(n266), .Y(n265) );
  INVX2 U36 ( .A(B[15]), .Y(n354) );
  BUFX4 U37 ( .A(n595), .Y(n939) );
  CLKBUFX8 U38 ( .A(n122), .Y(n977) );
  BUFX8 U39 ( .A(B[9]), .Y(n911) );
  BUFX8 U40 ( .A(B[7]), .Y(n833) );
  CLKBUFX8 U41 ( .A(B[5]), .Y(n913) );
  NAND2X1 U42 ( .A(n62), .B(n973), .Y(n67) );
  XNOR2X1 U43 ( .A(n259), .B(n258), .Y(PRODUCT[27]) );
  XNOR2X1 U44 ( .A(n793), .B(n792), .Y(PRODUCT[24]) );
  OAI21XL U45 ( .A0(n1089), .A1(n256), .B0(n255), .Y(n259) );
  BUFX4 U46 ( .A(n394), .Y(n1246) );
  OAI22X1 U47 ( .A0(n654), .A1(n432), .B0(n566), .B1(n427), .Y(n441) );
  AOI21XL U48 ( .A0(n487), .A1(n396), .B0(n395), .Y(n1242) );
  XNOR2XL U49 ( .A(n353), .B(n352), .Y(PRODUCT[25]) );
  XNOR2XL U50 ( .A(n1302), .B(n1298), .Y(PRODUCT[15]) );
  XNOR2XL U51 ( .A(n911), .B(A[2]), .Y(n162) );
  BUFX1 U52 ( .A(n654), .Y(n49) );
  XNOR2XL U53 ( .A(n920), .B(A[22]), .Y(n507) );
  XNOR2XL U54 ( .A(n765), .B(A[4]), .Y(n70) );
  XNOR2XL U55 ( .A(n765), .B(A[13]), .Y(n324) );
  XNOR2XL U56 ( .A(n920), .B(A[23]), .Y(n469) );
  BUFX3 U57 ( .A(n198), .Y(n5) );
  ADDFX2 U58 ( .A(n773), .B(n772), .CI(n771), .CO(n774), .S(n818) );
  INVX1 U59 ( .A(B[0]), .Y(n761) );
  XOR2XL U60 ( .A(n1197), .B(n1196), .Y(n1325) );
  XNOR2XL U61 ( .A(n1099), .B(n1098), .Y(n1319) );
  OAI21XL U62 ( .A0(n1093), .A1(n1092), .B0(n1063), .Y(mult_x_1_n291) );
  OAI22X1 U63 ( .A0(n323), .A1(n163), .B0(n977), .B1(n162), .Y(n173) );
  XOR2X1 U64 ( .A(n1179), .B(n1178), .Y(n1322) );
  XNOR2X1 U65 ( .A(n1182), .B(n1181), .Y(n1323) );
  INVX1 U66 ( .A(n1070), .Y(n1097) );
  NAND2X1 U67 ( .A(n245), .B(n244), .Y(n1071) );
  NAND2X1 U68 ( .A(n7), .B(n6), .Y(n483) );
  INVX1 U69 ( .A(n1180), .Y(n1175) );
  NAND2X1 U70 ( .A(n153), .B(n152), .Y(n1180) );
  OR2X2 U71 ( .A(n153), .B(n152), .Y(n151) );
  NAND2X1 U72 ( .A(n117), .B(n116), .Y(n1194) );
  NOR2X1 U73 ( .A(n1143), .B(n927), .Y(n980) );
  NOR2X1 U74 ( .A(n1143), .B(n1131), .Y(n1141) );
  NOR2X1 U75 ( .A(n1143), .B(n1122), .Y(n1135) );
  NOR2X1 U76 ( .A(n1143), .B(n969), .Y(n998) );
  NOR2X1 U77 ( .A(n1143), .B(n355), .Y(n378) );
  NOR2X1 U78 ( .A(n1143), .B(n453), .Y(n474) );
  BUFX8 U79 ( .A(n323), .Y(n979) );
  NOR2X1 U80 ( .A(n1143), .B(n403), .Y(n438) );
  NOR2BX1 U81 ( .AN(A[0]), .B(n937), .Y(n113) );
  XOR2X1 U82 ( .A(n426), .B(n21), .Y(PRODUCT[34]) );
  NOR2X1 U83 ( .A(n1235), .B(n1162), .Y(n1199) );
  NAND2X1 U84 ( .A(n486), .B(n396), .Y(n1235) );
  NAND2X1 U85 ( .A(n450), .B(n1263), .Y(n451) );
  INVX1 U86 ( .A(n1258), .Y(n1157) );
  INVX1 U87 ( .A(n1266), .Y(n527) );
  INVX1 U88 ( .A(n1252), .Y(n1201) );
  INVX1 U89 ( .A(n1294), .Y(n1035) );
  XNOR2X1 U90 ( .A(n1192), .B(n1191), .Y(n1324) );
  NAND2X1 U91 ( .A(n243), .B(n242), .Y(n1096) );
  INVX1 U92 ( .A(n589), .Y(n46) );
  ADDFHX2 U93 ( .A(n619), .B(n618), .CI(n617), .CO(n649), .S(n670) );
  NAND2XL U94 ( .A(n440), .B(n441), .Y(n6) );
  NOR2X1 U95 ( .A(n117), .B(n116), .Y(n1193) );
  ADDFHX1 U96 ( .A(n814), .B(n813), .CI(n812), .CO(n815), .S(n859) );
  NOR2X1 U97 ( .A(n1143), .B(n402), .Y(n416) );
  NOR2X1 U98 ( .A(n1143), .B(n357), .Y(n368) );
  NOR2X1 U99 ( .A(n1143), .B(n1107), .Y(n1120) );
  NOR2X1 U100 ( .A(n1143), .B(n372), .Y(n1105) );
  NOR2X1 U101 ( .A(n1143), .B(n728), .Y(n759) );
  NOR2X1 U102 ( .A(n1143), .B(n846), .Y(n880) );
  NOR2X1 U103 ( .A(n1143), .B(n430), .Y(n458) );
  XNOR2XL U104 ( .A(n1132), .B(A[24]), .Y(n1133) );
  XNOR2X1 U105 ( .A(n1210), .B(n1209), .Y(PRODUCT[39]) );
  XNOR2X1 U106 ( .A(n400), .B(n399), .Y(PRODUCT[35]) );
  NAND2X1 U107 ( .A(n257), .B(n1275), .Y(n258) );
  NAND2X1 U108 ( .A(n867), .B(n1285), .Y(n868) );
  NAND2X1 U109 ( .A(n592), .B(n1271), .Y(n593) );
  INVX1 U110 ( .A(n1282), .Y(n788) );
  OAI21XL U111 ( .A0(n1272), .A1(n1275), .B0(n1273), .Y(n40) );
  INVX1 U112 ( .A(n1278), .Y(n351) );
  INVX1 U113 ( .A(n1260), .Y(n1155) );
  XNOR2X1 U114 ( .A(n1301), .B(n1297), .Y(PRODUCT[16]) );
  XOR2X1 U115 ( .A(n1248), .B(n1299), .Y(PRODUCT[14]) );
  INVX1 U116 ( .A(mult_x_1_n309), .Y(mult_x_1_n308) );
  NAND2XL U117 ( .A(n19), .B(n18), .Y(n17) );
  NAND2XL U118 ( .A(n648), .B(n649), .Y(n16) );
  NAND2X1 U119 ( .A(n1066), .B(n1065), .Y(n1068) );
  INVXL U120 ( .A(n648), .Y(n19) );
  OR2XL U121 ( .A(n1152), .B(n1151), .Y(n1154) );
  INVXL U122 ( .A(n649), .Y(n18) );
  OAI2BB1XL U123 ( .A0N(n811), .A1N(n30), .B0(n26), .Y(n820) );
  INVXL U124 ( .A(n588), .Y(n45) );
  XOR2X1 U125 ( .A(n238), .B(n237), .Y(n54) );
  ADDFHX2 U126 ( .A(n308), .B(n307), .CI(n306), .CO(n347), .S(n309) );
  ADDFHX1 U127 ( .A(n951), .B(n950), .CI(n949), .CO(n954), .S(n1006) );
  ADDFHX1 U128 ( .A(n855), .B(n854), .CI(n853), .CO(n856), .S(n900) );
  ADDFHX1 U129 ( .A(n178), .B(n177), .CI(n176), .CO(n185), .S(n193) );
  ADDFHX1 U130 ( .A(n723), .B(n722), .CI(n721), .CO(n698), .S(n739) );
  ADDFHX1 U131 ( .A(n757), .B(n756), .CI(n755), .CO(n740), .S(n775) );
  OAI2BB1XL U132 ( .A0N(n835), .A1N(n836), .B0(n405), .Y(n436) );
  ADDFHX1 U133 ( .A(n681), .B(n680), .CI(n679), .CO(n668), .S(n697) );
  INVXL U134 ( .A(n30), .Y(n28) );
  ADDFHX1 U135 ( .A(n841), .B(n840), .CI(n839), .CO(n817), .S(n857) );
  ADDFHX1 U136 ( .A(n984), .B(n983), .CI(n982), .CO(n951), .S(n1017) );
  ADDFHX1 U137 ( .A(n996), .B(n995), .CI(n994), .CO(n1044), .S(n1026) );
  NAND2BX1 U138 ( .AN(n806), .B(n35), .Y(n34) );
  AND2XL U139 ( .A(n1217), .B(n1218), .Y(n1330) );
  NOR2X1 U140 ( .A(n1143), .B(n502), .Y(n563) );
  NOR2XL U141 ( .A(n1143), .B(n1142), .Y(n1149) );
  XNOR2XL U142 ( .A(n501), .B(A[17]), .Y(n402) );
  XNOR2XL U143 ( .A(n501), .B(A[23]), .Y(n1131) );
  XNOR2XL U144 ( .A(n501), .B(A[24]), .Y(n1142) );
  XNOR2XL U145 ( .A(n501), .B(A[21]), .Y(n1107) );
  XNOR2XL U146 ( .A(n501), .B(A[20]), .Y(n372) );
  XNOR2XL U147 ( .A(n501), .B(A[22]), .Y(n1122) );
  OR2XL U148 ( .A(n1216), .B(n1215), .Y(n1217) );
  XNOR2X1 U149 ( .A(n1166), .B(n1165), .Y(PRODUCT[36]) );
  XNOR2X1 U150 ( .A(n1173), .B(n1172), .Y(PRODUCT[37]) );
  XNOR2X1 U151 ( .A(n1186), .B(n1185), .Y(PRODUCT[38]) );
  INVXL U152 ( .A(n1243), .Y(n1244) );
  OR2XL U153 ( .A(n1235), .B(n1241), .Y(n1245) );
  NOR2X1 U154 ( .A(n40), .B(n39), .Y(n388) );
  INVX1 U155 ( .A(A[10]), .Y(n10) );
  INVXL U156 ( .A(A[3]), .Y(n15) );
  INVXL U157 ( .A(n1263), .Y(n37) );
  NAND2X1 U158 ( .A(n748), .B(n747), .Y(mult_x_1_n227) );
  OAI21X2 U159 ( .A0(n1288), .A1(n1291), .B0(n1289), .Y(n249) );
  XNOR2X2 U160 ( .A(n558), .B(n557), .Y(PRODUCT[30]) );
  OAI21X2 U161 ( .A0(n1276), .A1(n1279), .B0(n1277), .Y(n386) );
  OAI22X1 U162 ( .A0(n931), .A1(n169), .B0(n929), .B1(n201), .Y(n206) );
  OAI22X1 U163 ( .A0(n939), .A1(n165), .B0(n937), .B1(n204), .Y(n210) );
  NAND2X2 U164 ( .A(n65), .B(n72), .Y(n595) );
  XNOR2X1 U165 ( .A(n1132), .B(A[8]), .Y(n753) );
  OAI21XL U166 ( .A0(n440), .A1(n441), .B0(n439), .Y(n7) );
  XOR2X1 U167 ( .A(n8), .B(n439), .Y(n478) );
  XOR2X1 U168 ( .A(n440), .B(n441), .Y(n8) );
  XNOR2X4 U169 ( .A(B[12]), .B(B[11]), .Y(n198) );
  OAI22X2 U170 ( .A0(n1146), .A1(n719), .B0(n1147), .B1(n9), .Y(n722) );
  XOR2X2 U171 ( .A(n1132), .B(n10), .Y(n9) );
  NOR2X1 U172 ( .A(n245), .B(n244), .Y(n13) );
  NAND2XL U173 ( .A(n1071), .B(n11), .Y(n1072) );
  NAND2X1 U174 ( .A(n1097), .B(n11), .Y(n248) );
  INVX1 U175 ( .A(n13), .Y(n11) );
  NOR2X1 U176 ( .A(n246), .B(n12), .Y(n247) );
  NOR2X1 U177 ( .A(n13), .B(n1096), .Y(n12) );
  OAI22X1 U178 ( .A0(n979), .A1(n162), .B0(n977), .B1(n14), .Y(n209) );
  OAI22X1 U179 ( .A0(n979), .A1(n14), .B0(n219), .B1(n977), .Y(n227) );
  XOR2X1 U180 ( .A(n911), .B(n15), .Y(n14) );
  OAI2BB1X1 U181 ( .A0N(n17), .A1N(n647), .B0(n16), .Y(n636) );
  XOR2X2 U182 ( .A(n647), .B(n20), .Y(n673) );
  XOR2X2 U183 ( .A(n648), .B(n649), .Y(n20) );
  XNOR2X1 U184 ( .A(n968), .B(A[11]), .Y(n543) );
  AOI2BB1X2 U185 ( .A0N(n1095), .A1N(n1070), .B0(n1069), .Y(n1073) );
  XNOR2X1 U186 ( .A(n605), .B(n604), .Y(n626) );
  OAI22X1 U187 ( .A0(n1146), .A1(n621), .B0(n1147), .B1(n568), .Y(n604) );
  INVX1 U188 ( .A(n1143), .Y(n35) );
  OAI21XL U189 ( .A0(n1242), .A1(n1162), .B0(n1161), .Y(n1205) );
  INVXL U190 ( .A(n1239), .Y(n1161) );
  NAND2XL U191 ( .A(n66), .B(n890), .Y(n93) );
  XOR2XL U192 ( .A(B[2]), .B(B[3]), .Y(n66) );
  XNOR2X2 U193 ( .A(B[8]), .B(B[7]), .Y(n122) );
  BUFX4 U194 ( .A(n973), .Y(n835) );
  XNOR2XL U195 ( .A(B[2]), .B(B[1]), .Y(n890) );
  BUFX2 U196 ( .A(n93), .Y(n282) );
  INVXL U197 ( .A(n1261), .Y(n1158) );
  NAND2XL U198 ( .A(n1155), .B(n1157), .Y(n1160) );
  NAND2XL U199 ( .A(n1198), .B(n1201), .Y(n1233) );
  NOR2X1 U200 ( .A(n1278), .B(n1276), .Y(n637) );
  NOR2X1 U201 ( .A(n1274), .B(n1272), .Y(n387) );
  NOR2X1 U202 ( .A(n1286), .B(n1284), .Y(n785) );
  NOR2X1 U203 ( .A(n1282), .B(n1280), .Y(n254) );
  XNOR2XL U204 ( .A(n882), .B(A[13]), .Y(n288) );
  AOI21XL U205 ( .A0(n1202), .A1(n1201), .B0(n1200), .Y(n1236) );
  INVXL U206 ( .A(n1253), .Y(n1200) );
  INVXL U207 ( .A(n1233), .Y(n1204) );
  NAND2X1 U208 ( .A(n785), .B(n254), .Y(n385) );
  NAND2XL U209 ( .A(n1171), .B(n1255), .Y(n1172) );
  XNOR2X1 U210 ( .A(n885), .B(A[8]), .Y(n886) );
  XNOR2XL U211 ( .A(n882), .B(A[7]), .Y(n132) );
  ADDFX2 U212 ( .A(n175), .B(n174), .CI(n173), .CO(n230), .S(n186) );
  OAI22X1 U213 ( .A0(n926), .A1(n161), .B0(n160), .B1(n1085), .Y(n174) );
  NOR2BX1 U214 ( .AN(A[0]), .B(n929), .Y(n175) );
  NAND2XL U215 ( .A(n712), .B(n1277), .Y(n713) );
  OAI21XL U216 ( .A0(n1089), .A1(n711), .B0(n710), .Y(n714) );
  ADDFX2 U217 ( .A(n210), .B(n209), .CI(n208), .CO(n232), .S(n237) );
  OAI22XL U218 ( .A0(n654), .A1(n365), .B0(n566), .B1(n363), .Y(n369) );
  OAI22XL U219 ( .A0(n1146), .A1(n364), .B0(n1147), .B1(n361), .Y(n371) );
  OAI22XL U220 ( .A0(n1125), .A1(n401), .B0(n5), .B1(n362), .Y(n370) );
  OAI22X1 U221 ( .A0(n931), .A1(n764), .B0(n929), .B1(n729), .Y(n770) );
  NOR2X1 U222 ( .A(n48), .B(n47), .Y(n771) );
  INVXL U223 ( .A(n804), .Y(n47) );
  XNOR2XL U224 ( .A(n882), .B(A[4]), .Y(n98) );
  OAI22XL U225 ( .A0(n282), .A1(n167), .B0(n933), .B1(n170), .Y(n179) );
  OAI22X1 U226 ( .A0(n975), .A1(n164), .B0(n835), .B1(n168), .Y(n181) );
  OAI22X1 U227 ( .A0(n975), .A1(n133), .B0(n835), .B1(n164), .Y(n178) );
  OAI2BB1XL U228 ( .A0N(n5), .A1N(n1125), .B0(n1124), .Y(n1134) );
  INVXL U229 ( .A(n1123), .Y(n1124) );
  NAND2XL U230 ( .A(n1177), .B(n151), .Y(n157) );
  OAI22XL U231 ( .A0(n1146), .A1(n1133), .B0(n1147), .B1(n1144), .Y(n1150) );
  INVXL U232 ( .A(n390), .Y(n709) );
  INVX1 U233 ( .A(n385), .Y(n707) );
  NOR2XL U234 ( .A(n1256), .B(n1254), .Y(n1198) );
  NOR2X2 U235 ( .A(n1292), .B(n1294), .Y(n959) );
  INVXL U236 ( .A(n1199), .Y(n1164) );
  INVXL U237 ( .A(n1205), .Y(n1163) );
  INVXL U238 ( .A(n1256), .Y(n1168) );
  NAND2BXL U239 ( .AN(A[0]), .B(n885), .Y(n158) );
  XNOR2XL U240 ( .A(n882), .B(A[21]), .Y(n762) );
  XNOR2XL U241 ( .A(n882), .B(A[20]), .Y(n805) );
  XNOR2XL U242 ( .A(n882), .B(A[19]), .Y(n844) );
  XNOR2XL U243 ( .A(n882), .B(A[18]), .Y(n883) );
  XNOR2XL U244 ( .A(n882), .B(A[14]), .Y(n287) );
  XNOR2XL U245 ( .A(n882), .B(A[11]), .Y(n200) );
  XNOR2XL U246 ( .A(n913), .B(A[8]), .Y(n218) );
  XNOR2XL U247 ( .A(n913), .B(A[9]), .Y(n268) );
  XNOR2XL U248 ( .A(n911), .B(A[6]), .Y(n263) );
  XNOR2XL U249 ( .A(n882), .B(A[24]), .Y(n615) );
  XNOR2X1 U250 ( .A(n1108), .B(A[16]), .Y(n509) );
  XNOR2XL U251 ( .A(n882), .B(A[10]), .Y(n160) );
  AOI21XL U252 ( .A0(n36), .A1(n1155), .B0(n1158), .Y(n397) );
  INVXL U253 ( .A(n424), .Y(n36) );
  INVXL U254 ( .A(n1262), .Y(n450) );
  INVXL U255 ( .A(n1274), .Y(n257) );
  NAND2XL U256 ( .A(n1087), .B(n1287), .Y(n1088) );
  NOR2XL U257 ( .A(n1160), .B(n1262), .Y(n1234) );
  AOI21XL U258 ( .A0(n1158), .A1(n1157), .B0(n1156), .Y(n1159) );
  INVXL U259 ( .A(n1259), .Y(n1156) );
  NOR2XL U260 ( .A(n1233), .B(n1250), .Y(n1238) );
  NAND2XL U261 ( .A(n1199), .B(n1198), .Y(n1184) );
  XNOR2XL U262 ( .A(n913), .B(A[7]), .Y(n204) );
  INVXL U263 ( .A(n602), .Y(n574) );
  NOR2X1 U264 ( .A(n1143), .B(n686), .Y(n725) );
  XNOR2X1 U265 ( .A(n885), .B(A[12]), .Y(n729) );
  XNOR2X1 U266 ( .A(n885), .B(A[13]), .Y(n687) );
  XNOR2XL U267 ( .A(n913), .B(A[18]), .Y(n731) );
  XNOR2XL U268 ( .A(n913), .B(A[19]), .Y(n689) );
  XNOR2X1 U269 ( .A(n1132), .B(A[9]), .Y(n719) );
  NAND2BX1 U270 ( .AN(n763), .B(n35), .Y(n48) );
  OAI22X1 U271 ( .A0(n926), .A1(n805), .B0(n762), .B1(n761), .Y(n804) );
  INVXL U272 ( .A(n843), .Y(n33) );
  XNOR2XL U273 ( .A(n911), .B(A[13]), .Y(n803) );
  XNOR2X1 U274 ( .A(n885), .B(A[7]), .Y(n928) );
  XNOR2X1 U275 ( .A(n1132), .B(A[3]), .Y(n966) );
  OAI22XL U276 ( .A0(n926), .A1(n925), .B0(n924), .B1(n1085), .Y(n981) );
  NAND2BXL U277 ( .AN(A[0]), .B(n968), .Y(n927) );
  XNOR2XL U278 ( .A(n911), .B(A[7]), .Y(n322) );
  XOR2XL U279 ( .A(n885), .B(n43), .Y(n42) );
  INVXL U280 ( .A(A[4]), .Y(n43) );
  XNOR2XL U281 ( .A(n913), .B(A[10]), .Y(n285) );
  OAI22XL U282 ( .A0(n926), .A1(n199), .B0(n288), .B1(n1085), .Y(n271) );
  OAI22XL U283 ( .A0(n1125), .A1(n356), .B0(n5), .B1(n197), .Y(n270) );
  NAND2BXL U284 ( .AN(A[0]), .B(n1108), .Y(n197) );
  XNOR2XL U285 ( .A(n911), .B(A[23]), .Y(n429) );
  XNOR2XL U286 ( .A(n913), .B(A[25]), .Y(n454) );
  XNOR2X1 U287 ( .A(n1132), .B(A[15]), .Y(n470) );
  XNOR2X1 U288 ( .A(n1132), .B(A[14]), .Y(n506) );
  XNOR2XL U289 ( .A(n911), .B(A[19]), .Y(n564) );
  XNOR2XL U290 ( .A(n765), .B(A[25]), .Y(n503) );
  OAI22X1 U291 ( .A0(n935), .A1(n573), .B0(n933), .B1(n503), .Y(n562) );
  XNOR2XL U292 ( .A(n911), .B(A[20]), .Y(n508) );
  XNOR2X1 U293 ( .A(n1132), .B(A[13]), .Y(n544) );
  NAND2BXL U294 ( .AN(A[0]), .B(n913), .Y(n73) );
  XNOR2XL U295 ( .A(n882), .B(A[6]), .Y(n64) );
  XNOR2XL U296 ( .A(n882), .B(A[5]), .Y(n71) );
  XNOR2XL U297 ( .A(n913), .B(A[2]), .Y(n69) );
  XNOR2X1 U298 ( .A(n1054), .B(n1053), .Y(PRODUCT[17]) );
  NAND2XL U299 ( .A(n1234), .B(n1238), .Y(n1241) );
  NAND2XL U300 ( .A(n1199), .B(n1204), .Y(n1207) );
  INVXL U301 ( .A(n1236), .Y(n1203) );
  INVXL U302 ( .A(n1250), .Y(n1208) );
  NOR2XL U303 ( .A(n385), .B(n389), .Y(n393) );
  OAI2BB1XL U304 ( .A0N(n977), .A1N(n979), .B0(n360), .Y(n366) );
  INVXL U305 ( .A(n359), .Y(n360) );
  OAI22X1 U306 ( .A0(n836), .A1(n797), .B0(n835), .B1(n752), .Y(n802) );
  OAI22X2 U307 ( .A0(n1146), .A1(n798), .B0(n1147), .B1(n753), .Y(n801) );
  OAI22XL U308 ( .A0(n939), .A1(n849), .B0(n915), .B1(n809), .Y(n850) );
  OAI22X1 U309 ( .A0(n931), .A1(n847), .B0(n929), .B1(n807), .Y(n852) );
  OAI22XL U310 ( .A0(n939), .A1(n914), .B0(n915), .B1(n849), .Y(n891) );
  OAI22XL U311 ( .A0(n935), .A1(n889), .B0(n933), .B1(n848), .Y(n892) );
  OAI22X1 U312 ( .A0(n931), .A1(n886), .B0(n929), .B1(n847), .Y(n893) );
  OAI22X1 U313 ( .A0(n1146), .A1(n874), .B0(n1147), .B1(n837), .Y(n877) );
  OAI22X1 U314 ( .A0(n1146), .A1(n887), .B0(n1147), .B1(n874), .Y(n918) );
  INVX1 U315 ( .A(B[10]), .Y(n51) );
  INVXL U316 ( .A(n404), .Y(n405) );
  NOR2BXL U317 ( .AN(A[0]), .B(n122), .Y(n137) );
  NAND3X1 U318 ( .A(n241), .B(n240), .C(n52), .Y(n242) );
  NAND2XL U319 ( .A(n239), .B(n238), .Y(n52) );
  INVXL U320 ( .A(n1136), .Y(n1119) );
  OAI22XL U321 ( .A0(n1146), .A1(n1106), .B0(n1147), .B1(n1118), .Y(n1121) );
  OAI22XL U322 ( .A0(n1125), .A1(n375), .B0(n5), .B1(n1109), .Y(n1112) );
  OAI22XL U323 ( .A0(n1146), .A1(n376), .B0(n1147), .B1(n1106), .Y(n1111) );
  NAND2XL U324 ( .A(n27), .B(n810), .Y(n26) );
  NAND2BXL U325 ( .AN(n811), .B(n28), .Y(n27) );
  OAI22XL U326 ( .A0(n935), .A1(n95), .B0(n890), .B1(n94), .Y(n96) );
  NAND2BXL U327 ( .AN(A[0]), .B(n765), .Y(n94) );
  OAI22XL U328 ( .A0(n926), .A1(n99), .B0(n98), .B1(n1085), .Y(n112) );
  OAI22XL U329 ( .A0(n282), .A1(n100), .B0(n933), .B1(n81), .Y(n110) );
  CMPR32X1 U330 ( .A(n80), .B(n22), .C(n78), .CO(n118), .S(n117) );
  OAI22XL U331 ( .A0(n282), .A1(n81), .B0(n933), .B1(n70), .Y(n80) );
  BUFX1 U332 ( .A(n79), .Y(n22) );
  INVXL U333 ( .A(n1218), .Y(n1213) );
  NOR2X1 U334 ( .A(n243), .B(n242), .Y(n1070) );
  NOR2X1 U335 ( .A(n1075), .B(n1080), .Y(n59) );
  OAI21X1 U336 ( .A0(n1075), .A1(n1081), .B0(n1076), .Y(n55) );
  INVXL U337 ( .A(n1144), .Y(n1145) );
  INVXL U338 ( .A(n1150), .Y(n1140) );
  NOR2XL U339 ( .A(n97), .B(n96), .Y(n1223) );
  NAND2XL U340 ( .A(n97), .B(n96), .Y(n1224) );
  AOI21XL U341 ( .A0(n1212), .A1(n1213), .B0(n90), .Y(n1226) );
  INVXL U342 ( .A(n1211), .Y(n90) );
  INVXL U343 ( .A(n1187), .Y(n1196) );
  INVXL U344 ( .A(n144), .Y(n1177) );
  NOR2XL U345 ( .A(n155), .B(n154), .Y(n144) );
  NAND2X1 U346 ( .A(n195), .B(n194), .Y(n1081) );
  NOR2X1 U347 ( .A(n195), .B(n194), .Y(n1080) );
  INVXL U348 ( .A(n1234), .Y(n1162) );
  NAND2XL U349 ( .A(n1199), .B(n1168), .Y(n1170) );
  AOI21XL U350 ( .A0(n1205), .A1(n1168), .B0(n1167), .Y(n1169) );
  INVXL U351 ( .A(n1257), .Y(n1167) );
  INVXL U352 ( .A(n1254), .Y(n1171) );
  XNOR2XL U353 ( .A(n882), .B(A[22]), .Y(n727) );
  XNOR2XL U354 ( .A(n882), .B(A[17]), .Y(n924) );
  XNOR2XL U355 ( .A(n882), .B(A[15]), .Y(n338) );
  XNOR2XL U356 ( .A(n882), .B(A[16]), .Y(n925) );
  XNOR2XL U357 ( .A(n882), .B(A[12]), .Y(n199) );
  XNOR2XL U358 ( .A(n885), .B(A[14]), .Y(n653) );
  XNOR2XL U359 ( .A(n888), .B(A[22]), .Y(n655) );
  XNOR2XL U360 ( .A(n913), .B(A[20]), .Y(n656) );
  NAND2BXL U361 ( .AN(A[0]), .B(n911), .Y(n130) );
  XNOR2XL U362 ( .A(n882), .B(A[9]), .Y(n161) );
  NOR2XL U363 ( .A(n1242), .B(n1262), .Y(n38) );
  INVXL U364 ( .A(n1267), .Y(n488) );
  AOI21XL U365 ( .A0(n709), .A1(n641), .B0(n640), .Y(n642) );
  INVXL U366 ( .A(n1272), .Y(n644) );
  INVXL U367 ( .A(n1279), .Y(n708) );
  INVXL U368 ( .A(n1276), .Y(n712) );
  INVXL U369 ( .A(n1283), .Y(n787) );
  INVXL U370 ( .A(n1280), .Y(n791) );
  INVXL U371 ( .A(n1295), .Y(n1034) );
  AND2X2 U372 ( .A(n386), .B(n387), .Y(n39) );
  NAND2XL U373 ( .A(n637), .B(n387), .Y(n389) );
  NAND2XL U374 ( .A(n1168), .B(n1257), .Y(n1165) );
  INVXL U375 ( .A(n885), .Y(n159) );
  XNOR2XL U376 ( .A(n911), .B(A[16]), .Y(n682) );
  NOR2X1 U377 ( .A(n1143), .B(n616), .Y(n683) );
  ADDFX2 U378 ( .A(n692), .B(n691), .CI(n690), .CO(n701), .S(n742) );
  OAI22XL U379 ( .A0(n935), .A1(n688), .B0(n933), .B1(n655), .Y(n691) );
  OAI22XL U380 ( .A0(n939), .A1(n689), .B0(n915), .B1(n656), .Y(n690) );
  OAI22X1 U381 ( .A0(n49), .A1(n687), .B0(n929), .B1(n653), .Y(n692) );
  XNOR2XL U382 ( .A(n911), .B(A[14]), .Y(n758) );
  XNOR2XL U383 ( .A(n765), .B(A[19]), .Y(n766) );
  XNOR2XL U384 ( .A(n913), .B(A[16]), .Y(n809) );
  XNOR2X1 U385 ( .A(n885), .B(A[9]), .Y(n847) );
  XNOR2XL U386 ( .A(n888), .B(A[17]), .Y(n848) );
  XNOR2XL U387 ( .A(n913), .B(A[15]), .Y(n849) );
  XNOR2X1 U388 ( .A(n920), .B(A[15]), .Y(n797) );
  XNOR2XL U389 ( .A(n833), .B(A[14]), .Y(n834) );
  XNOR2XL U390 ( .A(n1108), .B(A[8]), .Y(n838) );
  XNOR2XL U391 ( .A(n833), .B(A[13]), .Y(n873) );
  XNOR2XL U392 ( .A(n1108), .B(A[7]), .Y(n875) );
  XNOR2XL U393 ( .A(n1108), .B(A[6]), .Y(n916) );
  XNOR2XL U394 ( .A(n913), .B(A[14]), .Y(n914) );
  XNOR2XL U395 ( .A(n913), .B(A[13]), .Y(n936) );
  XNOR2XL U396 ( .A(n1108), .B(A[5]), .Y(n970) );
  XNOR2XL U397 ( .A(n911), .B(A[9]), .Y(n976) );
  ADDFX2 U398 ( .A(n993), .B(n992), .CI(n991), .CO(n1005), .S(n1023) );
  OAI22X1 U399 ( .A0(n935), .A1(n934), .B0(n933), .B1(n932), .Y(n992) );
  OAI22XL U400 ( .A0(n939), .A1(n938), .B0(n937), .B1(n936), .Y(n991) );
  OAI22X1 U401 ( .A0(n931), .A1(n930), .B0(n929), .B1(n928), .Y(n993) );
  XNOR2X1 U402 ( .A(n765), .B(A[14]), .Y(n934) );
  XNOR2XL U403 ( .A(n1108), .B(A[4]), .Y(n971) );
  XNOR2XL U404 ( .A(n911), .B(A[8]), .Y(n978) );
  XNOR2XL U405 ( .A(n913), .B(A[12]), .Y(n938) );
  XNOR2X1 U406 ( .A(n885), .B(A[6]), .Y(n930) );
  XNOR2XL U407 ( .A(n913), .B(A[11]), .Y(n326) );
  CMPR22X1 U408 ( .A(n336), .B(n335), .CO(n1022), .S(n333) );
  OAI22X1 U409 ( .A0(n926), .A1(n287), .B0(n338), .B1(n1085), .Y(n336) );
  OAI22X1 U410 ( .A0(n1146), .A1(n354), .B0(n1147), .B1(n286), .Y(n335) );
  NAND2BXL U411 ( .AN(A[0]), .B(n1132), .Y(n286) );
  OAI22XL U412 ( .A0(n926), .A1(n288), .B0(n287), .B1(n1085), .Y(n292) );
  NOR2BXL U413 ( .AN(A[0]), .B(n266), .Y(n293) );
  OAI22XL U414 ( .A0(n1125), .A1(n290), .B0(n5), .B1(n289), .Y(n291) );
  CMPR32X1 U415 ( .A(n296), .B(n295), .C(n294), .CO(n301), .S(n304) );
  OAI22XL U416 ( .A0(n939), .A1(n218), .B0(n937), .B1(n268), .Y(n294) );
  OAI22XL U417 ( .A0(n979), .A1(n219), .B0(n977), .B1(n260), .Y(n296) );
  OAI22XL U418 ( .A0(n282), .A1(n217), .B0(n933), .B1(n262), .Y(n295) );
  OAI22XL U419 ( .A0(n975), .A1(n168), .B0(n835), .B1(n202), .Y(n207) );
  OAI22XL U420 ( .A0(n939), .A1(n204), .B0(n937), .B1(n218), .Y(n211) );
  OAI22XL U421 ( .A0(n282), .A1(n203), .B0(n933), .B1(n217), .Y(n212) );
  OAI22X1 U422 ( .A0(n1125), .A1(n215), .B0(n5), .B1(n290), .Y(n273) );
  OAI22XL U423 ( .A0(n975), .A1(n269), .B0(n835), .B1(n284), .Y(n276) );
  OAI22XL U424 ( .A0(n282), .A1(n262), .B0(n933), .B1(n281), .Y(n297) );
  OAI22X1 U425 ( .A0(n261), .A1(n931), .B0(n929), .B1(n42), .Y(n298) );
  OAI22X1 U426 ( .A0(n1146), .A1(n267), .B0(n1147), .B1(n339), .Y(n341) );
  XNOR2XL U427 ( .A(n1108), .B(A[18]), .Y(n466) );
  XNOR2XL U428 ( .A(n885), .B(A[19]), .Y(n471) );
  NOR2X1 U429 ( .A(n1143), .B(n468), .Y(n512) );
  OAI22XL U430 ( .A0(n1125), .A1(n509), .B0(n5), .B1(n467), .Y(n513) );
  CMPR32X1 U431 ( .A(n659), .B(n658), .C(n657), .CO(n665), .S(n700) );
  OAI22XL U432 ( .A0(n939), .A1(n656), .B0(n915), .B1(n608), .Y(n657) );
  OAI22X1 U433 ( .A0(n935), .A1(n655), .B0(n933), .B1(n607), .Y(n658) );
  OAI22XL U434 ( .A0(n654), .A1(n653), .B0(n929), .B1(n606), .Y(n659) );
  OAI22XL U435 ( .A0(n836), .A1(n542), .B0(n835), .B1(n507), .Y(n545) );
  OAI22X1 U436 ( .A0(n1146), .A1(n544), .B0(n1147), .B1(n506), .Y(n546) );
  OAI22XL U437 ( .A0(n979), .A1(n564), .B0(n977), .B1(n508), .Y(n550) );
  OAI22XL U438 ( .A0(n1125), .A1(n559), .B0(n5), .B1(n509), .Y(n549) );
  XNOR2XL U439 ( .A(n882), .B(A[8]), .Y(n131) );
  XNOR2XL U440 ( .A(n913), .B(A[6]), .Y(n165) );
  XNOR2XL U441 ( .A(n833), .B(A[4]), .Y(n168) );
  XNOR2XL U442 ( .A(n765), .B(A[8]), .Y(n170) );
  XNOR2XL U443 ( .A(n913), .B(A[5]), .Y(n166) );
  XNOR2XL U444 ( .A(n913), .B(A[4]), .Y(n125) );
  XNOR2XL U445 ( .A(n833), .B(A[2]), .Y(n133) );
  XNOR2XL U446 ( .A(n833), .B(A[3]), .Y(n164) );
  XNOR2XL U447 ( .A(n911), .B(A[1]), .Y(n163) );
  NAND2XL U448 ( .A(n1157), .B(n1259), .Y(n399) );
  OAI21XL U449 ( .A0(n1246), .A1(n398), .B0(n397), .Y(n400) );
  XNOR2X2 U450 ( .A(n452), .B(n451), .Y(PRODUCT[33]) );
  XNOR2X1 U451 ( .A(n646), .B(n645), .Y(PRODUCT[28]) );
  NAND2XL U452 ( .A(n644), .B(n1273), .Y(n645) );
  OAI21XL U453 ( .A0(n643), .A1(n1089), .B0(n642), .Y(n646) );
  OAI21XL U454 ( .A0(n1089), .A1(n385), .B0(n390), .Y(n353) );
  XNOR2X1 U455 ( .A(n829), .B(n828), .Y(PRODUCT[23]) );
  NAND2XL U456 ( .A(n788), .B(n1283), .Y(n828) );
  OAI21XL U457 ( .A0(n1089), .A1(n827), .B0(n826), .Y(n829) );
  XOR2X1 U458 ( .A(n1013), .B(n1012), .Y(PRODUCT[19]) );
  AOI21XL U459 ( .A0(n1239), .A1(n1238), .B0(n1237), .Y(n1240) );
  NAND2XL U460 ( .A(n1201), .B(n1253), .Y(n1185) );
  XNOR2XL U461 ( .A(n1108), .B(A[24]), .Y(n1109) );
  CMPR32X1 U462 ( .A(n611), .B(n610), .C(n609), .CO(n652), .S(n664) );
  OAI2BB1XL U463 ( .A0N(n761), .A1N(n845), .B0(n574), .Y(n609) );
  OAI22X1 U464 ( .A0(n836), .A1(n677), .B0(n835), .B1(n620), .Y(n681) );
  OAI22X1 U465 ( .A0(n836), .A1(n718), .B0(n835), .B1(n677), .Y(n723) );
  OAI22XL U466 ( .A0(n939), .A1(n731), .B0(n915), .B1(n689), .Y(n732) );
  OAI22X1 U467 ( .A0(n931), .A1(n729), .B0(n929), .B1(n687), .Y(n734) );
  OAI22X1 U468 ( .A0(n836), .A1(n752), .B0(n835), .B1(n718), .Y(n757) );
  OAI22X1 U469 ( .A0(n1146), .A1(n753), .B0(n1147), .B1(n719), .Y(n756) );
  NOR2X1 U470 ( .A(n34), .B(n33), .Y(n812) );
  CMPR32X1 U471 ( .A(n945), .B(n944), .C(n943), .CO(n946), .S(n1003) );
  OAI22XL U472 ( .A0(n935), .A1(n932), .B0(n890), .B1(n889), .Y(n982) );
  OAI22X1 U473 ( .A0(n931), .A1(n928), .B0(n929), .B1(n886), .Y(n984) );
  OAI22X1 U474 ( .A0(n1146), .A1(n966), .B0(n1147), .B1(n887), .Y(n983) );
  OAI22XL U475 ( .A0(n975), .A1(n284), .B0(n973), .B1(n328), .Y(n319) );
  OAI22XL U476 ( .A0(n282), .A1(n281), .B0(n933), .B1(n324), .Y(n321) );
  OAI22X1 U477 ( .A0(n929), .A1(n327), .B0(n931), .B1(n42), .Y(n320) );
  OAI22XL U478 ( .A0(n979), .A1(n429), .B0(n977), .B1(n409), .Y(n435) );
  OAI22XL U479 ( .A0(n1125), .A1(n428), .B0(n5), .B1(n411), .Y(n433) );
  INVXL U480 ( .A(n367), .Y(n412) );
  OAI22XL U481 ( .A0(n1146), .A1(n410), .B0(n1147), .B1(n364), .Y(n414) );
  OAI2BB1XL U482 ( .A0N(n915), .A1N(n595), .B0(n455), .Y(n472) );
  INVXL U483 ( .A(n454), .Y(n455) );
  OAI22XL U484 ( .A0(n979), .A1(n500), .B0(n977), .B1(n464), .Y(n475) );
  OAI22XL U485 ( .A0(n836), .A1(n469), .B0(n835), .B1(n462), .Y(n477) );
  OAI22XL U486 ( .A0(n1146), .A1(n470), .B0(n1147), .B1(n463), .Y(n476) );
  OR2XL U487 ( .A(n605), .B(n604), .Y(n578) );
  INVXL U488 ( .A(n562), .Y(n575) );
  OAI2BB1XL U489 ( .A0N(n933), .A1N(n935), .B0(n504), .Y(n561) );
  INVXL U490 ( .A(n503), .Y(n504) );
  ADDFX2 U491 ( .A(n600), .B(n599), .CI(n598), .CO(n583), .S(n618) );
  OAI22XL U492 ( .A0(n836), .A1(n567), .B0(n835), .B1(n542), .Y(n600) );
  ADDFX2 U493 ( .A(n665), .B(n664), .CI(n663), .CO(n671), .S(n703) );
  ADDFX2 U494 ( .A(n583), .B(n582), .CI(n581), .CO(n570), .S(n630) );
  XNOR2XL U495 ( .A(n882), .B(A[2]), .Y(n91) );
  XNOR2XL U496 ( .A(n765), .B(A[1]), .Y(n101) );
  XNOR2XL U497 ( .A(n882), .B(A[3]), .Y(n99) );
  XNOR2XL U498 ( .A(n913), .B(A[1]), .Y(n82) );
  XNOR2XL U499 ( .A(n765), .B(A[2]), .Y(n100) );
  XNOR2XL U500 ( .A(n765), .B(A[3]), .Y(n81) );
  OAI22XL U501 ( .A0(n926), .A1(n98), .B0(n71), .B1(n1085), .Y(n85) );
  INVXL U502 ( .A(n913), .Y(n74) );
  NAND2BXL U503 ( .AN(A[0]), .B(n833), .Y(n63) );
  ADDFX2 U504 ( .A(n140), .B(n139), .CI(n138), .CO(n146), .S(n148) );
  OAI22XL U505 ( .A0(n282), .A1(n70), .B0(n933), .B1(n124), .Y(n140) );
  OAI22X1 U506 ( .A0(n975), .A1(n68), .B0(n835), .B1(n134), .Y(n139) );
  OAI22XL U507 ( .A0(n282), .A1(n129), .B0(n933), .B1(n167), .Y(n184) );
  AND2X2 U508 ( .A(n1175), .B(n1177), .Y(n57) );
  NAND2XL U509 ( .A(n1208), .B(n1251), .Y(n1209) );
  NOR2BXL U510 ( .AN(A[0]), .B(n933), .Y(n88) );
  OAI22XL U511 ( .A0(n926), .A1(n86), .B0(n91), .B1(n1085), .Y(n89) );
  INVXL U512 ( .A(n373), .Y(n374) );
  OAI22XL U513 ( .A0(n1125), .A1(n411), .B0(n5), .B1(n401), .Y(n417) );
  INVXL U514 ( .A(n1104), .Y(n377) );
  OAI22XL U515 ( .A0(n1146), .A1(n361), .B0(n1147), .B1(n376), .Y(n379) );
  OAI22XL U516 ( .A0(n1125), .A1(n362), .B0(n5), .B1(n375), .Y(n382) );
  ADDFX2 U517 ( .A(n480), .B(n479), .CI(n478), .CO(n482), .S(n520) );
  XNOR2XL U518 ( .A(n882), .B(A[1]), .Y(n86) );
  INVX4 U519 ( .A(n61), .Y(n882) );
  INVX1 U520 ( .A(B[1]), .Y(n61) );
  BUFX3 U521 ( .A(n845), .Y(n926) );
  NAND2XL U522 ( .A(n89), .B(n88), .Y(n1211) );
  INVX1 U523 ( .A(n315), .Y(n41) );
  XNOR3X2 U524 ( .A(n46), .B(n588), .C(n587), .Y(n590) );
  OAI22XL U525 ( .A0(n1146), .A1(n1118), .B0(n1147), .B1(n1133), .Y(n1130) );
  ADDFX2 U526 ( .A(n1102), .B(n1101), .CI(n1100), .CO(n1114), .S(n383) );
  NAND2X1 U527 ( .A(n24), .B(n23), .Y(n795) );
  NAND2XL U528 ( .A(n822), .B(n823), .Y(n23) );
  OAI21XL U529 ( .A0(n822), .A1(n823), .B0(n821), .Y(n24) );
  NAND2X1 U530 ( .A(n32), .B(n31), .Y(n871) );
  NAND2X1 U531 ( .A(n905), .B(n904), .Y(n31) );
  XOR3X2 U532 ( .A(n905), .B(n904), .C(n903), .Y(n908) );
  NOR2X1 U533 ( .A(n350), .B(n349), .Y(n1092) );
  NAND2XL U534 ( .A(n350), .B(n349), .Y(n1063) );
  OAI21XL U535 ( .A0(n46), .A1(n45), .B0(n44), .Y(n554) );
  OAI21XL U536 ( .A0(n588), .A1(n589), .B0(n587), .Y(n44) );
  OAI22XL U537 ( .A0(n926), .A1(A[0]), .B0(n86), .B1(n1085), .Y(n1216) );
  NAND2XL U538 ( .A(n87), .B(n926), .Y(n1215) );
  NAND2BXL U539 ( .AN(A[0]), .B(n882), .Y(n87) );
  NAND2XL U540 ( .A(n1216), .B(n1215), .Y(n1218) );
  OAI21XL U541 ( .A0(mult_x_1_n308), .A1(n1067), .B0(n1068), .Y(mult_x_1_n301)
         );
  XNOR2XL U542 ( .A(n1214), .B(n1213), .Y(n1329) );
  NAND2XL U543 ( .A(n1212), .B(n1211), .Y(n1214) );
  INVXL U544 ( .A(n1095), .Y(n1099) );
  NAND2XL U545 ( .A(n1154), .B(n1153), .Y(mult_x_1_n58) );
  NAND2XL U546 ( .A(n1152), .B(n1151), .Y(n1153) );
  NOR2XL U547 ( .A(n1138), .B(n1137), .Y(mult_x_1_n109) );
  NAND2XL U548 ( .A(n1138), .B(n1137), .Y(mult_x_1_n110) );
  NOR2XL U549 ( .A(n1127), .B(n1126), .Y(mult_x_1_n120) );
  NAND2XL U550 ( .A(n1127), .B(n1126), .Y(mult_x_1_n121) );
  NOR2XL U551 ( .A(n1114), .B(n1113), .Y(mult_x_1_n129) );
  NAND2XL U552 ( .A(n1114), .B(n1113), .Y(mult_x_1_n130) );
  NAND2XL U553 ( .A(n636), .B(n635), .Y(mult_x_1_n198) );
  NOR2X1 U554 ( .A(n673), .B(n672), .Y(mult_x_1_n206) );
  NAND2XL U555 ( .A(n673), .B(n672), .Y(mult_x_1_n207) );
  NOR2XL U556 ( .A(n955), .B(n956), .Y(mult_x_1_n265) );
  NOR2XL U557 ( .A(n636), .B(n635), .Y(mult_x_1_n197) );
  NOR2BXL U558 ( .AN(A[0]), .B(n1085), .Y(n1331) );
  NAND2XL U559 ( .A(n1225), .B(n1224), .Y(n1227) );
  INVXL U560 ( .A(n1223), .Y(n1225) );
  NAND2XL U561 ( .A(n1220), .B(n1219), .Y(n1222) );
  NAND2XL U562 ( .A(n1230), .B(n1229), .Y(n1232) );
  INVXL U563 ( .A(n1228), .Y(n1230) );
  NAND2XL U564 ( .A(n1195), .B(n1194), .Y(n1197) );
  NAND2XL U565 ( .A(n1190), .B(n1189), .Y(n1191) );
  NAND2XL U566 ( .A(n1177), .B(n1176), .Y(n1178) );
  XOR2X1 U567 ( .A(n1084), .B(n1083), .Y(n1321) );
  OAI21X1 U568 ( .A0(n1284), .A1(n1287), .B0(n1285), .Y(n786) );
  AND2X1 U569 ( .A(n1155), .B(n1261), .Y(n21) );
  NOR2X1 U570 ( .A(n337), .B(n884), .Y(n922) );
  AOI21X1 U571 ( .A0(n393), .A1(n392), .B0(n391), .Y(n394) );
  AOI21X1 U572 ( .A0(n1054), .A1(n959), .B0(n958), .Y(n1013) );
  OAI21X2 U573 ( .A0(n157), .A1(n1174), .B0(n56), .Y(n1074) );
  OAI22X1 U574 ( .A0(n595), .A1(n74), .B0(n915), .B1(n73), .Y(n84) );
  NOR2X1 U575 ( .A(n1188), .B(n1193), .Y(n121) );
  OAI22X1 U576 ( .A0(n979), .A1(n842), .B0(n977), .B1(n803), .Y(n814) );
  OAI22X1 U577 ( .A0(n979), .A1(n912), .B0(n977), .B1(n879), .Y(n896) );
  CMPR22X1 U578 ( .A(n103), .B(n102), .CO(n105), .S(n97) );
  XNOR2X1 U579 ( .A(n34), .B(n843), .Y(n854) );
  OAI22X1 U580 ( .A0(n836), .A1(n462), .B0(n835), .B1(n404), .Y(n437) );
  CMPR22X1 U581 ( .A(n614), .B(n613), .CO(n627), .S(n661) );
  OAI22X1 U582 ( .A0(n979), .A1(n879), .B0(n977), .B1(n842), .Y(n855) );
  OAI22X1 U583 ( .A0(n979), .A1(n803), .B0(n977), .B1(n758), .Y(n773) );
  CMPR22X1 U584 ( .A(n128), .B(n127), .CO(n141), .S(n150) );
  OAI22X1 U585 ( .A0(n836), .A1(n283), .B0(n835), .B1(n63), .Y(n127) );
  CMPR22X1 U586 ( .A(n221), .B(n220), .CO(n226), .S(n208) );
  OAI22X1 U587 ( .A0(n654), .A1(n159), .B0(n929), .B1(n158), .Y(n220) );
  OAI22X1 U588 ( .A0(n979), .A1(n409), .B0(n977), .B1(n359), .Y(n367) );
  OAI22X1 U589 ( .A0(n935), .A1(n808), .B0(n933), .B1(n766), .Y(n811) );
  NOR2X2 U590 ( .A(n120), .B(n58), .Y(n1174) );
  XNOR2X1 U591 ( .A(n1132), .B(A[4]), .Y(n887) );
  XOR2X1 U592 ( .A(n1089), .B(n1088), .Y(PRODUCT[21]) );
  XNOR2X2 U593 ( .A(n869), .B(n868), .Y(PRODUCT[22]) );
  ADDFX2 U594 ( .A(n277), .B(n276), .CI(n275), .CO(n343), .S(n307) );
  CMPR22X1 U595 ( .A(n923), .B(n922), .CO(n894), .S(n944) );
  OAI22X1 U596 ( .A0(n939), .A1(n809), .B0(n915), .B1(n767), .Y(n810) );
  XNOR2X1 U597 ( .A(n48), .B(n804), .Y(n813) );
  XOR2X1 U598 ( .A(n1073), .B(n1072), .Y(n1318) );
  NAND2X1 U599 ( .A(n866), .B(n865), .Y(mult_x_1_n252) );
  XOR3X2 U600 ( .A(n823), .B(n821), .C(n822), .Y(n830) );
  NAND2X4 U601 ( .A(n198), .B(n25), .Y(n1125) );
  XOR2X1 U602 ( .A(B[12]), .B(B[13]), .Y(n25) );
  NAND2XL U603 ( .A(n956), .B(n955), .Y(mult_x_1_n266) );
  XOR2X1 U604 ( .A(n29), .B(n810), .Y(n860) );
  XOR2X1 U605 ( .A(n811), .B(n30), .Y(n29) );
  OAI22X4 U606 ( .A0(n931), .A1(n807), .B0(n764), .B1(n929), .Y(n30) );
  NOR2X1 U607 ( .A(n38), .B(n37), .Y(n424) );
  NAND2BX2 U608 ( .AN(n316), .B(n41), .Y(n1091) );
  NAND2X4 U609 ( .A(n50), .B(n566), .Y(n654) );
  XNOR2X4 U610 ( .A(B[9]), .B(B[10]), .Y(n566) );
  XNOR2X2 U611 ( .A(B[11]), .B(n51), .Y(n50) );
  NAND2XL U612 ( .A(n316), .B(n315), .Y(n1086) );
  OAI22X1 U613 ( .A0(n931), .A1(n327), .B0(n929), .B1(n930), .Y(n995) );
  OAI22X1 U614 ( .A0(n939), .A1(n326), .B0(n937), .B1(n938), .Y(n996) );
  AOI21X1 U615 ( .A0(n254), .A1(n786), .B0(n253), .Y(n390) );
  XNOR2X2 U616 ( .A(B[15]), .B(B[16]), .Y(n337) );
  CMPR22X1 U617 ( .A(n881), .B(n880), .CO(n853), .S(n895) );
  NOR2X2 U618 ( .A(n156), .B(n57), .Y(n56) );
  XNOR2X1 U619 ( .A(n1079), .B(n1078), .Y(n1320) );
  NAND2X1 U620 ( .A(n196), .B(n53), .Y(n1076) );
  NOR2X2 U621 ( .A(n196), .B(n53), .Y(n1075) );
  XOR2X2 U622 ( .A(n54), .B(n239), .Y(n53) );
  AOI21X2 U623 ( .A0(n59), .A1(n1074), .B0(n55), .Y(n1095) );
  AND2X2 U624 ( .A(n121), .B(n1187), .Y(n58) );
  NAND2X2 U625 ( .A(n122), .B(n60), .Y(n323) );
  XOR2X1 U626 ( .A(B[8]), .B(B[9]), .Y(n60) );
  XNOR2X2 U627 ( .A(B[13]), .B(B[14]), .Y(n266) );
  BUFX8 U628 ( .A(n654), .Y(n931) );
  XOR2X2 U629 ( .A(n1246), .B(n593), .Y(PRODUCT[29]) );
  CMPR22X1 U630 ( .A(n684), .B(n683), .CO(n660), .S(n694) );
  CMPR22X1 U631 ( .A(n726), .B(n725), .CO(n693), .S(n736) );
  OAI22XL U632 ( .A0(n654), .A1(n606), .B0(n929), .B1(n572), .Y(n611) );
  BUFX4 U633 ( .A(n67), .Y(n975) );
  OAI21XL U634 ( .A0(n390), .A1(n389), .B0(n388), .Y(n391) );
  INVX1 U635 ( .A(n911), .Y(n358) );
  XNOR2XL U636 ( .A(n882), .B(A[23]), .Y(n685) );
  XNOR2X1 U637 ( .A(n885), .B(A[15]), .Y(n606) );
  XNOR2X1 U638 ( .A(n920), .B(A[16]), .Y(n752) );
  XNOR2X1 U639 ( .A(n885), .B(A[16]), .Y(n572) );
  OAI22X1 U640 ( .A0(n1146), .A1(n506), .B0(n1147), .B1(n470), .Y(n515) );
  BUFX3 U641 ( .A(n890), .Y(n933) );
  ADDFX2 U642 ( .A(n541), .B(n540), .CI(n539), .CO(n537), .S(n571) );
  NAND2X1 U643 ( .A(B[1]), .B(n761), .Y(n845) );
  BUFX3 U644 ( .A(n761), .Y(n1085) );
  OAI22X1 U645 ( .A0(n926), .A1(n64), .B0(n132), .B1(n1085), .Y(n128) );
  XOR2X1 U646 ( .A(B[6]), .B(B[7]), .Y(n62) );
  XNOR2X4 U647 ( .A(B[6]), .B(B[5]), .Y(n973) );
  BUFX3 U648 ( .A(n67), .Y(n836) );
  INVX4 U649 ( .A(n833), .Y(n283) );
  NOR2BX1 U650 ( .AN(A[0]), .B(n835), .Y(n77) );
  OAI22X1 U651 ( .A0(n926), .A1(n71), .B0(n64), .B1(n1085), .Y(n76) );
  XOR2X1 U652 ( .A(B[4]), .B(B[5]), .Y(n65) );
  XNOR2X1 U653 ( .A(B[4]), .B(B[3]), .Y(n72) );
  BUFX3 U654 ( .A(n72), .Y(n937) );
  OAI22X1 U655 ( .A0(n939), .A1(n82), .B0(n937), .B1(n69), .Y(n75) );
  BUFX3 U656 ( .A(B[3]), .Y(n888) );
  INVX4 U657 ( .A(n888), .Y(n95) );
  INVX8 U658 ( .A(n95), .Y(n765) );
  XNOR2X1 U659 ( .A(n765), .B(A[5]), .Y(n124) );
  XNOR2XL U660 ( .A(n833), .B(A[0]), .Y(n68) );
  XNOR2XL U661 ( .A(n833), .B(A[1]), .Y(n134) );
  XNOR2XL U662 ( .A(n913), .B(A[3]), .Y(n126) );
  OAI22XL U663 ( .A0(n939), .A1(n69), .B0(n937), .B1(n126), .Y(n138) );
  BUFX3 U664 ( .A(n72), .Y(n915) );
  ADDFHX1 U665 ( .A(n77), .B(n76), .CI(n75), .CO(n149), .S(n78) );
  NOR2X1 U666 ( .A(n119), .B(n118), .Y(n1188) );
  XNOR2XL U667 ( .A(n913), .B(A[0]), .Y(n83) );
  OAI22XL U668 ( .A0(n939), .A1(n83), .B0(n937), .B1(n82), .Y(n109) );
  ADDHXL U669 ( .A(n85), .B(n84), .CO(n79), .S(n108) );
  OR2X2 U670 ( .A(n89), .B(n88), .Y(n1212) );
  OAI22X1 U671 ( .A0(n926), .A1(n91), .B0(n99), .B1(n1085), .Y(n103) );
  XNOR2X1 U672 ( .A(n765), .B(A[0]), .Y(n92) );
  OAI22X1 U673 ( .A0(n282), .A1(n92), .B0(n933), .B1(n101), .Y(n102) );
  BUFX3 U674 ( .A(n93), .Y(n935) );
  OAI21XL U675 ( .A0(n1226), .A1(n1223), .B0(n1224), .Y(n1221) );
  OAI22XL U676 ( .A0(n282), .A1(n101), .B0(n933), .B1(n100), .Y(n111) );
  NOR2XL U677 ( .A(n106), .B(n105), .Y(n104) );
  INVXL U678 ( .A(n104), .Y(n1220) );
  NAND2XL U679 ( .A(n106), .B(n105), .Y(n1219) );
  INVXL U680 ( .A(n1219), .Y(n107) );
  AOI21XL U681 ( .A0(n1221), .A1(n1220), .B0(n107), .Y(n1231) );
  CMPR32X1 U682 ( .A(n110), .B(n109), .C(n108), .CO(n116), .S(n115) );
  CMPR32X1 U683 ( .A(n113), .B(n112), .C(n111), .CO(n114), .S(n106) );
  NOR2XL U684 ( .A(n115), .B(n114), .Y(n1228) );
  NAND2XL U685 ( .A(n115), .B(n114), .Y(n1229) );
  OAI21XL U686 ( .A0(n1231), .A1(n1228), .B0(n1229), .Y(n1187) );
  NAND2XL U687 ( .A(n119), .B(n118), .Y(n1189) );
  OAI21XL U688 ( .A0(n1188), .A1(n1194), .B0(n1189), .Y(n120) );
  XNOR2XL U689 ( .A(n911), .B(A[0]), .Y(n123) );
  OAI22X1 U690 ( .A0(n979), .A1(n123), .B0(n977), .B1(n163), .Y(n177) );
  OAI22XL U691 ( .A0(n939), .A1(n125), .B0(n937), .B1(n166), .Y(n176) );
  XNOR2X1 U692 ( .A(n765), .B(A[6]), .Y(n129) );
  OAI22X1 U693 ( .A0(n282), .A1(n124), .B0(n933), .B1(n129), .Y(n143) );
  OAI22X2 U694 ( .A0(n939), .A1(n126), .B0(n937), .B1(n125), .Y(n142) );
  XNOR2X1 U695 ( .A(n765), .B(A[7]), .Y(n167) );
  OAI22X1 U696 ( .A0(n926), .A1(n131), .B0(n161), .B1(n1085), .Y(n172) );
  OAI22X4 U697 ( .A0(n979), .A1(n358), .B0(n977), .B1(n130), .Y(n171) );
  OAI22X1 U698 ( .A0(n926), .A1(n132), .B0(n131), .B1(n1085), .Y(n136) );
  OAI22XL U699 ( .A0(n975), .A1(n134), .B0(n835), .B1(n133), .Y(n135) );
  CMPR32X1 U700 ( .A(n137), .B(n136), .C(n135), .CO(n182), .S(n147) );
  ADDFHX1 U701 ( .A(n147), .B(n146), .CI(n145), .CO(n154), .S(n153) );
  CMPR32X1 U702 ( .A(n150), .B(n149), .C(n148), .CO(n152), .S(n119) );
  NAND2XL U703 ( .A(n155), .B(n154), .Y(n1176) );
  INVXL U704 ( .A(n1176), .Y(n156) );
  OAI22X1 U705 ( .A0(n926), .A1(n160), .B0(n200), .B1(n1085), .Y(n221) );
  BUFX8 U706 ( .A(B[11]), .Y(n885) );
  BUFX8 U707 ( .A(n566), .Y(n929) );
  OAI22X2 U708 ( .A0(n939), .A1(n166), .B0(n937), .B1(n165), .Y(n180) );
  XNOR2XL U709 ( .A(n833), .B(A[5]), .Y(n202) );
  XNOR2X1 U710 ( .A(n885), .B(A[0]), .Y(n169) );
  XNOR2X1 U711 ( .A(n885), .B(A[1]), .Y(n201) );
  XNOR2X1 U712 ( .A(n765), .B(A[9]), .Y(n203) );
  OAI22XL U713 ( .A0(n282), .A1(n170), .B0(n933), .B1(n203), .Y(n205) );
  CMPR22X1 U714 ( .A(n172), .B(n171), .CO(n187), .S(n183) );
  CMPR32X1 U715 ( .A(n184), .B(n183), .C(n182), .CO(n189), .S(n191) );
  CMPR32X1 U716 ( .A(n187), .B(n186), .C(n185), .CO(n239), .S(n188) );
  CMPR32X1 U717 ( .A(n190), .B(n189), .C(n188), .CO(n196), .S(n195) );
  INVX4 U718 ( .A(B[13]), .Y(n356) );
  INVX8 U719 ( .A(n356), .Y(n1108) );
  NOR2BX1 U720 ( .AN(A[0]), .B(n5), .Y(n224) );
  OAI22X2 U721 ( .A0(n926), .A1(n200), .B0(n199), .B1(n1085), .Y(n223) );
  XNOR2X1 U722 ( .A(n885), .B(A[2]), .Y(n216) );
  OAI22XL U723 ( .A0(n931), .A1(n201), .B0(n929), .B1(n216), .Y(n222) );
  XNOR2X1 U724 ( .A(n833), .B(A[6]), .Y(n214) );
  OAI22XL U725 ( .A0(n975), .A1(n202), .B0(n835), .B1(n214), .Y(n213) );
  XNOR2X1 U726 ( .A(n765), .B(A[10]), .Y(n217) );
  ADDFHX1 U727 ( .A(n207), .B(n206), .CI(n205), .CO(n233), .S(n228) );
  CMPR32X1 U728 ( .A(n213), .B(n212), .C(n211), .CO(n278), .S(n231) );
  XNOR2X1 U729 ( .A(n833), .B(A[7]), .Y(n269) );
  OAI22XL U730 ( .A0(n975), .A1(n214), .B0(n973), .B1(n269), .Y(n274) );
  XNOR2X1 U731 ( .A(n1108), .B(A[0]), .Y(n215) );
  XNOR2X1 U732 ( .A(n1108), .B(A[1]), .Y(n290) );
  XNOR2X1 U733 ( .A(n885), .B(A[3]), .Y(n261) );
  OAI22XL U734 ( .A0(n931), .A1(n216), .B0(n929), .B1(n261), .Y(n272) );
  XNOR2XL U735 ( .A(n911), .B(A[4]), .Y(n219) );
  XNOR2XL U736 ( .A(n911), .B(A[5]), .Y(n260) );
  XNOR2X1 U737 ( .A(n765), .B(A[11]), .Y(n262) );
  CMPR32X1 U738 ( .A(n227), .B(n226), .C(n225), .CO(n303), .S(n236) );
  ADDFHX1 U739 ( .A(n230), .B(n229), .CI(n228), .CO(n235), .S(n238) );
  CMPR32X1 U740 ( .A(n236), .B(n235), .C(n234), .CO(n244), .S(n243) );
  NAND2XL U741 ( .A(n239), .B(n237), .Y(n241) );
  NAND2XL U742 ( .A(n237), .B(n238), .Y(n240) );
  INVXL U743 ( .A(n1071), .Y(n246) );
  NOR2X4 U744 ( .A(n1288), .B(n1290), .Y(n250) );
  NAND2X2 U745 ( .A(n250), .B(n959), .Y(n252) );
  AOI21X4 U746 ( .A0(n1296), .A1(n1303), .B0(n1300), .Y(n957) );
  OAI21X2 U747 ( .A0(n1292), .A1(n1295), .B0(n1293), .Y(n958) );
  AOI21X4 U748 ( .A0(n250), .A1(n958), .B0(n249), .Y(n251) );
  OAI21X4 U749 ( .A0(n252), .A1(n957), .B0(n251), .Y(n392) );
  INVX4 U750 ( .A(n392), .Y(n1089) );
  NAND2XL U751 ( .A(n707), .B(n637), .Y(n256) );
  OAI21XL U752 ( .A0(n1280), .A1(n1283), .B0(n1281), .Y(n253) );
  INVXL U753 ( .A(n386), .Y(n639) );
  AOI21XL U754 ( .A0(n709), .A1(n637), .B0(n386), .Y(n255) );
  OAI22XL U755 ( .A0(n323), .A1(n260), .B0(n977), .B1(n263), .Y(n299) );
  XNOR2X1 U756 ( .A(n765), .B(A[12]), .Y(n281) );
  OAI22XL U757 ( .A0(n323), .A1(n263), .B0(n977), .B1(n322), .Y(n342) );
  XOR2X1 U758 ( .A(B[14]), .B(B[15]), .Y(n264) );
  INVX8 U759 ( .A(n354), .Y(n1132) );
  XNOR2XL U760 ( .A(n1132), .B(A[0]), .Y(n267) );
  XNOR2X1 U761 ( .A(n1132), .B(A[1]), .Y(n339) );
  XNOR2X1 U762 ( .A(n1108), .B(A[2]), .Y(n289) );
  XNOR2X1 U763 ( .A(n1108), .B(A[3]), .Y(n325) );
  OAI22XL U764 ( .A0(n1125), .A1(n289), .B0(n5), .B1(n325), .Y(n340) );
  OAI22XL U765 ( .A0(n939), .A1(n268), .B0(n937), .B1(n285), .Y(n277) );
  XNOR2X1 U766 ( .A(n833), .B(A[8]), .Y(n284) );
  ADDHXL U767 ( .A(n271), .B(n270), .CO(n275), .S(n280) );
  ADDFHX1 U768 ( .A(n274), .B(n273), .CI(n272), .CO(n308), .S(n305) );
  ADDFHX1 U769 ( .A(n280), .B(n279), .CI(n278), .CO(n306), .S(n314) );
  XNOR2X1 U770 ( .A(n885), .B(A[5]), .Y(n327) );
  INVX8 U771 ( .A(n283), .Y(n920) );
  XNOR2X1 U772 ( .A(n920), .B(A[9]), .Y(n328) );
  OAI22X1 U773 ( .A0(n939), .A1(n285), .B0(n937), .B1(n326), .Y(n334) );
  CMPR32X1 U774 ( .A(n293), .B(n292), .C(n291), .CO(n332), .S(n302) );
  CMPR32X1 U775 ( .A(n299), .B(n298), .C(n297), .CO(n345), .S(n300) );
  CMPR32X1 U776 ( .A(n305), .B(n304), .C(n303), .CO(n310), .S(n312) );
  ADDFHX1 U777 ( .A(n311), .B(n310), .CI(n309), .CO(n315), .S(n1066) );
  INVXL U778 ( .A(n1068), .Y(n318) );
  INVXL U779 ( .A(n1086), .Y(n317) );
  AOI21X2 U780 ( .A0(n1091), .A1(n318), .B0(n317), .Y(n1093) );
  CMPR32X1 U781 ( .A(n321), .B(n320), .C(n319), .CO(n1028), .S(n331) );
  OAI22XL U782 ( .A0(n323), .A1(n322), .B0(n977), .B1(n978), .Y(n990) );
  OAI22XL U783 ( .A0(n935), .A1(n324), .B0(n933), .B1(n934), .Y(n989) );
  OAI22XL U784 ( .A0(n1125), .A1(n325), .B0(n5), .B1(n971), .Y(n988) );
  XNOR2XL U785 ( .A(n920), .B(A[10]), .Y(n974) );
  OAI22XL U786 ( .A0(n975), .A1(n328), .B0(n973), .B1(n974), .Y(n994) );
  NOR2BX1 U787 ( .AN(A[0]), .B(n1143), .Y(n987) );
  OAI22X1 U788 ( .A0(n926), .A1(n338), .B0(n925), .B1(n761), .Y(n986) );
  XNOR2X1 U789 ( .A(n1132), .B(A[2]), .Y(n967) );
  OAI22XL U790 ( .A0(n1146), .A1(n339), .B0(n1147), .B1(n967), .Y(n985) );
  ADDFHX1 U791 ( .A(n342), .B(n341), .CI(n340), .CO(n1020), .S(n344) );
  CMPR32X1 U792 ( .A(n345), .B(n344), .C(n343), .CO(n1045), .S(n348) );
  CMPR32X1 U793 ( .A(n348), .B(n347), .C(n346), .CO(n349), .S(n316) );
  NAND2XL U794 ( .A(n351), .B(n1279), .Y(n352) );
  XNOR2X1 U795 ( .A(n1132), .B(A[20]), .Y(n361) );
  XNOR2X1 U796 ( .A(n1132), .B(A[21]), .Y(n376) );
  BUFX3 U797 ( .A(B[16]), .Y(n501) );
  XNOR2XL U798 ( .A(n501), .B(A[19]), .Y(n355) );
  XNOR2X1 U799 ( .A(n885), .B(A[24]), .Y(n363) );
  XNOR2XL U800 ( .A(n885), .B(A[25]), .Y(n373) );
  OAI22X1 U801 ( .A0(n654), .A1(n363), .B0(n566), .B1(n373), .Y(n1104) );
  XNOR2X1 U802 ( .A(n1108), .B(A[22]), .Y(n362) );
  XNOR2X1 U803 ( .A(n1108), .B(A[23]), .Y(n375) );
  XNOR2X1 U804 ( .A(n501), .B(A[18]), .Y(n357) );
  XNOR2XL U805 ( .A(n911), .B(A[24]), .Y(n409) );
  XNOR2XL U806 ( .A(n911), .B(A[25]), .Y(n359) );
  XNOR2X1 U807 ( .A(n1132), .B(A[19]), .Y(n364) );
  XNOR2X1 U808 ( .A(n1108), .B(A[21]), .Y(n401) );
  XNOR2X1 U809 ( .A(n885), .B(A[23]), .Y(n365) );
  XNOR2XL U810 ( .A(n1132), .B(A[18]), .Y(n410) );
  XNOR2X1 U811 ( .A(n885), .B(A[22]), .Y(n427) );
  OAI22XL U812 ( .A0(n654), .A1(n427), .B0(n566), .B1(n365), .Y(n413) );
  CMPR32X1 U813 ( .A(n368), .B(n367), .C(n366), .CO(n381), .S(n407) );
  CMPR32X1 U814 ( .A(n371), .B(n370), .C(n369), .CO(n380), .S(n406) );
  OAI2BB1X1 U815 ( .A0N(n566), .A1N(n654), .B0(n374), .Y(n1103) );
  XNOR2X1 U816 ( .A(n1132), .B(A[22]), .Y(n1106) );
  CMPR32X1 U817 ( .A(n379), .B(n378), .C(n377), .CO(n1110), .S(n420) );
  CMPR32X1 U818 ( .A(n382), .B(n381), .C(n380), .CO(n1100), .S(n419) );
  NOR2XL U819 ( .A(n384), .B(n383), .Y(mult_x_1_n136) );
  NAND2XL U820 ( .A(n384), .B(n383), .Y(mult_x_1_n137) );
  NOR2XL U821 ( .A(n1270), .B(n1268), .Y(n486) );
  NOR2XL U822 ( .A(n1266), .B(n1264), .Y(n396) );
  NOR2XL U823 ( .A(n1235), .B(n1262), .Y(n423) );
  NAND2XL U824 ( .A(n423), .B(n1155), .Y(n398) );
  OAI21XL U825 ( .A0(n1268), .A1(n1271), .B0(n1269), .Y(n487) );
  OAI21XL U826 ( .A0(n1264), .A1(n1267), .B0(n1265), .Y(n395) );
  XNOR2X1 U827 ( .A(n1108), .B(A[20]), .Y(n411) );
  XNOR2X1 U828 ( .A(n501), .B(A[16]), .Y(n403) );
  XNOR2X1 U829 ( .A(n920), .B(A[24]), .Y(n462) );
  XNOR2XL U830 ( .A(n920), .B(A[25]), .Y(n404) );
  CMPR32X1 U831 ( .A(n408), .B(n407), .C(n406), .CO(n418), .S(n446) );
  XNOR2X1 U832 ( .A(n1132), .B(A[17]), .Y(n431) );
  OAI22XL U833 ( .A0(n1146), .A1(n431), .B0(n1147), .B1(n410), .Y(n434) );
  XNOR2X1 U834 ( .A(n1108), .B(A[19]), .Y(n428) );
  CMPR32X1 U835 ( .A(n414), .B(n413), .C(n412), .CO(n408), .S(n443) );
  CMPR32X1 U836 ( .A(n417), .B(n416), .C(n415), .CO(n447), .S(n442) );
  CMPR32X1 U837 ( .A(n420), .B(n419), .C(n418), .CO(n384), .S(n421) );
  NOR2XL U838 ( .A(n422), .B(n421), .Y(mult_x_1_n151) );
  NAND2XL U839 ( .A(n422), .B(n421), .Y(mult_x_1_n152) );
  INVXL U840 ( .A(n423), .Y(n425) );
  OAI21XL U841 ( .A0(n1246), .A1(n425), .B0(n424), .Y(n426) );
  XNOR2X1 U842 ( .A(n885), .B(A[21]), .Y(n432) );
  OAI22XL U843 ( .A0(n1125), .A1(n466), .B0(n5), .B1(n428), .Y(n461) );
  XNOR2XL U844 ( .A(n911), .B(A[22]), .Y(n464) );
  OAI22XL U845 ( .A0(n979), .A1(n464), .B0(n977), .B1(n429), .Y(n460) );
  INVXL U846 ( .A(n437), .Y(n459) );
  XNOR2X1 U847 ( .A(n501), .B(A[15]), .Y(n430) );
  XNOR2X1 U848 ( .A(n1132), .B(A[16]), .Y(n463) );
  OAI22XL U849 ( .A0(n1146), .A1(n463), .B0(n1147), .B1(n431), .Y(n457) );
  XNOR2XL U850 ( .A(n885), .B(A[20]), .Y(n465) );
  OAI22XL U851 ( .A0(n654), .A1(n465), .B0(n566), .B1(n432), .Y(n456) );
  CMPR32X1 U852 ( .A(n435), .B(n434), .C(n433), .CO(n444), .S(n480) );
  CMPR32X1 U853 ( .A(n438), .B(n437), .C(n436), .CO(n415), .S(n479) );
  CMPR32X1 U854 ( .A(n444), .B(n443), .C(n442), .CO(n445), .S(n481) );
  CMPR32X1 U855 ( .A(n447), .B(n446), .C(n445), .CO(n422), .S(n448) );
  NOR2XL U856 ( .A(n449), .B(n448), .Y(mult_x_1_n160) );
  NAND2XL U857 ( .A(n449), .B(n448), .Y(mult_x_1_n161) );
  OAI21XL U858 ( .A0(n1246), .A1(n1235), .B0(n1242), .Y(n452) );
  XNOR2XL U859 ( .A(n501), .B(A[14]), .Y(n453) );
  XNOR2XL U860 ( .A(n913), .B(A[24]), .Y(n505) );
  OAI22X1 U861 ( .A0(n939), .A1(n505), .B0(n915), .B1(n454), .Y(n473) );
  CMPR32X1 U862 ( .A(n458), .B(n457), .C(n456), .CO(n439), .S(n495) );
  CMPR32X1 U863 ( .A(n461), .B(n460), .C(n459), .CO(n440), .S(n494) );
  XNOR2XL U864 ( .A(n911), .B(A[21]), .Y(n500) );
  OAI22XL U865 ( .A0(n654), .A1(n471), .B0(n566), .B1(n465), .Y(n499) );
  XNOR2X1 U866 ( .A(n1108), .B(A[17]), .Y(n467) );
  OAI22XL U867 ( .A0(n1125), .A1(n467), .B0(n5), .B1(n466), .Y(n498) );
  XNOR2X1 U868 ( .A(n501), .B(A[13]), .Y(n468) );
  INVXL U869 ( .A(n473), .Y(n511) );
  OAI22X1 U870 ( .A0(n836), .A1(n507), .B0(n835), .B1(n469), .Y(n516) );
  XNOR2X1 U871 ( .A(n885), .B(A[18]), .Y(n510) );
  OAI22XL U872 ( .A0(n654), .A1(n510), .B0(n566), .B1(n471), .Y(n514) );
  CMPR32X1 U873 ( .A(n474), .B(n473), .C(n472), .CO(n496), .S(n534) );
  CMPR32X1 U874 ( .A(n477), .B(n476), .C(n475), .CO(n519), .S(n533) );
  CMPR32X1 U875 ( .A(n483), .B(n482), .C(n481), .CO(n449), .S(n484) );
  NOR2XL U876 ( .A(n485), .B(n484), .Y(mult_x_1_n169) );
  NAND2XL U877 ( .A(n485), .B(n484), .Y(mult_x_1_n170) );
  INVXL U878 ( .A(n486), .Y(n526) );
  NAND2XL U879 ( .A(n486), .B(n527), .Y(n490) );
  INVXL U880 ( .A(n487), .Y(n525) );
  AOI21XL U881 ( .A0(n487), .A1(n527), .B0(n488), .Y(n489) );
  OAI21X1 U882 ( .A0(n1246), .A1(n490), .B0(n489), .Y(n493) );
  INVXL U883 ( .A(n1264), .Y(n491) );
  NAND2X1 U884 ( .A(n491), .B(n1265), .Y(n492) );
  XNOR2X2 U885 ( .A(n493), .B(n492), .Y(PRODUCT[32]) );
  CMPR32X1 U886 ( .A(n496), .B(n495), .C(n494), .CO(n522), .S(n532) );
  CMPR32X1 U887 ( .A(n499), .B(n498), .C(n497), .CO(n518), .S(n538) );
  OAI22XL U888 ( .A0(n979), .A1(n508), .B0(n977), .B1(n500), .Y(n541) );
  XNOR2XL U889 ( .A(n501), .B(A[12]), .Y(n502) );
  XNOR2X1 U890 ( .A(n765), .B(A[24]), .Y(n573) );
  XNOR2XL U891 ( .A(n913), .B(A[23]), .Y(n560) );
  OAI22XL U892 ( .A0(n595), .A1(n560), .B0(n915), .B1(n505), .Y(n547) );
  XNOR2X1 U893 ( .A(n920), .B(A[21]), .Y(n542) );
  XNOR2X1 U894 ( .A(n1108), .B(A[15]), .Y(n559) );
  XNOR2XL U895 ( .A(n885), .B(A[17]), .Y(n565) );
  OAI22XL U896 ( .A0(n654), .A1(n565), .B0(n566), .B1(n510), .Y(n548) );
  ADDFHX1 U897 ( .A(n513), .B(n512), .CI(n511), .CO(n497), .S(n552) );
  CMPR32X1 U898 ( .A(n519), .B(n518), .C(n517), .CO(n521), .S(n530) );
  CMPR32X1 U899 ( .A(n522), .B(n521), .C(n520), .CO(n485), .S(n523) );
  NOR2XL U900 ( .A(n524), .B(n523), .Y(mult_x_1_n176) );
  NAND2XL U901 ( .A(n524), .B(n523), .Y(mult_x_1_n177) );
  OAI21X1 U902 ( .A0(n1246), .A1(n526), .B0(n525), .Y(n529) );
  NAND2X1 U903 ( .A(n527), .B(n1267), .Y(n528) );
  XNOR2X2 U904 ( .A(n529), .B(n528), .Y(PRODUCT[31]) );
  CMPR32X1 U905 ( .A(n532), .B(n531), .C(n530), .CO(n524), .S(n555) );
  CMPR32X1 U906 ( .A(n535), .B(n534), .C(n533), .CO(n517), .S(n589) );
  XNOR2X1 U907 ( .A(n920), .B(A[20]), .Y(n567) );
  BUFX3 U908 ( .A(B[16]), .Y(n968) );
  NOR2XL U909 ( .A(n1143), .B(n543), .Y(n599) );
  XNOR2XL U910 ( .A(n1132), .B(A[12]), .Y(n568) );
  OAI22XL U911 ( .A0(n1146), .A1(n568), .B0(n1147), .B1(n544), .Y(n598) );
  CMPR32X1 U912 ( .A(n547), .B(n546), .C(n545), .CO(n539), .S(n582) );
  CMPR32X1 U913 ( .A(n550), .B(n549), .C(n548), .CO(n553), .S(n581) );
  CMPR32X1 U914 ( .A(n553), .B(n552), .C(n551), .CO(n536), .S(n569) );
  NOR2XL U915 ( .A(n555), .B(n554), .Y(mult_x_1_n183) );
  NAND2XL U916 ( .A(n555), .B(n554), .Y(mult_x_1_n184) );
  OAI21X2 U917 ( .A0(n1246), .A1(n1270), .B0(n1271), .Y(n558) );
  INVXL U918 ( .A(n1268), .Y(n556) );
  NAND2X1 U919 ( .A(n556), .B(n1269), .Y(n557) );
  XNOR2X1 U920 ( .A(n1108), .B(A[14]), .Y(n597) );
  OAI22XL U921 ( .A0(n1125), .A1(n597), .B0(n5), .B1(n559), .Y(n577) );
  XNOR2XL U922 ( .A(n913), .B(A[22]), .Y(n594) );
  OAI22XL U923 ( .A0(n595), .A1(n594), .B0(n915), .B1(n560), .Y(n576) );
  CMPR32X1 U924 ( .A(n563), .B(n562), .C(n561), .CO(n540), .S(n585) );
  XNOR2XL U925 ( .A(n911), .B(A[18]), .Y(n601) );
  OAI22XL U926 ( .A0(n979), .A1(n601), .B0(n977), .B1(n564), .Y(n580) );
  OAI22XL U927 ( .A0(n654), .A1(n572), .B0(n566), .B1(n565), .Y(n579) );
  XNOR2X1 U928 ( .A(n920), .B(A[19]), .Y(n620) );
  OAI22X1 U929 ( .A0(n836), .A1(n620), .B0(n835), .B1(n567), .Y(n605) );
  XNOR2X1 U930 ( .A(n1132), .B(A[11]), .Y(n621) );
  ADDFHX2 U931 ( .A(n571), .B(n570), .CI(n569), .CO(n587), .S(n633) );
  XNOR2XL U932 ( .A(n765), .B(A[23]), .Y(n607) );
  OAI22XL U933 ( .A0(n935), .A1(n607), .B0(n933), .B1(n573), .Y(n610) );
  XNOR2XL U934 ( .A(n882), .B(A[25]), .Y(n602) );
  CMPR32X1 U935 ( .A(n577), .B(n576), .C(n575), .CO(n586), .S(n651) );
  CMPR32X1 U936 ( .A(n580), .B(n579), .C(n578), .CO(n584), .S(n650) );
  CMPR32X1 U937 ( .A(n586), .B(n585), .C(n584), .CO(n634), .S(n629) );
  NOR2XL U938 ( .A(n591), .B(n590), .Y(mult_x_1_n194) );
  NAND2XL U939 ( .A(n591), .B(n590), .Y(mult_x_1_n195) );
  INVXL U940 ( .A(n1270), .Y(n592) );
  XNOR2XL U941 ( .A(n913), .B(A[21]), .Y(n608) );
  OAI22XL U942 ( .A0(n595), .A1(n608), .B0(n915), .B1(n594), .Y(n625) );
  XNOR2XL U943 ( .A(n968), .B(A[10]), .Y(n596) );
  NOR2XL U944 ( .A(n1143), .B(n596), .Y(n624) );
  XNOR2X1 U945 ( .A(n1108), .B(A[13]), .Y(n622) );
  OAI22XL U946 ( .A0(n1125), .A1(n622), .B0(n5), .B1(n597), .Y(n623) );
  XNOR2XL U947 ( .A(n911), .B(A[17]), .Y(n612) );
  OAI22XL U948 ( .A0(n979), .A1(n612), .B0(n977), .B1(n601), .Y(n628) );
  OAI22X1 U949 ( .A0(n845), .A1(n615), .B0(n602), .B1(n1085), .Y(n614) );
  XNOR2X1 U950 ( .A(n968), .B(A[9]), .Y(n603) );
  NOR2X1 U951 ( .A(n1143), .B(n603), .Y(n613) );
  OAI22XL U952 ( .A0(n979), .A1(n682), .B0(n977), .B1(n612), .Y(n662) );
  OAI22X1 U953 ( .A0(n845), .A1(n685), .B0(n615), .B1(n1085), .Y(n684) );
  XNOR2X1 U954 ( .A(n968), .B(A[8]), .Y(n616) );
  XNOR2X2 U955 ( .A(n920), .B(A[18]), .Y(n677) );
  XNOR2X1 U956 ( .A(n1108), .B(A[12]), .Y(n678) );
  OAI22XL U957 ( .A0(n1125), .A1(n678), .B0(n5), .B1(n622), .Y(n679) );
  CMPR32X1 U958 ( .A(n625), .B(n624), .C(n623), .CO(n619), .S(n667) );
  CMPR32X1 U959 ( .A(n628), .B(n627), .C(n626), .CO(n617), .S(n666) );
  ADDFHX1 U960 ( .A(n631), .B(n630), .CI(n629), .CO(n632), .S(n647) );
  INVXL U961 ( .A(n637), .Y(n638) );
  NOR2XL U962 ( .A(n638), .B(n1274), .Y(n641) );
  NAND2XL U963 ( .A(n641), .B(n707), .Y(n643) );
  OAI21XL U964 ( .A0(n639), .A1(n1274), .B0(n1275), .Y(n640) );
  XNOR2X1 U965 ( .A(n765), .B(A[21]), .Y(n688) );
  CMPR32X1 U966 ( .A(n662), .B(n661), .C(n660), .CO(n663), .S(n699) );
  CMPR32X1 U967 ( .A(n668), .B(n667), .C(n666), .CO(n669), .S(n702) );
  ADDFHX4 U968 ( .A(n671), .B(n670), .CI(n669), .CO(n648), .S(n674) );
  XNOR2X1 U969 ( .A(n920), .B(A[17]), .Y(n718) );
  XNOR2X1 U970 ( .A(n1108), .B(A[11]), .Y(n720) );
  OAI22XL U971 ( .A0(n1125), .A1(n720), .B0(n5), .B1(n678), .Y(n721) );
  XNOR2XL U972 ( .A(n911), .B(A[15]), .Y(n724) );
  OAI22XL U973 ( .A0(n979), .A1(n724), .B0(n977), .B1(n682), .Y(n695) );
  OAI22X1 U974 ( .A0(n845), .A1(n727), .B0(n685), .B1(n1085), .Y(n726) );
  XNOR2X1 U975 ( .A(n968), .B(A[7]), .Y(n686) );
  XNOR2X1 U976 ( .A(n765), .B(A[20]), .Y(n730) );
  OAI22XL U977 ( .A0(n935), .A1(n730), .B0(n933), .B1(n688), .Y(n733) );
  CMPR32X1 U978 ( .A(n695), .B(n694), .C(n693), .CO(n696), .S(n741) );
  CMPR32X1 U979 ( .A(n698), .B(n697), .C(n696), .CO(n717), .S(n745) );
  NOR2XL U980 ( .A(n706), .B(n705), .Y(mult_x_1_n215) );
  NAND2XL U981 ( .A(n706), .B(n705), .Y(mult_x_1_n216) );
  NAND2XL U982 ( .A(n707), .B(n351), .Y(n711) );
  AOI21XL U983 ( .A0(n709), .A1(n351), .B0(n708), .Y(n710) );
  XNOR2X1 U984 ( .A(n714), .B(n713), .Y(PRODUCT[26]) );
  ADDFHX1 U985 ( .A(n717), .B(n716), .CI(n715), .CO(n705), .S(n748) );
  XNOR2X1 U986 ( .A(n1108), .B(A[10]), .Y(n754) );
  OAI22XL U987 ( .A0(n1125), .A1(n754), .B0(n5), .B1(n720), .Y(n755) );
  OAI22XL U988 ( .A0(n979), .A1(n758), .B0(n977), .B1(n724), .Y(n737) );
  OAI22X1 U989 ( .A0(n926), .A1(n762), .B0(n727), .B1(n761), .Y(n760) );
  XNOR2XL U990 ( .A(n968), .B(A[6]), .Y(n728) );
  XNOR2X1 U991 ( .A(n885), .B(A[11]), .Y(n764) );
  OAI22XL U992 ( .A0(n935), .A1(n766), .B0(n933), .B1(n730), .Y(n769) );
  XNOR2X1 U993 ( .A(n913), .B(A[17]), .Y(n767) );
  OAI22X1 U994 ( .A0(n939), .A1(n767), .B0(n915), .B1(n731), .Y(n768) );
  CMPR32X1 U995 ( .A(n734), .B(n733), .C(n732), .CO(n743), .S(n778) );
  CMPR32X1 U996 ( .A(n737), .B(n736), .C(n735), .CO(n738), .S(n777) );
  CMPR32X1 U997 ( .A(n740), .B(n739), .C(n738), .CO(n751), .S(n781) );
  CMPR32X1 U998 ( .A(n743), .B(n742), .C(n741), .CO(n746), .S(n780) );
  CMPR32X1 U999 ( .A(n746), .B(n745), .C(n744), .CO(n716), .S(n749) );
  NOR2XL U1000 ( .A(n748), .B(n747), .Y(mult_x_1_n226) );
  ADDFHX1 U1001 ( .A(n751), .B(n750), .CI(n749), .CO(n747), .S(n784) );
  XNOR2X1 U1002 ( .A(n1132), .B(A[7]), .Y(n798) );
  XNOR2X1 U1003 ( .A(n1108), .B(A[9]), .Y(n799) );
  OAI22XL U1004 ( .A0(n1125), .A1(n799), .B0(n5), .B1(n754), .Y(n800) );
  CMPR22X1 U1005 ( .A(n760), .B(n759), .CO(n735), .S(n772) );
  XNOR2XL U1006 ( .A(n968), .B(A[5]), .Y(n763) );
  XNOR2X1 U1007 ( .A(n885), .B(A[10]), .Y(n807) );
  XNOR2X1 U1008 ( .A(n765), .B(A[18]), .Y(n808) );
  CMPR32X1 U1009 ( .A(n768), .B(n769), .C(n770), .CO(n779), .S(n819) );
  CMPR32X1 U1010 ( .A(n776), .B(n775), .C(n774), .CO(n796), .S(n822) );
  CMPR32X1 U1011 ( .A(n779), .B(n778), .C(n777), .CO(n782), .S(n821) );
  CMPR32X1 U1012 ( .A(n782), .B(n781), .C(n780), .CO(n750), .S(n794) );
  NOR2XL U1013 ( .A(n784), .B(n783), .Y(mult_x_1_n233) );
  NAND2XL U1014 ( .A(n784), .B(n783), .Y(mult_x_1_n234) );
  NAND2XL U1015 ( .A(n785), .B(n788), .Y(n790) );
  AOI21XL U1016 ( .A0(n786), .A1(n788), .B0(n787), .Y(n789) );
  OAI21XL U1017 ( .A0(n1089), .A1(n790), .B0(n789), .Y(n793) );
  NAND2X1 U1018 ( .A(n791), .B(n1281), .Y(n792) );
  OAI22X1 U1019 ( .A0(n836), .A1(n834), .B0(n835), .B1(n797), .Y(n841) );
  XNOR2X1 U1020 ( .A(n1132), .B(A[6]), .Y(n837) );
  OAI22XL U1021 ( .A0(n1125), .A1(n838), .B0(n5), .B1(n799), .Y(n839) );
  XNOR2XL U1022 ( .A(n911), .B(A[12]), .Y(n842) );
  OAI22X1 U1023 ( .A0(n926), .A1(n844), .B0(n805), .B1(n1085), .Y(n843) );
  XNOR2XL U1024 ( .A(n968), .B(A[4]), .Y(n806) );
  OAI22XL U1025 ( .A0(n935), .A1(n848), .B0(n933), .B1(n808), .Y(n851) );
  CMPR32X1 U1026 ( .A(n820), .B(n819), .C(n818), .CO(n823), .S(n862) );
  NOR2XL U1027 ( .A(n825), .B(n824), .Y(mult_x_1_n244) );
  NAND2XL U1028 ( .A(n825), .B(n824), .Y(mult_x_1_n245) );
  INVXL U1029 ( .A(n785), .Y(n827) );
  INVXL U1030 ( .A(n786), .Y(n826) );
  ADDFHX1 U1031 ( .A(n832), .B(n831), .CI(n830), .CO(n824), .S(n866) );
  OAI22XL U1032 ( .A0(n836), .A1(n873), .B0(n835), .B1(n834), .Y(n878) );
  XNOR2X1 U1033 ( .A(n1132), .B(A[5]), .Y(n874) );
  OAI22XL U1034 ( .A0(n1125), .A1(n875), .B0(n5), .B1(n838), .Y(n876) );
  XNOR2XL U1035 ( .A(n911), .B(A[11]), .Y(n879) );
  OAI22X1 U1036 ( .A0(n845), .A1(n883), .B0(n844), .B1(n1085), .Y(n881) );
  XNOR2XL U1037 ( .A(n968), .B(A[3]), .Y(n846) );
  XNOR2X1 U1038 ( .A(n888), .B(A[16]), .Y(n889) );
  CMPR32X1 U1039 ( .A(n852), .B(n851), .C(n850), .CO(n861), .S(n901) );
  CMPR32X1 U1040 ( .A(n858), .B(n857), .C(n856), .CO(n872), .S(n904) );
  CMPR32X1 U1041 ( .A(n861), .B(n860), .C(n859), .CO(n864), .S(n903) );
  CMPR32X1 U1042 ( .A(n864), .B(n863), .C(n862), .CO(n831), .S(n870) );
  NOR2XL U1043 ( .A(n866), .B(n865), .Y(mult_x_1_n251) );
  OAI21X1 U1044 ( .A0(n1089), .A1(n1286), .B0(n1287), .Y(n869) );
  INVXL U1045 ( .A(n1284), .Y(n867) );
  ADDFHX1 U1046 ( .A(n872), .B(n871), .CI(n870), .CO(n865), .S(n907) );
  XNOR2XL U1047 ( .A(n920), .B(A[12]), .Y(n921) );
  OAI22XL U1048 ( .A0(n975), .A1(n921), .B0(n973), .B1(n873), .Y(n919) );
  OAI22XL U1049 ( .A0(n1125), .A1(n916), .B0(n5), .B1(n875), .Y(n917) );
  ADDFHX1 U1050 ( .A(n878), .B(n877), .CI(n876), .CO(n858), .S(n898) );
  XNOR2XL U1051 ( .A(n911), .B(A[10]), .Y(n912) );
  OAI22X1 U1052 ( .A0(n926), .A1(n924), .B0(n883), .B1(n1085), .Y(n923) );
  XNOR2XL U1053 ( .A(n968), .B(A[2]), .Y(n884) );
  XNOR2X1 U1054 ( .A(n888), .B(A[15]), .Y(n932) );
  CMPR32X1 U1055 ( .A(n893), .B(n892), .C(n891), .CO(n902), .S(n950) );
  CMPR32X1 U1056 ( .A(n902), .B(n901), .C(n900), .CO(n905), .S(n952) );
  NOR2XL U1057 ( .A(n907), .B(n906), .Y(mult_x_1_n262) );
  NAND2XL U1058 ( .A(n907), .B(n906), .Y(mult_x_1_n263) );
  CMPR32X1 U1059 ( .A(n910), .B(n909), .C(n908), .CO(n906), .S(n956) );
  OAI22XL U1060 ( .A0(n979), .A1(n976), .B0(n977), .B1(n912), .Y(n942) );
  OAI22X1 U1061 ( .A0(n939), .A1(n936), .B0(n915), .B1(n914), .Y(n941) );
  OAI22XL U1062 ( .A0(n1125), .A1(n970), .B0(n5), .B1(n916), .Y(n940) );
  ADDFHX1 U1063 ( .A(n919), .B(n918), .CI(n917), .CO(n899), .S(n947) );
  XNOR2XL U1064 ( .A(n920), .B(A[11]), .Y(n972) );
  OAI22XL U1065 ( .A0(n975), .A1(n972), .B0(n973), .B1(n921), .Y(n945) );
  CMPR32X1 U1066 ( .A(n942), .B(n941), .C(n940), .CO(n948), .S(n1004) );
  ADDFHX1 U1067 ( .A(n954), .B(n953), .CI(n952), .CO(n909), .S(n963) );
  CLKINVX3 U1068 ( .A(n957), .Y(n1054) );
  OAI21XL U1069 ( .A0(n1013), .A1(n1290), .B0(n1291), .Y(n962) );
  INVXL U1070 ( .A(n1288), .Y(n960) );
  NAND2XL U1071 ( .A(n960), .B(n1289), .Y(n961) );
  XNOR2X1 U1072 ( .A(n962), .B(n961), .Y(PRODUCT[20]) );
  CMPR32X1 U1073 ( .A(n965), .B(n964), .C(n963), .CO(n955), .S(n1010) );
  OAI22X1 U1074 ( .A0(n1146), .A1(n967), .B0(n1147), .B1(n966), .Y(n999) );
  XNOR2XL U1075 ( .A(n968), .B(A[1]), .Y(n969) );
  OAI22XL U1076 ( .A0(n1125), .A1(n971), .B0(n5), .B1(n970), .Y(n997) );
  OAI22XL U1077 ( .A0(n975), .A1(n974), .B0(n973), .B1(n972), .Y(n1002) );
  OAI22XL U1078 ( .A0(n979), .A1(n978), .B0(n977), .B1(n976), .Y(n1001) );
  ADDHXL U1079 ( .A(n981), .B(n980), .CO(n943), .S(n1000) );
  CMPR32X1 U1080 ( .A(n990), .B(n989), .C(n988), .CO(n1024), .S(n1027) );
  CMPR32X1 U1081 ( .A(n999), .B(n998), .C(n997), .CO(n1019), .S(n1043) );
  CMPR32X1 U1082 ( .A(n1002), .B(n1001), .C(n1000), .CO(n1018), .S(n1042) );
  NOR2XL U1083 ( .A(n1010), .B(n1009), .Y(mult_x_1_n273) );
  NAND2XL U1084 ( .A(n1010), .B(n1009), .Y(mult_x_1_n274) );
  INVXL U1085 ( .A(n1290), .Y(n1011) );
  NAND2XL U1086 ( .A(n1011), .B(n1291), .Y(n1012) );
  CMPR32X1 U1087 ( .A(n1016), .B(n1015), .C(n1014), .CO(n1009), .S(n1033) );
  CMPR32X1 U1088 ( .A(n1019), .B(n1018), .C(n1017), .CO(n1016), .S(n1041) );
  ADDFHX1 U1089 ( .A(n1022), .B(n1021), .CI(n1020), .CO(n1050), .S(n1046) );
  ADDFHX1 U1090 ( .A(n1025), .B(n1024), .CI(n1023), .CO(n1031), .S(n1049) );
  CMPR32X1 U1091 ( .A(n1028), .B(n1027), .C(n1026), .CO(n1048), .S(n1060) );
  ADDFHX1 U1092 ( .A(n1031), .B(n1030), .CI(n1029), .CO(n1015), .S(n1039) );
  NOR2XL U1093 ( .A(n1033), .B(n1032), .Y(mult_x_1_n276) );
  NAND2XL U1094 ( .A(n1033), .B(n1032), .Y(mult_x_1_n277) );
  AOI21X1 U1095 ( .A0(n1054), .A1(n1035), .B0(n1034), .Y(n1038) );
  INVXL U1096 ( .A(n1292), .Y(n1036) );
  NAND2X1 U1097 ( .A(n1036), .B(n1293), .Y(n1037) );
  XOR2X1 U1098 ( .A(n1038), .B(n1037), .Y(PRODUCT[18]) );
  CMPR32X1 U1099 ( .A(n1041), .B(n1040), .C(n1039), .CO(n1032), .S(n1052) );
  ADDFHX1 U1100 ( .A(n1044), .B(n1043), .CI(n1042), .CO(n1030), .S(n1057) );
  NOR2XL U1101 ( .A(n1052), .B(n1051), .Y(mult_x_1_n281) );
  NAND2XL U1102 ( .A(n1052), .B(n1051), .Y(mult_x_1_n282) );
  NAND2X1 U1103 ( .A(n1035), .B(n1295), .Y(n1053) );
  CMPR32X1 U1104 ( .A(n1057), .B(n1056), .C(n1055), .CO(n1051), .S(n1062) );
  CMPR32X1 U1105 ( .A(n1060), .B(n1059), .C(n1058), .CO(n1061), .S(n350) );
  NOR2XL U1106 ( .A(n1062), .B(n1061), .Y(mult_x_1_n286) );
  NAND2XL U1107 ( .A(n1062), .B(n1061), .Y(mult_x_1_n287) );
  INVXL U1108 ( .A(n1092), .Y(n1064) );
  NAND2XL U1109 ( .A(n1064), .B(n1063), .Y(mult_x_1_n82) );
  OR2X2 U1110 ( .A(n1066), .B(n1065), .Y(n1090) );
  INVXL U1111 ( .A(n1090), .Y(n1067) );
  NAND2XL U1112 ( .A(n1090), .B(n1068), .Y(mult_x_1_n84) );
  INVXL U1113 ( .A(n1096), .Y(n1069) );
  INVX1 U1114 ( .A(n1074), .Y(n1084) );
  OAI21XL U1115 ( .A0(n1084), .A1(n1080), .B0(n1081), .Y(n1079) );
  INVXL U1116 ( .A(n1075), .Y(n1077) );
  NAND2XL U1117 ( .A(n1077), .B(n1076), .Y(n1078) );
  INVXL U1118 ( .A(n1080), .Y(n1082) );
  NAND2XL U1119 ( .A(n1082), .B(n1081), .Y(n1083) );
  NAND2XL U1120 ( .A(n1091), .B(n1086), .Y(mult_x_1_n83) );
  INVXL U1121 ( .A(n1286), .Y(n1087) );
  NAND2XL U1122 ( .A(n1091), .B(n1090), .Y(n1094) );
  NOR2XL U1123 ( .A(n1094), .B(n1092), .Y(mult_x_1_n290) );
  OAI21XL U1124 ( .A0(mult_x_1_n308), .A1(n1094), .B0(n1093), .Y(mult_x_1_n294) );
  NAND2XL U1125 ( .A(n1097), .B(n1096), .Y(n1098) );
  CMPR32X1 U1126 ( .A(n1105), .B(n1104), .C(n1103), .CO(n1117), .S(n1102) );
  XNOR2X1 U1127 ( .A(n1132), .B(A[23]), .Y(n1118) );
  XNOR2XL U1128 ( .A(n1108), .B(A[25]), .Y(n1123) );
  OAI22X1 U1129 ( .A0(n1125), .A1(n1109), .B0(n5), .B1(n1123), .Y(n1136) );
  CMPR32X1 U1130 ( .A(n1112), .B(n1111), .C(n1110), .CO(n1115), .S(n1101) );
  CMPR32X1 U1131 ( .A(n1117), .B(n1116), .C(n1115), .CO(n1127), .S(n1113) );
  CMPR32X1 U1132 ( .A(n1121), .B(n1120), .C(n1119), .CO(n1129), .S(n1116) );
  CMPR32X1 U1133 ( .A(n1130), .B(n1129), .C(n1128), .CO(n1138), .S(n1126) );
  XNOR2XL U1134 ( .A(n1132), .B(A[25]), .Y(n1144) );
  CMPR32X1 U1135 ( .A(n1136), .B(n1135), .C(n1134), .CO(n1139), .S(n1128) );
  CMPR32X1 U1136 ( .A(n1141), .B(n1140), .C(n1139), .CO(n1152), .S(n1137) );
  OAI2BB1X1 U1137 ( .A0N(n1147), .A1N(n1146), .B0(n1145), .Y(n1148) );
  XOR3X2 U1138 ( .A(n1150), .B(n1149), .C(n1148), .Y(n1151) );
  OAI21XL U1139 ( .A0(n1160), .A1(n1263), .B0(n1159), .Y(n1239) );
  OAI21XL U1140 ( .A0(n1246), .A1(n1164), .B0(n1163), .Y(n1166) );
  OAI21XL U1141 ( .A0(n1246), .A1(n1170), .B0(n1169), .Y(n1173) );
  INVXL U1142 ( .A(n1174), .Y(n1182) );
  AOI21XL U1143 ( .A0(n1182), .A1(n151), .B0(n1175), .Y(n1179) );
  NAND2XL U1144 ( .A(n151), .B(n1180), .Y(n1181) );
  OAI21XL U1145 ( .A0(n1254), .A1(n1257), .B0(n1255), .Y(n1202) );
  AOI21XL U1146 ( .A0(n1205), .A1(n1198), .B0(n1202), .Y(n1183) );
  OAI21XL U1147 ( .A0(n1246), .A1(n1184), .B0(n1183), .Y(n1186) );
  OAI21XL U1148 ( .A0(n1196), .A1(n1193), .B0(n1194), .Y(n1192) );
  INVXL U1149 ( .A(n1188), .Y(n1190) );
  INVXL U1150 ( .A(n1193), .Y(n1195) );
  AOI21XL U1151 ( .A0(n1205), .A1(n1204), .B0(n1203), .Y(n1206) );
  OAI21XL U1152 ( .A0(n1246), .A1(n1207), .B0(n1206), .Y(n1210) );
  XNOR2XL U1153 ( .A(n1222), .B(n1221), .Y(n1327) );
  XOR2XL U1154 ( .A(n1227), .B(n1226), .Y(n1328) );
  XOR2XL U1155 ( .A(n1232), .B(n1231), .Y(n1326) );
  OAI21XL U1156 ( .A0(n1236), .A1(n1250), .B0(n1251), .Y(n1237) );
  OAI21XL U1157 ( .A0(n1242), .A1(n1241), .B0(n1240), .Y(n1243) );
  OAI21XL U1158 ( .A0(n1246), .A1(n1245), .B0(n1244), .Y(n1247) );
  XNOR2XL U1159 ( .A(n1247), .B(n1249), .Y(PRODUCT[40]) );
endmodule

